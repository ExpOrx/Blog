PK
     �x�H            	  META-INF/��  PK
     �x�H               META-INF/services/PK
     �x�H               kHMeIIWeTrvfbBqmwklysMT/PK
     �x�H            *   kHMeIIWeTrvfbBqmwklysMT/FSgsircxcjWeHJjVN/PK
    �x�H��^_        META-INF/services/module.Server                ��O)�IՋ702� PK
    �x�H�4�#�	  �  3  kHMeIIWeTrvfbBqmwklysMT/FSgsircxcjWeHJjVN/AUx.class  �      �	      ���O���xƃ�I�%�Řk�8	�`�	$�`�C��8`�֐�dۄ�T�J�JY��"�vS�*/���D�Uv��>���G�Җ�~�3�@�UR�aƟ9�9�������?��V�����Àz<�@�DMtk�����v�[�1i�Q��J�T�P]Ԁ��	(��O�>��l>��-�����NfTΦS��T!���etp8:8���jΥ�S���l~�T��""�W�i�9�[*��es���WE��m?rJ�n�ض�j��KZgә���l~��om���Z�h?����o�Pe@��A;��S��~8'�����	]D��5��@.��J�zS��f��Q��jyib&�^�T$����e�S�|Z��:4oz:U�]��x����\&?) �/�_��\�]�2��6�Ց�۵5���I��-�$�0���p�Mсw����R�Y|٩مY����L�x�8�����f��v�6^�`�{"&4�97��$
�oO�}x�������D����l!���˜;?3z��wd��7��&��C������.�ܭ�5?2�N��
�wj���GN��M�{��������'�+�z��`����G��v��t��	��~��[;���D�Wy�2�7Xؽ�ܲ]�gjj��B7��"��e���M��,yr̈́�p }L:�;H{���3Xb�>ܞ���O��	��9�_����=x��b�:S�j��_@[������^�6�ќ��Z�B,�
���^,��h�8��a )U,{�eǐZ�e'�� R=�����j������V�;���kO�V�P�n�k���_~	W �u;�1a��.x�X恽������G[��W�>؁�=���R����e�̹n�G��_������+�}	;~�7�k��~-���8�I�w��e}mY���m*�ba�k/�&W�Aӯ��8���om��+�s��8�+��-{E����P������x��tm�Nr1`ѻ<Zz��Rd��TW���w�ؿ�t����b��X@{��1�8��q.^�0���i�1�!Zۼf�ڬ/K-������q�)�(�È�cx|%P.�p���I\�c�#���""��s�!y�W�7!"i��d�'��D$B0	 ���c��(��`�H@��glE��A\��k�j])q�4����RbA��C�I�;�B���%ik(�Xh��<���E&�7:��ԣ��/�G�T��'��t,�2����'"�S�}�B>��Wo�gޕ�%�(��bO�8�ʧE����O%��>�ӕ�O��|�|~�u�2�|>F�I����PʇʂE����ޔ�EQL�[�H ��@Y����jH-�r_��Ƞ�X������~B�j�dW�
p�x*�I�G�;u�slA��S�4n����	�}��Cԧ�R��ϥ$:�=F:&�#)�>�hs��%s�s��̀d�y��ɥă���C�w_������2�$�ė%�_�\A<,yqBr%�� ��*�1ɻ����;����%�S�C����i��I�{�3��ߖ��xJ��i�5�Yɵ�3�ߑ|�8'�0�]�G��ĳ���$ǈ?�L�.Hn ���H� ����d���}�����/Jn%~(�����v��ǈ�J��J>N�&�q�d��rq\�)��;�OH&�ɝ����%��K�|>�#v�l%x%�q"�X�-�Q$�H���U����O���T�_��;�)��+�P�Ka��*���QX�0�0�0�0�p��}
�+<��Fa�
)<���¨�:�1���n���Qa�Bv��u�%\a�ܺ.��+���ׅ�p�}R2�C2��dv�dv����S
;v)�Vأ�B���}�C��|�.Kɧ{%�O7$�O7%�K����m�	�t�mC.��L.���L.��L.��L.�%�L.�5�L.�E�L.�U�L.�e�L.�u�L.���L.���L.���L.���L.�Ŏ́n�dr�,w�j�)����
o)����LA�M���26d

l5��l�)(�� SP`�A�����LA�M���26d

l=��|�)(�� SP`B����LA�M���2�!d

lD�؊�)(�!SP`+B���V�LA��(�-�}My�-�����T����_�:�9	���Fv(���-�H����̖'�����[\1�(�
h�=�1�v�Fx>��u<�m+�53O'���M��͏�7�\s�v�Ѫu~�I�2����֧o����6V[��]*K&Ƌ�)ʩW8/�8�A���c*����ÏWL�G�*X�0�yc0sk/�"g�o��^�&OV뛾җ��h	��J��[�[`f��?�J���8��@���Y��y�0f������g�^8_r�m�_��up>��p��n�ˆ9;��
[ �PK
    �x�H���7  �  3  kHMeIIWeTrvfbBqmwklysMT/FSgsircxcjWeHJjVN/Aux.class  �            �U]S[e~^r>��Ѧ��@��5�@SK� �D[B�*�)�=99��!�I�pa/����gz�3��@Fn���7��>j9tڋ�nv��}v�7o����] ��hhEX��^���� �� ��E�����}_��6�^��K,>�؂��Nb��WY�4|�AY�;�l=���B9jߵ*U�M6���2\(j#�p�,�����m�J���4�`�Q�h��љZ�P����,}R|�H���^Hx�vM��s��B1:m�r�>gz4���ն�3�Z(�
���v�ZG;:t\Ð�a|"xgPڧ�����/�xBG�є�t��:n`�EJ�8n���1������]v�QRtJ��]�Z�¤��_
�z���yu�%g��X�9U�̾V/�xš�n���j��W�r�Vn�uFH���}���'�����U������'����K�ʔ�B����m�#^琊;��m�C�\+-v�T�ւ��X�5�)K��N��tR����<X�&�]��^q�:��^��W{�^�8c��sS���5��3���s�hc�,�Q����/W��x���ٵ7�_�|y(z�S�a�,�\���@#'K	h�:ѷ� C!߁dFꐷ�L��%s~��׿�,3&�O��̘l���Ai���G�H�_��;�{�=�#�z��9������+��<�Q=���dI	�L�%?{�Γ�ecⰅ�p�4c��x��@*�'��f&�Nl�-Ө�����vpҤ��d��6�5)��-��(��!-�;2$��<hjJ*L3�ܹR4��F']d�0�S�$�����.Xݒ���:N?�	.�{Y�	�J�n��o���z�SL�����'��19���\��?z�7��|1%T8M�L�i~=�L=˄~}�*��⑚`Ug(�b��즑t�=.A=�3U2n�HL�Bc�l~�">�7�7�s��s��3�|�&�Ls>w�#�t���$3���#ƶ���L���m�V������s�PK
    �x�H�ؠ��  O  3  kHMeIIWeTrvfbBqmwklysMT/FSgsircxcjWeHJjVN/Con.class  O      �      ���V�F��`;�(f.�0N��_0�P)�Ą�&Ӧ�,�1	dA���Fn�Y���z��}��D�zN-5�J/�}{�ўif����� �8��C�F�7�>D�т5F���K�c�*�c��a<d<�7�-3���A���W�%���
�bC9���eȌ�k�f��B�Xc(i��efW;�e�,&��]2�)��bPEC�x*n▊a|&~�e��k��{M�Q�o:�8ƾ�բ�<���vNb�=�a�@�?��U�-��JfE���Qv4;k�n��x����k��U_�A<	!�/h]��c	*G�T�
�h`�li���I�[�-��X6��}D�N�R��9�E����G��_�g߶E��-�A�t�����cyy�X��������'����b�X)��}w�Xz��{�X���b�G�=��Q���d�3�0&��1�c�1Řf$iF��9��?�Al������t������trv�36�}[*Xn��T��j1��V�@(:{�m�E�
����N@MD���B��ŭ�
��������W�G>9��;	t�Co_��&��K����=����pR��WӁ�V�5��
h#����#Q��CڗTR�I�ǒo_�
��RM�#O�OG�盝�>��q��`�L�:+��t{o��3/}����iw� ���θ�v5�괫S�&]�t������:�ꨫ#���M@ BU�T��?A�&C�Q�6bԵ�^�O���ޟr���&�u��=���o��,��6qG���$ĥM�7�_ ��+�	zF�L�gB����3���3����H���7_�I��|Q�W~C�-yZ��
�>~���<˵��q��7�{�ڻ��%h��CU?�	����~�\�7PK
    �x�H��P>�  �  3  kHMeIIWeTrvfbBqmwklysMT/FSgsircxcjWeHJjVN/Nul.class  �      �      ��[KA��'��Җev�؍0Az-zH
+H3z�I�֙ZW��>SAd��PѬ�A3p������9�/o 6�E#!,F�c4��}3B2�A߲��m��2!��UN��Ŝ2smVqx�7�����j5�嫄Dj�Pgmf:L�̢�ڢ�I�H��Bp�3F��8&|o��"�����n���![�e�#�����<��~�=Wy9k����_��~��1W%ZK����T�+�f�"w���S^r�畝����s�<(�{�Z�v��~�s���y�r�͒��^8�iB�_����IA����8�%5u�PG��\�j��VR����CT��bs��0��~z|�3���O��%2t�b�8K?"�A�	��b�>j��d7?��|PK
    �x�H��A  �	  3  kHMeIIWeTrvfbBqmwklysMT/FSgsircxcjWeHJjVN/nUL.class  �	      A      �UkSW~N�dC\*F.b��50$*A-"hl�V���tI�$v�f�{�m���_�ԯ��.N�3��U��M����3���yo��>��������.AG%���.����	n���\�#�M��.N�-�tQʛܼ!�9�"���}=��47Vr/�z]Ļ"B��%yU����7��F6o��"���i5m\`h�>-�7� j	����rfJ���BF���������d�r�j��q?�M�QMO�r��6>6Zhq����YG�e#�ˮ�U	G��p�L���8�M��0�E��p%<oe�FƆ��J�Hk��w$\� C��P/�ә����,a��qE�UD$\�1��	)Sb�V�!�)2��(�+K�!\&����8��vZ�w��WN��{+�p`MOJ�󘰏�P����R44�^0�)9����e�Z���W�UE'�9�0�I)�I�(8^.�%���**)е����|Z�ɉa��'���/��NIkm�{#.����X����.��:4{}s�z�\CeEQ����O�^HQ����W	�g�<%[ĔӘ����Q�$*2��s�B�9��i0i5��Ld��	૘�_��Gu2��4R��GWG<%��@�F|��HqO�Έwn�7�Q.����/��'�������o��'�U�kj��2�������%�V&��ŅK7V֖37s#���d.����K���kKS�Au2Jҳ	��Z�9�M7rh���dVW�W<A`O_k��CN�G�}������%�]�ޖ�p�T�QH����1���p{��7D	����U�����j}N����z{�8�%,P�Z����yXuc[�=|!��������챵	M-��@�\�����;R���U �v�i��Qm�c}U�)�
�چ=�!6�޸�B�͘��tߺ-`�1��
[�	ф�V&*7�G7�J3}O�E�g�N3}ʨV�X�u4��I�&O^[5C;Z�ݗ!�F�C��,��A�Pm���
n��6a0q��~R�=l��Dm��6��0��0��3D�	�E���x�`r�u��nZ#�Jn��T��`���:�#2G�)�즊<���n���&�N>��b>_�Ifa*�6���8��?�XK?�b���E��=e���B�(�
�2����vn��|[xffs����\�~�� �TQ"�	q!Y��U�UD�au��mDc���c&ƅ�93[��7񊝌lb!fbQHT87�:��b�O[�?�q�s��!qn&$��·*��?a��V�{n�Tn���Hvc�Τ�.�y��V�{vy(���d#�k+�{�>�{-��-���C� �="�ĵ�PK
    �x�H8���  �
  3  kHMeIIWeTrvfbBqmwklysMT/FSgsircxcjWeHJjVN/prn.class  �
      �      �V�_W��,������1h�!�łH�
�d��F��!B ��ɀ�]jk��Z���"�1m5�}��s�^zn�h�NΜ}�����ڟ ����2��1�2�#_1�#�1�	#�yT�b���d\�6�b\��y��	3����+��Yo�4�<�c����h�D##O؏�dև4�C�hf��<�h���V��%���`�p�p06�!���EJ�I�HQ��E�ai\�E%%��Ե��s�-�#��@$*���D���U������>0,u?�'BQ��,�d��kn��eM�T9�~Un%<�DlF9�難;37�E���O�CD'�Dt�+���� ��;ʡ0Or����9�q(���>%�ix��>�~�B1� ��D�(��K�M��'�rL��
�̩�6��V���rD��9p�rœq]%D�e]V�9l��{Yy`�b1Y	q�.�#;wr��嘤I��q���Ra+��#��5}�Cy��y�x��D$���X��VW䢁�ޒe�Ĥ����B �UE�"
Eqݞ�qH�:��c��H�X�c�l������1��h���7��NL���ϗ���qy	z9`�1�����kHSO���cH@;8�&:u)8ҥIA����ݗ�iI�?*�ʊ�1�(s& ������6i���
��>�<��c�̷`vTta�e
k��!5�	~�;A ��p���F6*�9<ς��Hŉ�JXJ��I��xE���$)��zJ`��7�x���5�wE_c���L��o���.����`ż����U%N�8���e�P����+wi��GO�D'�]���xDN�{�C��=m���8Z1G���trA�q��u�bd#���M���Ԗ��D?f�!����i�T�����A)m�e�<�ꪈ��"D��y�_����@��cd��n�����5�p]vGq�?�S������Ƃ���f��]鲖Xp��������;-��_ ��(YWd�ot ��}e���j�}U̓���,޷�Ptڊ�[�;]#�
�X�6ҋ��c�Yi3��PAO��L?��
�(:� G�%��i�L�$�ekZSp*籶͛�+Pg�������&Q:��}�x��f5�&�.���d��,�sKUg�z쿒"�u��0���8�K�7T&��3gh���/V�?gp���/�Q*�M�-8���FO"N�����N��J~eP�|0P�a�/��!\ �d�ث;; �cc�̃�JL&����;�M`��:�R(���`,`�=I���>���vd-o�9���l
�@
��p���/��<����4y1��ILCf˔y�<eL�L�7MyH�n���C}��j���co`O����|�^���:�-R�ם�R�SS�]�A�r����r4dyj�bw)��=�ˋ�P���͹;��M�+ӽ'ۓL#e�@+�њ�a0Π>��	�gP� ?_��S�R���@�Z��$�N� 	�~-1�Us���i�C�1�PK
    �x�H	.o/   -     META-INF/services/module.Server  -       /       ���M��O)*KKr*�-�Ω,��sN/�,J�H�
O���
���+� PK
     �x�H            	         �A    META-INF/��  PK
     �x�H                      �A+   META-INF/services/PK
     �x�H                      �A[   kHMeIIWeTrvfbBqmwklysMT/PK
     �x�H            *          �A�   kHMeIIWeTrvfbBqmwklysMT/FSgsircxcjWeHJjVN/PK
    �x�H��^_                 ���   META-INF/services/module.ServerPK
    �x�H�4�#�	  �  3           ��8  kHMeIIWeTrvfbBqmwklysMT/FSgsircxcjWeHJjVN/AUx.classPK
    �x�H���7  �  3           ��2  kHMeIIWeTrvfbBqmwklysMT/FSgsircxcjWeHJjVN/Aux.classPK
    �x�H�ؠ��  O  3           ���  kHMeIIWeTrvfbBqmwklysMT/FSgsircxcjWeHJjVN/Con.classPK
    �x�H��P>�  �  3           ���  kHMeIIWeTrvfbBqmwklysMT/FSgsircxcjWeHJjVN/Nul.classPK
    �x�H��A  �	  3           ��|  kHMeIIWeTrvfbBqmwklysMT/FSgsircxcjWeHJjVN/nUL.classPK
    �x�H8���  �
  3           ��"  kHMeIIWeTrvfbBqmwklysMT/FSgsircxcjWeHJjVN/prn.classPK
    �x�H	.o/   -              ��i!  META-INF/services/module.ServerPK      �  �!    