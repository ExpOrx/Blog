PK
     �d=I            	  META-INF/��  PK
     �d=I               NLPaDgKCzmcxbojyd/PK
     �d=I            ,   NLPaDgKCzmcxbojyd/afoRIZwlznmSLehmfLSBTAPbP/PK
    �d=Ia?ݘ  �  5  NLPaDgKCzmcxbojyd/afoRIZwlznmSLehmfLSBTAPbP/AUX.class  �            �U]SU~�d�����h+V!@1�Rm��|�)D���V�$'a1��dS>��g�\w�K�Lu����{/�����l� �:Ӌ}�s��=������~�3�|��}��bSFLE }*�1 cP��e�xWE�hŰ
#�W�F�𡀏�T����[>�1.|ܖQ�q��[�4�q�_�l�Pw*u'�T�Ycݲl�g��?��i�����5�+f�23E�$�!P�ۄ1a�~��hڅ8���b9�K���|�Wyn��9^^}ִ���,���4t����Ә[N\73�J��0�i���h��'����I�YoC'cBç�L�L
��a��9�XА���ְ�e�Vd�jX��a=��>���0����*��:����A��K�N}B�X��D=W�iN.���S6�B�o�,C,�)�>�Β�c�`�������@�W�I�#㗻.���Y�l*�����@"BY�Vm�Tqv�S���U�����	�{[k�L͛�v%}����.8^�$�X�߮��
մU���);��P��|�^#�g<Mc�H���뉜�g�J��+�H��*��Ei�|��Z�aX��S�tavj���Δ7wrq3_^L�ow�RZ�����\�HeR��5qGM����n0:5R֬q�B��.��k��o���5�޵�+]��
��-����}�
�!2<B����{ԩ�7ԻK�*<���U��ze;��e�H�XK��M�3\!��s���� `�Cb���X{�� ��O�Uڐ�����Qaq<*�PP�~ �8@�1�B�l�tg���]wq֘�߇\��x�ÿ�"��wNH�P3v"8�D��r� (�,*�0"r��ӞHLFT$���GT9�a��q� �=�#Z�D���q�����yb..F�.:�h�׽Û�	�HT�e�p(�in�d*��#�Y6�F���,!F����E��U���������F���ğ���т
�@����;<GoA��x�� �a7.7�����'/���`?���q/Ni�����'k��]4�PK
    �d=I;����  
	  5  NLPaDgKCzmcxbojyd/afoRIZwlznmSLehmfLSBTAPbP/Aux.class  
	      �      �UkOg~^_��=����.w3��0�7BH��8& ��-;؃156��%M�*����j�~�~m�։�j7j����͞1d��J�yϜs�sg����� ���p`�;T+lXDȊ�0j��u2��&un��4�����jf��C�+E�����C���w�㮶��U�(�0��7�Z�aT�-���j��2�����x����^C��	���P�5�0�f��q(&�b�]�;�����z�4\���`lw�D��.�D���aV����ufN��n����E�<�n>���Z�Eμ]�ސO��j�#�Wkj��1�΍7����i���L,5U��v��#�U~i��t�J��|� �hߒ���4��ڬi�~�1����1�'��5)c����Ƽ��v�k���z��e���0��tC������W����u��VS-�����q�������C֊F�ԧM�|��V*�]cbd�Bb�U7��Բ
X���N�wU�U-)G���H1~��7��o�׊>>��jC�tN}�!��|B=�7;j�� �k�M��&P�E��}�tB�u��r��W�FB��cC�l�pĝ��;�@�<d_�,���_�o�*�M���W���)��c�Z,�)7jwV�U�����~��ڣ�Ɠ��FQ=8�/n\�\��wO^�>�`�������d��ek�w"(.u(=����E]��2�����\b9�=��/$�Y����<��l��1cw,�	��څP�;�LL$E�}N��m1vc'/��1�,�C���rp2$��g�094����<Kl<�O	����ޭ���$ũI�L�mCW��m���D�3qə�}�My
�N�����Rt>��p�}��O,�3م�d��;���������vܼ�Ř�U��������u3��E�����S�B(Z;d�l�/Ϙ��o8�_����i�#N[��QK�(;�-9��V����&��f'��?z��ty�r*���)�~����I���#�o�
�ل�\����ǦR�lxl~�G���b��;O��М5��ف���;�v�S��%���-��b�t%b�9A�3?�)�<4�ӆ:���\n}��3��Z�^s��gp0�y7���]w�5�`���d�?�P.�-Jo*o�0@\�x|��g�ח3&�W���/���0"�k�2 �o�O/]�;�RX=������>ҙq����p��$� ,���>r�[D�tw�v_��W(�>�������1�7lWK!\<���tZcQ��a8GQ:�Y(E�/��I��w��*���o�)�A��
�VLɝn��������p���LU����?7<�1ϣ$-�l�.;�R���N�v��)�nf�;�H>S4���#�[�� ���������|\4pAC�/ﶂ����o����e�����ʚ*��s�7PK
    �d=ICY�V  ]  5  NLPaDgKCzmcxbojyd/afoRIZwlznmSLehmfLSBTAPbP/COn.class  ]      V      �V�wU��&�L�ڡXZ����� A��� ��֦RP��C��fj2����"�w-˴WD���_�9~�x�<�O��ea)���λ���~���0r�s �����X]�%x��'��`垵�E�D��f#W�%l������,�E��<��+���$q�m�J(F;Wd�Pn�(����q�	�<R΍�%Tp���%��&��xN��G�h���'�z\�������7cW~���[�"�6��m<x�����0�۫�T�A���٫��p��M�a�>*�3.ۖ�Ac%�2�������z�Ơx��ڤF�jgHk����I;x��.R��n�������v�F��{���)���:�Tn�Q�Z��ѵ�c�P��]��z���&c����WƝ���j�pt��cl��$��~w����De��؉]��2�ؼf ��A=��*.��R��&�X���]����^g�m���]���XHs���N-� F5à��ݚ����ʱx����Z�
ϻ&D�]���ݬ�1f����"ACko[K?�X;Ӝ��Ţ=��$��YI�G�qq�l�Kc�g�F�(j���=�W�x�%|k,l�h�%*јrE7�`�� ���!�%��h�f�̱i����q����pl��-�[t��u���`8�qF�;s�
�p/[���N=H�e�Qb��$D�Bo��E]ݽ�aO_`�S����Vw譍�B{�}>��ӷ��o�k�lq74���I5��nZu�Z!@d��4�x����L��fp��M��@Έ�X(GD]l G�ڞ+��=�ڷ���̮�+�Aoʙ+:GA�"�۹��r�x��p��W��߫d7�,-)�x�f~���"ޠ�����-^�]���̛#�m2eo`y�}ƴj�`�9D�O�ҩ����R�bɂ�"N�b�g���y{��P��55"���"�,y*]v�|�=����m"���N^\��8�CE"���&勸@w�|U��B�9W�������E�����d)���+T���K��<�B�U��
��&�������!�[N¦��&���øǄȽ'�^�D�	�@&�s�F�	�KL�&0�_5�I����)XỴ)�劤���$H����k$�HΓ��ν\�;ɟ$�m#��@�ߥ��ne������	������>��yJ2��&J�Ɏ�O5F�i&�Ǔ�(Ϥ�`bF<�I�"�ibV<9+��~�n41'�,N��	�5�'-.�QT�2>�k���_	TeR\&��G~�|��N�=���������w��RS拏r)dϵȿL6቏����¶�~���;���b"v%��g�~H<���Z��8�:���Z�0��CƃxraQ�#�?  ����G�n:�IǠ�%��g�@�o!�Rs>��O�S����ש�I����x�P*"�"�d#"�$R�B[*�Y6T�S�/�1���C�T�~��u������ep�7i�f��f≏�9�^�������u�3'�C>,���rvT9��� �,��Y��

3��~0E)_=Lw��V�m�#"\$� �%N�vN�mq�^"��ˈ�q\�~��������:����PK
    �d=I�`���    5  NLPaDgKCzmcxbojyd/afoRIZwlznmSLehmfLSBTAPbP/CoN.class        �      �T�NQ]�����R
� r��B)rk��IcB(��i;�C�ӦL��/�_x&�B$�D��	�uO�	`����>g�Y�\�돏g �x�@=�츎i70���<:����t���a������1��6C{l[ڕD%/.&�唾X�%=�e)f�&Mѧ:}�Zؿ�`���2�+�OI�TT��*���\,i}�:W�H���HpE��w7/�z�gK����ah&����bF�䢒�YYU��eh�)�>��0�f� �.���1�8_N�]ɓn���,�M3������'
�F��E�K2�]�������QM�}�E�m�n���,���C��<?�U�5V�߲j��qz�Kn��]�)���):eM�c`�x(�[��2�"��T9��~����rtcO��r��m��+3K�%1�_ q,E-IM"g)iG0�!�p2�W�)������_A�zz���\�|f���G�&�����&�-,ύ{��6�2�Ԕs�[O�9]�-�L�.��>l3L�;��``:2V��b3�0��x�fG���4W�Ou��)̉cX\�W`}|
����`"d9��-���(綾C����!>��+���k�#����ß����a"�g�)eN���)��A1PA]Bm��fY=�/G!E���YZ�.^���p@���׌�a1$c�j̉�@+�m���>H�0Z�~PK
    �d=I�P�*   �  5  NLPaDgKCzmcxbojyd/afoRIZwlznmSLehmfLSBTAPbP/NUl.class  �             �U[WU�N2�$�҄Q���6܌P/5�V�h�) �P�L�	��I��������4�쪮�.���擯>���3iJt-�>����˷g��翿��0>�ЁA�ź�WqQ�%�_VWѫ��Th�cP��4(HH�CRk��7�xS�����*��(�xG�Ժ��L���Lf��:35g�椝�e�	�G��\�����Ee���"�r�,,����y)��Z�2.�E�
fi5Aw���<
AQ z��1zD9[)g�j�ڮÂ�k��U�rs���*�tt�[��
�����:nt4w�=3L�6l*�:�Ř�0.ń��������#�-L�� �U�t����t�Ň:��M2��g&��ֆc�KǊ�_c������j%�.��ڪ���{S'���Z[VV o��ަ�1�t>}�3��ojh���?����Kj�s�.�B�1
�C����↳�Ѳ���Q����&y��Q�Z�T݃��T�,/�����͊�XS%fU�ϲ}�B��&��Z>2����KR�Y�_&�K͊>�RQ�0[�}��ɽdm
���Pj:5k�\�=�S�ne��۹��/�M-ovJ�t�Z+�S������lbz�@v���	���\�\�,HC�3"��� 8��#�dͪ�ciK�H�&�Xm����)=�M�s�# R�)m��p |����Wn�ߴ7��������d'x@v� X��	`���v��ሤI�	�uD78T�����؇WU��'P(/E����������n��Im���%�Im��c���P��:�M^�Cpڝ�:Z����`��pk�lӫ���;�sR0VVVxS����G}������������0'�nP
M�)t�qR1��(�kЉ��dk�W����}�
���q�2�ZG�q��~xt0x7�Fk����y/)GwS��
E�� [9 ��N4"F��F����6c�<�
>��X������{���ex�?�S"�E&��E"���D��rDYDA�4�������0�<���!�B�1�O�2?���-�A|Ϯ,߭���1�_vuA�wr�?PK
    �d=Iu�~?  �  5  NLPaDgKCzmcxbojyd/afoRIZwlznmSLehmfLSBTAPbP/Nul.class  �      ?      �U[WW��LƂZԨ�F/oH�h�Ė���1�m�F���^��з�����g�j����Y��[W��k��ikԶ���>����{����>��0J�qۆ&���#�^>�y�	��a����4�$#ꎀ!f�Ǩ�3fE�X���+i��&�C[t[�@�Ԝ���VR�RIϗ��^P�0�eB�T}����O��5n6�V��\Jή�UNf�U�0���YY�H�Q�L��
i��ӤG���*3�u�ߟ.�}ھ��EeE)��:��.�2�
%��׷&n���q�<&D�`���U�LIͦ���x(bo�x�x$bQ�D,`Q�����2D<�
CcM���ý����U�*�jV�U�tn�(�(%����V�H�4�/���(C�գa�e�&��9\1�p���whmL���e���hF9�W4�h�R�+��V^�3nP�b(�X�\-��4��{Y�Wumڒ�W��e�-���HJ�
�l�̖��j��͸���8�%:+·�CC��S��R��Ao�:�x�5�]xJ-i�.՛���%�M���btY~���=�I�%s��iI�̭D��m'U�v6������䲴X�R����Y���0&�H`�07E��:�tV���5T��H������D�������\��m#�a��-�u6�{�4I]����ͱ�p���9�L<k�ׇ<V�}�s�qH�)��ch��%�
���?.���|�+�#a|V�Wg��d��H[9��)��p���Ê���\g�������g:�(�z����g�!'y&C���J�!p���-¹}��c���Ȁ����P��x �-g�a�����c��P���N�k�sU�d*�9��V��>�%�N�;�)���R�2�E_pnn��|�,�c�2֝Z%�:��ʰ�S�@`g�
=��x�w*+���?E]<d��O��s���Y3����l�H�A�8���Uß�!,O��2����uz��y���7q���٣�#�'�S��_����g���3�&I���ܢ33~�3���v|�w�ALnbzN#����cR�<�PK
    �d=I6$�S�  7  5  NLPaDgKCzmcxbojyd/afoRIZwlznmSLehmfLSBTAPbP/aUX.class  7      �      �U]Sg~ްɆ�"!)D��!����ѦD!�tټ���n\6���a����W�֙60��tzы�����/�=/6v�"�={���<�����	@?*��͸� ��
�਌7�qL�q2:�xS�Na��-'pRFLFYF7C8}[��%L�*%2�cX�a���a�y�Hl��{�AJ�E.�m]3g4��L�����Z$c"n؉+�ɩr�.C�1\���MF\Eze��8�U�*"�fh{ԥ�a��4�U����Q1(꾫�,���K]_�y�5l��Vv��Z���a&J�⎡'njV�.34����ޝ��T�~������ʺ<���0�����<w-��Ap@�T�E������6OT,��;m����"^_1��9~��-��!� �_7�ej�u7uU��Xvv�=M�1�sq�;2�1t�a0m�O�n�Z�؎ˋϦ(cD�(:�hHW��dM��ź���q����-�v�.��1�%'MmyyR+sI0D�'YƸ�+�,��a�����]􊼏s�FeX��qŨR/7+A���(~]�N�cr��.m�b)7�ٵ�^��i3�R�N��k%�֤�Y䅇h��
�����|�p⥖hX���#�&���N�'�S��ҵ�jY_Y�o?(&�E�fjj�3i�T^Lg.eǦ���,-��GCb��L'���L��W���ī����b��K�RCG�%��G�T����Q�u-�{��0�5Rw[�BVi�n��ph��б��]�#��W{o\��w�<�-��Oh>w������Z��	�g8N_�}�Y(,�%�!�(��G��;��j��M���q��KR����H�אn 1UÍ|9�ؤ����J`-�_���B���ɗ��/�g�badrP.���|n>?:�?�c})}ĞR�B{�0ɵ�/���AΓ}9���G��Ӈ��F?�e3��u|��h�*�\���m^c���'��!�@m�!lo@ۀ��1L��=er�|�:礞M���\~�x��RF���/{z�Ы�^�R�k�[��=o�[����?�+�鋢����{ۥ�Yޔ{�K?�b�O��ۜx}cE:[�Jx�|�K��C'~�NZ��}MܵC"��������ѩ���������3������[��-�	ÿPK
    �d=I`�^  �  5  NLPaDgKCzmcxbojyd/afoRIZwlznmSLehmfLSBTAPbP/aUx.class  �      ^      �TKsG�F��,����q ;deG�@�v�m��� �-IFڱ���.�]�6�T%��r�\��*���UAN�*~ ?
ҳ.���������{���y���� ��R1���8�E�S�>�(�@E����]N��UL�C��+�H�C.�8�sr�D��
>SPW�9C�����x�q�V��4�D3,2�MڮN3�{"r���%2����-�ۼ��0���K�.q� �~�p�\�?p��n˨�^SAQ� ҶC�1J�ϷL;�'x� z�m;������=X�[�0�!_h���������=rh�´�/qQ�J
f4�bN�%�Q���]f��aW\�PƤ�k��a{F�ri�)G���SvC���{��� �W��U_p�=X��qZK�] ]�b����*�z�D7���F�Dl�S�=���;��ܲ��˶��gz��&���T��6w�r��|1��Z��p�&��bC�j��cd�e�\�;r@ɠlp;�����D�ޖ�%�Aq�ؠ&k0�5��*�k]�����lxk[��W���羻^3����Y�Y(UU��ܔ���[���`DkҬ4�(7Q���ƛ�]zc�M*c䘑q�(f3c)ܑ���_H2��ЇJ�B"��hH��O�L��S��л��yT���4�M�AAi�����av7��R}j�����	��]���'nw�t��G������Kyq�p��6F#s3mc �%G�'���].$N$:x�^H�;x{�����Br}�B���y�<B?�~Ñ��;2T�	*bz�|�
��!n4��F'�o?c#�������|�xI"f�����:Nx@�_�{��#Ic�g�,4d�_�t�䟥?�PK
    �d=I\q��    5  NLPaDgKCzmcxbojyd/afoRIZwlznmSLehmfLSBTAPbP/cOn.class        �      �T[S�P�m	�(�TAQ�� ^A�-�J�
���顄I�NHy�?1#�#3� ��
��>�C�l��~���&���`_e���AhB,�x�'zd�-�S!ze<�s	/d�x)�+!�d�#"a@²�(CH���t��킺湦]�`h�4mӛb��_�[��I'��c�ֺ�z��!|n�&~�jᦣΙ�\�+����;��]b
1��y=e�lZy�*��`����8UP'��(x�w
��
>�rw\��Vf^�L�
^f�l�\ϓc�3-��m���y���V�^M�U�p?�hH�^*q���Zq��x�v8�Z��_�נ�=���R�0~�^K{�E�.�/�]6ށ�a9�t��VٮU"�Z�&Cߍ����$������]�a8���
>cZ|"q�I�����9&͆�ڲ��g
��âq�sv��U}�YMm�[�vqM���-m-���si�X��*��G'C��
R�T�DH�B�m ��[FP	�}�+���� 4�HЙ癥]������s&(��ߪ�"�=A�/��b��D�'�*�*h��U;������Rl0K7�
�
�Vqo�hC;"L`	������6f1Ggz0��t7�0�謖�k��i¿m0�������#2]��V��	m�Zbg�iM�?PK
    �d=I��w�.  �  5  NLPaDgKCzmcxbojyd/afoRIZwlznmSLehmfLSBTAPbP/con.class  �      .      �U[WU�N2�t�4J(Zi(����E� 
����$Lf�Ʉ�����|��}f�6�lե��K}�g��}@.i��e�={����Ϝ?���G g�0:t!R�V��� �n	=b=-�W�+
bxUA=�(�qV�s
�8/�!^ �+x�g��~��$\��Ix��]�7����&����&J^��%<��~�p�]�\������]�|�˶�K'"��N3��gi�i��2�9>%��-�$#b_�
�3�L��-;Cy�nԴ�0�]���"Y[�O2TJ���S��Hq�_E;:$���	o�x�24�EV1��-�a��-Ǩ�]b�'aP�5h"Ә�*&W��H���uӘ�0�b��9ܐpS���@Ň�P�*n;��Ȓ���ػ;���)�#�H`8��ec�gf���y6�� �N�`�v�F��}��8�d���<a(�m4G�ھ=�K�d�Dj�7Z����v�gzw?�Dj:Č5��ڜa���eӁ��:���H���U������Q�E�p���eE�5j�MR~��v��n��*q��5H���V\^�&��:�ޡ�'�+r���U+��j{�=&�]��6!"����t�T��U<՘=$T�D����$	�������X4�,�pF��ƕ̵ᕼ��t�S1#�L��-�V�|B��|ZKMƓ���ct[5�	��i�
[\�4�Tdp�!v����#���0�}��N����O�d��Vb�:O^��	)��d|F�]�q��)wɜ8��%:����kd�V�1$
ߴ�H~� �D/��:�}���I��a&�N��:xB��a-C�C��^�)CYá5�c��xN��{�h���8|��Ч]F�}�}N�����[?m<�S�B_T|M}���}�/��M�D�2��VF3�p����WX���Ʒ3}2)a��w���*���xBe=�ϕ��}���%�cX��rx�|#�y���� ����B�<N!H����*m�D>Z[z��B_u��Q	��=����fj�]4��eUl̈́�F+�PK
    �d=Ih��s  �  5  NLPaDgKCzmcxbojyd/afoRIZwlznmSLehmfLSBTAPbP/nuL.class  �      s      ��[S�@��mӆ Xnr��mEx�"��j�2Q�A�4��t�iR�<�=��a��?����> 2�<��={~��lv����4Ve��;B�G�-�Jx��>���`�7���!ܑ0,aQ�]�м�mo��9�b$E�b�j�4�-�h���CX�U^�s���2t��Z�84T��9U��6��1DO
�-�Spm
F0*aL�8�)�!� ���ބ�~�C�&L������j*�Z6����� �%�Ru�xh���<�s�4Q̩yWp���^Kg�$Mut\�N���]�<�C����DQ�ڿ*j\�wS�e(sH��j����t�_���]��:�?���E����hѤ�J�Uny��:��kzu��z��EiLG�th�Wu|�%aA�#�Kx!�	���0��i��J�u�`�3"�9�{b#���9�]��{������YWyI��X�Q.���Lõ�a�Am7޼k�X*�$��	j�~�/�7�Xb�vgZF�Ca$1L7��h���`h��(���Pt���ь�&Y���3<���uN����)X��]u`�^�&'��)�r��'h����l'���p��)�m�����1"'�+�Z��1LЅm9������A�K�͂�Z��6T��KC�4�/PK
    �d=I��1R  r  5  NLPaDgKCzmcxbojyd/afoRIZwlznmSLehmfLSBTAPbP/prn.class  r      R      �T]Sg~^����#�"��Q�H����(Qы�+���APk�io�Wz�L�N3��uT&g%Nk䢙�=���x�9Ͼ����Ͽ İ��	�<��C<|���a��Q���Ÿ���#�prX�0����'�T�����j�Ze����jj+�����f0f�eE/�����T�bU�낡���H�<{�\�KkjU!�;����R����4���ǐ�~��9�0��P+m�Z��Q��1+`��':�S	�3��xٗ�g%��R�4��_��aS�˔�n�U��hJS-I��V���ձ;=uv�S���;8�P"ؖ�Wj��c��]x��;W�G'�,7�F3G���{�/<��U�]�/�uөN9�R�~L��.+m��׼��ͷ�0���Z��c:7�r����܏��y�E�V:+֏~.K�A}3�wZ=�j[9�v��Z�?�(nH��F33���ϒ|�XAR@
.�[��׻�XAݩ��т�~��ܘ8�<^}��.1cLy�z�*�ѡ���w�ۊ��gĐ�l�$g�El�kQn>e�L�o�����B�r��G���OA�;��_�cB2o�7�&L�%�y�J�J�{ۢ5��ጎ����L�s����y_"a�v��.�?�6�CcR��I�h�Kˇۭ�dB�̈?�-/�b��Ѿ	�i��7x�)��%O�(���-x�Q�v�t1'��%�@� A���~�=�_:���5z��_c���G�
�+����M��vW����%��?` ��u>/�_�v	��;;���_���~�G:m�K�]H��b�t,�s3�◱b�m ͇C{W``�З�A����n|V�w��>PK
     �d=I               META-INF/services/PK
    �d=IBx1   /     META-INF/services/module.Server  /       1       ��	HtI�v��M�H�ϪL�KL��*ϩ���I��M�	v
qH
��+� PK
     �d=I            	         �A    META-INF/��  PK
     �d=I                      �A+   NLPaDgKCzmcxbojyd/PK
     �d=I            ,          �A[   NLPaDgKCzmcxbojyd/afoRIZwlznmSLehmfLSBTAPbP/PK
    �d=Ia?ݘ  �  5           ���   NLPaDgKCzmcxbojyd/afoRIZwlznmSLehmfLSBTAPbP/AUX.classPK
    �d=I;����  
	  5           ��   NLPaDgKCzmcxbojyd/afoRIZwlznmSLehmfLSBTAPbP/Aux.classPK
    �d=ICY�V  ]  5           ��;  NLPaDgKCzmcxbojyd/afoRIZwlznmSLehmfLSBTAPbP/COn.classPK
    �d=I�`���    5           ���  NLPaDgKCzmcxbojyd/afoRIZwlznmSLehmfLSBTAPbP/CoN.classPK
    �d=I�P�*   �  5           ��4  NLPaDgKCzmcxbojyd/afoRIZwlznmSLehmfLSBTAPbP/NUl.classPK
    �d=Iu�~?  �  5           ���  NLPaDgKCzmcxbojyd/afoRIZwlznmSLehmfLSBTAPbP/Nul.classPK
    �d=I6$�S�  7  5           ��a  NLPaDgKCzmcxbojyd/afoRIZwlznmSLehmfLSBTAPbP/aUX.classPK
    �d=I`�^  �  5           ��W#  NLPaDgKCzmcxbojyd/afoRIZwlznmSLehmfLSBTAPbP/aUx.classPK
    �d=I\q��    5           ��'  NLPaDgKCzmcxbojyd/afoRIZwlznmSLehmfLSBTAPbP/cOn.classPK
    �d=I��w�.  �  5           ��*  NLPaDgKCzmcxbojyd/afoRIZwlznmSLehmfLSBTAPbP/con.classPK
    �d=Ih��s  �  5           ���.  NLPaDgKCzmcxbojyd/afoRIZwlznmSLehmfLSBTAPbP/nuL.classPK
    �d=I��1R  r  5           ���1  NLPaDgKCzmcxbojyd/afoRIZwlznmSLehmfLSBTAPbP/prn.classPK
     �d=I                      �A?5  META-INF/services/PK
    �d=IBx1   /              ��o5  META-INF/services/module.ServerPK        �5    