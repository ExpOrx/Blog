PK
     �n�H            	  META-INF/��  PK
     �n�H               QVPVaobWbVTFtfGqxSePn/PK
     �n�H            )   QVPVaobWbVTFtfGqxSePn/sDYozveMUDUjWPEYCF/PK
    �n�H$7�	  {  2  QVPVaobWbVTFtfGqxSePn/sDYozveMUDUjWPEYCF/Con.class  {      	      �Wi`W��%kW�ڱ�S���4I%Y�rծ%��v���R��T�B��F�+K��r���rS�&B�e��V�h�R(-��\�j9���h���rp�}���f�̬���>`33����؂'\i��8i��ǉ߄����*{t�`�
]���=|�ˉ&�gB {��>W��5&�����D^�-�Z�܋�~NL�b�~Ͱa�����u���AČ(F��b��7U@���6��A�}\���C&����^�|W��*ۇ�1���w�+��:�P;՘"�x��HHm`��]L��ào�*����c!�?�tq�P��ˑ��tB���cY�&��h,��G#�]���)w�/��?h���C���l�X"B��ERFnpFG�-aeD�p��y|?�@L������w���ݣr,����с�mJ�J�UP�1�t���آ�=���S�
s��,iʊ۾XNB�3eɝ��vNn�p3�!��ޅwKx���Ѷ�e|@UCQ�Z�B�x�W��P/���E��A	�G��%|�p+3Hs�p����6	��)�oK��%|G%|����)�!�-��]��v	�`J�[%|�J�>+�m>�����/☄i���a	_���t,������a������hd(���<s�R:���r~����^gc��#	�q"�f-�s�
.p�����R�g�-�V�_Qj�l����)S³�M-E�Oݑ�Z��K4o�Ҿ�I�-�-��L.�mY���b���`>�J�d�0�8���?��1�Da�ݩ��x�ĸ���%�`*j��l3-4�<:�D�f]��H_�Z����:�(�U�EX:b�Q%�ҽ_q��^�nH�/1��zr�D�.[�J�A�ʉk��,�#���H\�#T;���-s�ZHyQ�[�R�Վ.\Uf�ڗ�
6�MO�ݱ/��0F��9� Ť�>�7ꒃ~yD��$��>��ڕHP�rG_ }H��[�b%R�#�F���'T�^� *�0�e}�7=�����&K�Ms���� ���G'(��@B�ۂ��Y��7�%��*ZX�4в�`���!�N��y����X�ƚɣ��0��H7�ʠ+�`k{5�'�$���}� �|��2�~UOG������jU��<0ީtD����Ę����=���hnu�׃���G�'L�u��C�0�l?=�6(��<��6N�8�pr9�ʲ��ïF��{�^ߣ�3�U箬�n��֊�!���y?&Gp�Y�f����)�D��D��X\X�[+���1:6��*�+��*��򺪍r �~}~�J�PG�V^��"~sA(:_�w�ro�V�g�\~�X��\��ٸ��>;�ZYSdU���]��k��n����p���ʊK+����VQ��yt"��Mc�m}��*�E�sb���Шݡ��W\��+�o�l)��)�Юq�^L��%�HoOÿ�ΘØSg '��:=&���"�0��z�{vr��E���-"c�\�)+�%XLG�(����Y.�'ꍆڢ�"��~�o��"��«��r�z�My���K��j�v�=� r��4ꈖ�	���xX�q�,�#����-�#��ՎĺN���|g�t�`�����B��g���X���'��1���ԫ�d��-䉯)$�B>�Mx�m�tVHr��Dz�PE蚠��^��)t9wÀ<���#p?rN�8Iw�,O��$�x��#�u��$�]�DA�������-?'r�~�3���&Yt5'Q�<��X~M�q��2�G��ϫ3��z���f���]X�!�CF�0%�lڴ�,L�$�nC����,�>	+�V�?����$*I�5���a�.a4��Hx�r�6��@�hf����iJ��gp)}���I���Y�[MڭY���Z�)(V����8��V�,l�I��>��,��'���I���_������i[���0]V)	G_ߍ"+�^	���>�*��8�S(��S�hTҨ�h�I��}���{�=��>������4LTϱ�iM��$^(��V�W�{�5*6�g�:*�s̈f4P�<��Z�(_�3�:Za`x��N���x�JTd�8J%�#�F��f���¸�J�f���J�RA��醺����9���әl������N"�U����L9�� �GHB�K,e���w���y��3V��i-P8�)\��h!-��-�{}I�S���a>�@g+hVp�:�'�0���V���L���k�h'��qH�i��)�)��)�����u���j(�i�vJ`+yh�.m�����Pz��Ԣ����?PK
    �n�H��d�
  \  2  QVPVaobWbVTFtfGqxSePn/sDYozveMUDUjWPEYCF/NUl.class  \      
      �SMS�P=�QbT
bP�J����B��QZ�t���Q�%�4 :�:���u�3Nq�q�?J�� ���Yܼ�s���w��ǧ/ ���	�PѤ��´T1���A-��&C�N3Hq'��f��UL[n�Z)�Ea;��6�zǞ�}���^"��b�g֭-+V��|l�sv~DG4m8)N�:N!����'�Y��nq�:q6�Ǜ��������:U���!�6F���Bđ��n�q�3�d$�S.y�K��=Nl��rW�i������<Uti��	j��.xV�ѢkeIx�����4U���H�Y��s:%ǋV�4gmp�hd�#Y��!�>��Q;�pZ��N����ro����h�1�i�.q�:j$��R��gA�_  �L7�9>�cH�vb�x���{k�[��q���T�h�
ϮY���E\�M��m�#��LO���ork]bGk�-�}j�s�ޙ�00� �L[���Jzq�[��d{�'�Xi�t�o���dj})9eƧcs�"龋)���I��p�}���� �p��@<2��&�ͥ�z3�쀽�-Y�w"�{�s�	�������*C9�8vX�k?��8>z<DEֶ�:3��;�̀d>�@�@��h;�h�<��F�Է��4w�m��L��L�2�\��z2W*�jV0&�@Y�Vʊ�-�eq����2^�r�ѹa5�4,--�c����ƣA)z���u�]� [.�J�^���hP���@(�e�^���<z��u�ft��3|K���t~PK
     �n�H               META-INF/services/PK
    �n�H�sv.   ,     META-INF/services/module.Server  ,       .       K�O
O
q+Is/�N��+v�̯*K�u	�
p�tv��� PK
     �n�H            	         �A    META-INF/��  PK
     �n�H                      �A+   QVPVaobWbVTFtfGqxSePn/PK
     �n�H            )          �A_   QVPVaobWbVTFtfGqxSePn/sDYozveMUDUjWPEYCF/PK
    �n�H$7�	  {  2           ���   QVPVaobWbVTFtfGqxSePn/sDYozveMUDUjWPEYCF/Con.classPK
    �n�H��d�
  \  2           ��
  QVPVaobWbVTFtfGqxSePn/sDYozveMUDUjWPEYCF/NUl.classPK
     �n�H                      �A�  META-INF/services/PK
    �n�H�sv.   ,              ���  META-INF/services/module.ServerPK      #  7    