PK
     kZ�H               HIrcfOqUnFBvR/PK
     kZ�H            )   HIrcfOqUnFBvR/sJmCBUeyDQLXFWznuAJJuRXoiu/PK
     kZ�H            	  META-INF/��  PK
    kZ�H��G�(  �	  2  HIrcfOqUnFBvR/sJmCBUeyDQLXFWznuAJJuRXoiu/AUX.class  �	      (      �U�SW��d���Z�b�`���,bZ��i��
�|��K�!��.&A�Z���z�[g|���2#I)��t�/��J��T2�$�{>�s����O ���Amě���L�gr��w2��qHF���4"�;x���6!�#Lޓq��c�e����|����+�''��#�K�U-lX���%=c�*�t��K�V�%��@�c2.[3.k�邞�j�)�>��Z�0u2��0L��H`_p(yY�И�4heu�����
cZ��&�(��y�,���޺��+Y��JEͦ���ڬb댘9��׵b��I
���O�f�i۰Lr�*��'=�`7:vo�����`�6?R������D��*8�0�J
N�S��(8���a� ���ڶڥHl�C�ّ4s*<���e���7�X0�T?X����M[�~��ȵ��d����n�+�����7ɚ֩���A���m�dӚ)Xeʽ�PTr9�4b\ם1�{"�� ��vn<�M3%��]�@�'�
�̹B����TKs�M/��j�V{a�pse|��.�[�\-iº'JG����:]Ћ�i�*�(;�]�s�����"9o��두�8�/	*#@�u���� @_(�әN��K$�U���0�:��;���{D/�,�&����Lq��l�ݜ��
.��s���(P�e2��R?���]5Ӭ�Bm
��*�,!���|Q��[�T��)�+S���^��M��\�!�����^���2�ؕ�94p�b�<\���N]�&�Ư������ńeT���?�t���	T�����)����5���+t(��v�L�c����Eʫ��^����W����!Z)*���)�����~������H�ݧϘ���䤚|��#H�#��d�+����KhL��jh:���_,`�o�Z�V�Y�k��Q�����d3Oy@�Y4��x��ܢu�&�&�0�b���8 Os#�tu韄���K�%�p!Y��*Ƥ#�*>�ab��I/�\F�
S���$�,���SI�|�UMH���=r:�#M$�z|�����*��w�2�+��;����o�R�n����4dy׳� }�������K(&�k��F �R��T�5�_�Y)&O:���$5��CM�A��Y�w�|�ϯE;J��sp�ݡ����z�&q^��Mc!Q�k�>HGψU��h~�Fr��@�9�s��j-4�_q���"��u�@��L�$�]�'��.�m�]U��RŎ����?��U��n@$����+Pv����	}*���PK
    kZ�H��6\�  0  2  HIrcfOqUnFBvR/sJmCBUeyDQLXFWznuAJJuRXoiu/coN.class  0      �      ��]OA���n�.��~����%�M�CUb���B�LۡYlgt�m�&MI��(�ٖ�E1D������yϙ���,�`!��&�0���#��ᡉ�&��}�˄Q��IHuKr�n�Φ|���/q d�*j�d3$d���i�-�R��w
޾�	�#Tۭ����K6��l<�O�,^Nؘ�E��VԑnU=����El=1p�[i�s�R�f;)�Kܯ�¾lrHV���;�������P\cι��l�Ĭ��!� ��>���^�{M���6܃r��Z��ֽ��֑�V��h����m��ܪ���_mL�9���+��m�\�6ry�&~�T3��+~;�_j����fx$��S�/�l�� �����	0����x,/"���?�����1Fw��:�q��0�O�{��g��K�ߘ�9D�p	PK
    kZ�H��&�  �  2  HIrcfOqUnFBvR/sJmCBUeyDQLXFWznuAJJuRXoiu/nuL.class  �      �      �V�Sg�}�a�(�bbKS/!$�Ֆ*�m@�� 
Xi�K�$����{Ѧh�ӷv|�3}�VC�q:N|�C�����%�"Zy��=�߹~����o�8�oE�b_=��N>�_��K (b��k��aD89("�W�*��9��k>��s�9����pD�UG��YeA��������2���|�1U��f�mPǵ���c9-g�`�
>��i����zZe�&���S��2�WG9!���FQ#��^/�h�(��eҜЍLt��k����A;R�?-z��|Z5tI��^	�p\�	�)�-��H��I	��'�4�04nDah�$(�I�q�s�m		�BS��SK)u���TP���y�P��>���2y(�h�Z�fh���żQ��`�TӤ|�O�լ%�?�x��7�[��W5�<��z���c�`;��B�~���}�șjr��ƷYd��k&_,dZ��]"�-ߘ��P�ԗ�f>!P�!���oQ]S1d��-����4Ptm^�"_cC"�b�Κ���8j()Z�`��#	�T��Ꜫ��we���^eN�0��ϧ8�!c\� ۱T3��m�w��w�;9����"���m /�r��{\ᤃp�1��E�KHCрR���� �`��WB9����'{���M�sɜHߪ�>k"�*�L��'����|!��H8�3q#53t)���,G�s�=Iu���D��e���/O�b4���Ea�-9i�w��G�b�iU.J�̿&��І��vK0�cox+�<]���w�E�=(QF��0��u�uz1}]u�#;<��:�' ���������;Y�p�7�͢�~��"/h��2��j�4��X0�@oP�?V0(WpV^ù2��C�e�_��TD��H�ed�i���^r����⼫"�|��'����c����x�s|J>���r�"iv�|+�J�[�~���wI�M��@�Y�ѐ�J]5�'}���f��
����)W��JtR�X��T��vM�n8H�WH�GN*�����_��!�ax�Y��K?�I=eԗ!�Sυ�>l�;ְ]�~n�6�D�@O����r~��r���mv=������ol�`k�����h*c�j��q�?T��7,Y�j��#�
g�^i@��_�=���hY�D�]-�H�\����I��u�?��O<�e�=:�Z����p�������sK�@�▩PJ�PK
     lZ�H               META-INF/services/PK
    lZ�H��.   ,     META-INF/services/module.Server  ,       .       ��,JN�/�ss*�+��uv
M�t	�p��+u��*���,�K�� PK
     kZ�H                      �A    HIrcfOqUnFBvR/PK
     kZ�H            )          �A,   HIrcfOqUnFBvR/sJmCBUeyDQLXFWznuAJJuRXoiu/PK
     kZ�H            	         �As   META-INF/��  PK
    kZ�H��G�(  �	  2           ���   HIrcfOqUnFBvR/sJmCBUeyDQLXFWznuAJJuRXoiu/AUX.classPK
    kZ�H��6\�  0  2           ��*  HIrcfOqUnFBvR/sJmCBUeyDQLXFWznuAJJuRXoiu/coN.classPK
    kZ�H��&�  �  2           ��;  HIrcfOqUnFBvR/sJmCBUeyDQLXFWznuAJJuRXoiu/nuL.classPK
     lZ�H                      �Av  META-INF/services/PK
    lZ�H��.   ,              ���  META-INF/services/module.ServerPK      {  %    