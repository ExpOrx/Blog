PK
     8��H            	  META-INF/��  PK
     8��H               oztTSYbRWxqJcGzRjtLf/PK
     8��H            %   oztTSYbRWxqJcGzRjtLf/ybpKxWXLYBLlRFO/PK
    8��H�b�[W  6  .  oztTSYbRWxqJcGzRjtLf/ybpKxWXLYBLlRFO/AUX.class  6      W      �V�wU�^3�L��`J[�X[���R+tC([ ��-��i2MS�II&P��V�q7�%�B������?�w�_x4�7i�BM{�}o޽�{w��;�㟟~ЌeTas1��E.���blA���hq���G+_���6���E��t�x_�jtq�C�{2��Í2�]��M.���u�r���"ޕQ��x�� �n�e���G�;ՁI����}�c�F���)��J�T;C�u�ޔ�5;��ꈚQ����s���41�����CzlHOD���1�鬉h���H�$=ܜ�����͈���f�]A�"�*؇�"�
� C����R�X�H(����*��E�)�ǀ�A�2� �a�)8��fX������3�.f���32��h��u��h�1L#��'�XLA`(���S1��o$�	)iX�F��≈o27}�{{�%�r�.�M�й�gi9�=���2l\�f��T��6�0�� ��r��d�[�Y���D ���e�A>�y�x,��`��!�D��i�l!��횴􄵠����!})�䄳�iX����*_Z��q#!��"'�?��E<(C�fb��=��@B��<ם���3��"z���d��swLO&{�)CA�S��&�"�2&1��: c�| �k"΃�8�m�D���4x��a�9S�ǐ��I.�N�0#z��\����'q�Czb���U�����<J]�t7�O����w��t��*4�<?yxg��$���f��g�bT
�x�� 1����5Я��g��훴㾓c�g��mW ַ�׷sp�?�c4tr7J�Q_��x<ʧ��U�Eb��)v9���_�X���b�p�6(x�<���B�)Դ���PSs0V�i��ѹe]iiK�8�q��S�j����歑M�Kf757������p��n����l߾��Mw4*$|T�����]�%|BWFi�zt�Ve����t?�=���귴$f���k�{v;%|NLu��X��^U?[1��w]I��/��Zڻ:[�$|M�c_�Q�/�	���7J�D&�m{?��������u㩺�e��]�r	W��W��Y����W�c�����zKs�,i�5ŜM����wC���y�j�е,�2�G2x(����$�RZ�B�%͹f\s.mF�s�sN%���SІG��HGO�8l��Zg�s�͕�No��V�a9B=U�!97wn��"H��-��k4dy�(7XC�2gg���o�8�y�x�;���I�f�/�ggG\^�i?�l��^F��ͣ�Ҫwxs�^
.�||O�;ס�����znE�O��~�"�++�~���P�"X@e�
��{8���P�X�
�6|E�v�<D��;�8������2߽��+g�*��2(�@ܢu|����h�� ��F��i��z��X��d�&�[ӹ���V
ȭ�	Y�f�6�{ۡfQ�Ν��<�;KSE:�$M��s�ҹKy��6�<���՚Z�ʂ�oϠ6�	\�����߱P�8yQ�/��/�.ҽ�<G�"|�Z����?QiS�E�zq�ve�����j�g�OW�AsE�zd�C=��F]��
�� �Ȍ'��� _��;���tˋ�PK
    8��H]�6 �  �  .  oztTSYbRWxqJcGzRjtLf/ybpKxWXLYBLlRFO/CON.class  �      �      �R�J�@=�.њ��}ߗX�� >(�5�ں<%1���h�J��
n���Q�V�R���;��s�f>>��,b�"�x������SD��i�"z:Լ~�+���#�`�������C0�]Z��3u'�l�p�c��KQ��HhCLD��>�K� CgU���]m�lZ7��Qw�n�y��I��K�[�N�}���H������C���e2�ʍ��M8,x�U,!dzn��H�ރ|tf����=s�!���+�޸�/gOճM�Iok���)wqK�ð.7O�g�3�vNi��t	#�H�0��,��Z��
!��
 �$B�E�3�#FU�NKh�W����V�j�ʠw�"LY�r���0A� �6�~K,#� �-$�/��� � P!�F�!�9Ʃ�l�&!�/PK
    8��H���V�    .  oztTSYbRWxqJcGzRjtLf/ybpKxWXLYBLlRFO/Con.class        �      ��]OA��C��v]K��mo6���5�&�-_dڎ�6�,S�.�M�!���QƳ-ًbH������9?�~XF�A�m,`���Ic(%a��K��P��!�7	�Uݖ�b�["�q(��\O!בf�M(y�+��	���&U�!��{5P�Z�JɖqQ���!�x�'�r�����n�"��e|$c.���!L��گ6�\b-I��{�b���f�d�~>խx���MN!whD���͍�g�6<�<���3�^o4k['�Z�j]|�O���O���ƻ �}��|@�fF�c/������hT);�*}��ͽ|������K�#����wx5�#�\�~���rtI�1�q�X���w���C����2���_kT���#{��OXÎ�����}n����PK
    8��H��=́    .  oztTSYbRWxqJcGzRjtLf/ybpKxWXLYBLlRFO/nUL.class        �      �R[OQ�N[���VQ�{��*^���Mq��TJ}b�.����v�³�c|2�c|�	B�	?����✭ DB�df��|3g�7��קu ��G�2E�q�"<hцvo��q'E��i��,W�8,�s:�	8�������^O(�1N�A3�13��UKW�-��ۚ7H�8��2�ʬ��Fէv4ifM;&��.H��"C���K�,�S�\pM�u�pSB����G�-����ө�rN��u�:�A5���KS�\c�%[+2�s�vJ/j	�P�KN�[}9��j�	�j�͢��oߛ0�KZܘ2)iZ���akV�u�}��H��q/?C=���^�'?��2�C<�I|E�J�\�9ԅ�ά\�92r�Q�@:�s�N�e��t��h��Rr�V���ٹ���P
ɑ�Q�BW�,�*����&�nɴ� �<�N.���A#�up���~��w��d&f>�U�Ih&�L ����dP!Fe#X+Úॕ6�p�}�'���{tn��+p=��Ux!<~�/�����M�J2B2K�2�~�b�U�+����-Kr�UX�|����;�g�ݘ�����W��j�uW�PQ*�T�;~��bڝ�7p�!ƃoD��I�J���PK
    8��H,�;  �  .  oztTSYbRWxqJcGzRjtLf/ybpKxWXLYBLlRFO/nUl.class  �      ;      �T[S[U�vrNNH�m�A.��$c)F���jh�5�K��'�&	��CO��3�����K^�F:u����+ĵ����q�9Y{�u�����g��ϯ/ ����Mh��Az�y �ۃ+�����xQp]����!��s<�PZ@APAH$��ూX��5Z2J�m).�3�%a�4}A�JZV�)!�֦A2 ��4�7��=�"ږI�Y�apdb*|�TV�!"��(�H�MPvݱi��HR3�fY�-���*�B|�O|��㋩��߰K&���u�(D��-ks���� C�|�I=*U���?c�۩ؼ�М۴,nةR�ϔt�T��9}6ضJF��mƊ�5nYڎh[0cP�m�F���u����B��:�*�C��s�!¦E�C��Ll��rK�0C��-1	�������l-���������^�&u^�GT��]�<�H��v���jeJn�3���1��T���1I�
�.��`�O����Z�"�T��=�:C�dT�E��o 9gj���=�#��9��6>sw)�չQ���y�U,`Q|2K�ȉ!��ed��Q k��JXV��T�y��l�lx��X9gڐeB	s�Nͥ�����ӹ���5;���n<�^\J�'zr�aĘ�	�iD��[��ҟF�����4m����_z�Pښ��y�w���s���X�|�5"]+������%7,����JW��9��û���t%��y�R��lK��\�Y{x�g8�~�e��^JGe���1t���ҋ�����
g���R!x�ھ����\=�c��.VO��*܉*�����A$,<����/�L�m�=��@��o�?�TT��N�S��x�|A�b���1�0����Mb/��MT.��1F��#��k��25|v�+5�:I$k�Oא��{Orm�C�^�L��2��"�3��Q%��V�cQye�U�x�'������pu����n� r�������"�'�]���c���ߏq%>��?����Wi%�TL�����F1CT�hZ�?�|��������ir;�I=)�m�zO�_PK
     9��H               META-INF/services/PK
    9��HpK=\*   (     META-INF/services/module.Server  (       *       ˯*		�L

�(�Jv�
�*�IӫL*����t��	r��s�� PK
     8��H            	         �A    META-INF/��  PK
     8��H                      �A+   oztTSYbRWxqJcGzRjtLf/PK
     8��H            %          �A^   oztTSYbRWxqJcGzRjtLf/ybpKxWXLYBLlRFO/PK
    8��H�b�[W  6  .           ���   oztTSYbRWxqJcGzRjtLf/ybpKxWXLYBLlRFO/AUX.classPK
    8��H]�6 �  �  .           ��X  oztTSYbRWxqJcGzRjtLf/ybpKxWXLYBLlRFO/CON.classPK
    8��H���V�    .           ��J	  oztTSYbRWxqJcGzRjtLf/ybpKxWXLYBLlRFO/Con.classPK
    8��H��=́    .           ��Q  oztTSYbRWxqJcGzRjtLf/ybpKxWXLYBLlRFO/nUL.classPK
    8��H,�;  �  .           ��2  oztTSYbRWxqJcGzRjtLf/ybpKxWXLYBLlRFO/nUl.classPK
     9��H                      �A�  META-INF/services/PK
    9��HpK=\*   (              ���  META-INF/services/module.ServerPK    
 
 *  x    