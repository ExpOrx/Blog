PK
     2R�H            	  META-INF/��  PK
     2R�H               _005_/PK
     2R�H               _005_/resources/PK
     2R�H               ghIcrdbadKKutXgMjTlYNdzfxIM/PK
     2R�H            +   ghIcrdbadKKutXgMjTlYNdzfxIM/pojBrCRxzxSdwP/PK
    2R�H�=:N'  �    _005_/Capture.class  �      '      u��n�P��M�	�M���B)���:!�.��EKT�E�+u�ڕ� ʆ��$*$eǂ��9�:&�Yܙ;�33����og �hf�AM��4��Y�AúCCC�}��oy�9�Z�o����S�\�b�u��t��9Yjy���G��P��c��6�[��>2̥�6��섒t�J��r_3��؎�5:�Yގ�2S�}�59�q�T�ۗ��F���2���g=f[�o[�Үv�8g��;F������I�T%Ռ?ɨ��M� ��v�`#�d�eM�r��@n�y}�-��b��|c�Ŝ��4i���q����\��C�/z�V?XS�kl�;���Gc��E��*���~�0����{>��C���\�-12��Z��1�_�̈́�Y\���Z�(�ZT�AuJ�k�S�ϓ�\�-�f>�P���&��� �8H)d)$YdMy
H>�����,%��LI�An�fe
H!Y��<��)������@�P� 5�ԧ�ȿD��z0�
5�j
I�`�NVڈd�K��;m�S��TWBU�PK
    2R�H���ՙ  �    _005_/CaptureMaster.class  �      �      uR�NQ]�---S�B�����[�DkLТ ^ȡL��253Sy�ů�4�$��o~��`\�t,��s.�����k��?_ ��Bq�H��O�b�M ��^�'ps:|3�[1܎��	�v���ڮ����Ň�@�Tw<_:���5��ϩ���} з+�S����k�.�[i�<�tyG�����j���+ߔ���˪��f�d7�|y�P�����&E<�G|_��K-��L�?�R}����r짍�M�]��5FR�z�J��{����ܦ�$=�vI��.ӭ��r�� �dW�/�����v�yI�LG����.�=n~���%:\��p$���!]m���r���?N�ʶS��M�?/�\o���2��6���0�!0naI��.�Z��b��q��I�����6�5�T��6w�/0dB��_6ӥ����iMϔ;3���d�if��8��S��也�� ?V�sJ��x�ć��+����2+�Ӽ�y�{r��t, ��3\�& gq�{��<ct��&y����s����!�v����-��I"$��b�G�@@�".�+�q��MA�Enma�b�$e���Y����lx����>M�E�;��@a������{ė0���Ǹ�-�(�R�+�\�u���^�t�Rp����C���ǎ�ٮ�Wj�/PK
    2R�H�j��      _005_/resources/a.png        �      ��s���b``���p	� ��$��� R,�N�!@PÑ��sxD30p} aF�5&3��2%�%��i%�E��)�I�
n�E���E��
���3��1Չ��9�&�d��)�d�2���8|�&R��c�����2H�"���ƾ� 19;�D!)5=3�VIAAAI!3�V)������95#ӣ�(5��/$�*;�2E�ގ˦�
�97�$Q�"7'�ت�V	l���WR +)ɶU��:�7@�9�(U�D�P7���D��L������LG!8�D�+1O��\��� HYZ�*@����)JI�
rq��	��*e��X�뗗������ZZZ���U�W�$V��+C���Z�\�Y /?1)���VI�K	@=�X �(�x�`�J����M��D~QH~~��H��GW�M������Y�XZD!�(B���V����������I,\���� KI��WAiQ8ZR��SsRsS�J��af�f)�Vi�E��%v�����y�6�A��0Y��ӥ��h��%_�_000�y�8�xt�vЯ�A�m�jOݸ&ۊ�������|��\��jH��(	~���Ӻ&�4�������vl�6���3��RS�m�8s�$��ݳmf����Ss��{C��J�Bi�.�1ux�0kܲ�I�w�	*lBS]'���u7Y�)��2�=p¾�k��<U�'�˞��qF�e��*1&�m]�_jsMZv���M��s�׋"��	O?pf���/�4�Y����+##-����sC@ǚ��=Q�W��1����u�")Z/v0�5V{>5����Q8d��}�ψ�~�)<1qIp�O�-�E�O��ܹD8����فU�|�~��ӑ]빲��������|?�y~J�lVۿܟ,#����R,�<]�\�9%4 PK
    2R�H�>���  �  4  ghIcrdbadKKutXgMjTlYNdzfxIM/pojBrCRxzxSdwP/COn.class  �      �      ��[S�@���&-Q˥x	"(B[,ETT.*T�BAG.R���Y�bH�4h�����/<�3Zqt�G?�~�,E�6Θdv6����ɞ��_�� �İ^���@\���㩏ުT�P�ZC
l��ӛ�r�-w04� ��g�N�Ӻ9��9}���b�{�RQ	UEN24������[�h�r�m/-:�,�����[
N�8���7p<ks�`�&狔/8$��{Yp��+�f��cw윕X��㶂35�T�/�"��p~�c�9z�ٸ��i��P*�W�k���rzT�C�����w�ycT_ �6J\	�̠�CTA����M���AC�A��1S/DJ��,��P�*p�a��G�2�?-/��}���ɗ}*�]WI��V��n�|\E��߇m@�M�q���Y��wĖ�C1���9���k�#,�-GU{�$�����-�͋���Б�d�iۘՍ��%g*32?n&G�Ws��Ht1??`�_ǌ����U?C��ah�c���.!@3�z�TPS�[?\tZ�\oPW��5�OP�k[?��)T��*xhv��L��DkV�ʵA������`Rr�#\�E�]�c����ް�(�;������ �nBKn�lr%��:S%��6SB�����%K��bY���r�L��2囑�T�h����f�}]�L�g����V���>�qy�����l�����C�+���z��>��ַMt'#�xw��U*����PK
    2R�H��9l  �  4  ghIcrdbadKKutXgMjTlYNdzfxIM/pojBrCRxzxSdwP/Con.class  �      l      �V{xSg���N��a	���m�V =�
+��"����hK����IIsJr��Wt^�yٜ��9��m��	�8�T�y���]��L�������'Io�H������/��~9/N?��Z��E�@	��E�q�[��w���'�r��Ì��Њ6�.܋#":Dt�L��.2�m!��S�L���[���^`o_w�N<�r���5ω����c�U������(%䢗A��(�A����PP�_\����-�e�=�*�������<W�}G�^M'�cO<כ��\C�ZN��
����*��"J⨒�+�	��� k*�$�a9w�PBI��H=��ʂZ��7�֒�Cm�yD�y�#hEH�3}�O��f�.&�x���W����:��2��Y¾P�ш:��5��������Q5%b@�	4JH`PB��!���BZ��1	S���X�D���`t~�f��:%�4�$�-x+�o���eM�jm���s�O(�t���2�謈�w�I��b�n�p?�����2�}hZ}g�n<*`���"���[E���Z4�P}jjXM	p�U]������z�:=W�I�R��P���$ETs]��#E�����,i�9���jW����[`�:�ޗȤc\\�|����6���$�e�Q��=�ݹ�Z��%e�y2��I4�qK
b�C,x��پj��i]I�p�Qנ�I����&�'�S�)5M���5�*i�N�>NQĦp�6�Ғ��ʯ��:��x��_��b�i#�t�x��s8@mc��9љR"d��Sݽ �"�@BTi�%| d�(
R�π2�J�0N�3yeu�a|ą����nQ����?����8]i<�V�h5���u�K�}�d�b�Bvj�_��od@�g���YbDbJj��	�>�,s.p�t���SL�����E\��zc�O�e�|���	�&[2�HpG�4�#��8��`,IE{�����X�@g"�=�7h�i�S�#��G;�#��T�_����5SM�E�}ZJ���c�fo�0ɧI��+5�`�5A3�D�
�bt��g��J��Pڒ+T�V�@5��i����۽^'~HiW;�c�����ȵ�vn��8�s��;jwVmp�$�͉_ѶՉ�cc��R���J�wU��ܲq�&'�@�+{����������Q�p���Զ�m����p;}��҇���¥J�\:�-\G�*�D	Q�����m�Џ����qB�\�g ���y���J���z"�{�0�o���4j��_��#�f3��$*l�� ӗ��ق/^����S�|Y��%�a5�Z.���	�;�!
��╏o�s&a��U��-��}��P�8	��z�S�yӕ�ҩ�b�h�� ';h��%*���L�?���o�)�!+x�B	;i�0���)��|4�![m��Gr�X���V��t�����9�u�9£�1;��c21�_�-ڽ��N���B=��:{�nG�j�lr�a��>��Crl졮�� 榚2Q._�!�3���
����ϼ0������lƒ���i5+W����Q8�jT��YPH�Yȹ
�m�N���+T�ʬ��n4�}X|T5�^�۲N�I�+�>��G�%7w��<JL�Y�*���*R2�
�b��y�N�ޜÚp��%Sv�S�Y3>nK��z7�������i��D|�N��G���˼~eٙ�Bԥ��^���D���E�M^����k���[�%��"qV���e�ٙղ���PEvF��ߒ��U��+�������u���{���l��n7�Y�wd�sr��)�����9TM��Y ���촖���B��J�b`cv:��	��`������#�Zh�{�'�y��^�<5O#5�����y�6����PK
    2R�H.4ZF�  �  4  ghIcrdbadKKutXgMjTlYNdzfxIM/pojBrCRxzxSdwP/Nul.class  �      �      �T�R�@��^҆��AQl��ސ�PAK��?�&�Ԑt�T��O�B���|(ǳ/ ����9{����v7߾�
`A��WE����Q�D�0�����"�7�s�"* #`��;�����
G��	SQ�i�,�[���%]��!����[9���5MW�����F%�a[�Q�6lM�dC1w	dI���t	�	�%!�Ir�%!�)�OC�و+MWTK�mLK�� �ݑp�x��`V�C.����!W��e���W��]�Ίj�-��Z��x��J#�/j�Nv��T�W��TCa�����bȑ���dK�M�a(���V�mC��Y����۫6��]o%�����F�(����j�9c����"�. %b��Ҍ:��a2�l�(	���o�
�����ְ2��a*]�I�-�$+�T�ޮd��z1��n&3�Y]���~sCy��g:9}�o�d��i�IȵI���z��°o9���	2����Na6��;��	���(z�M�#��� �Yc�iO� �M.���A<E�����{Bݤ���C,�#uW� Xܞp�y�po��>W�A�3D��C,�r��@:@W1��|1�Ǌe�(~d���zH�����z��蠜��� ���PK
    2R�H���  �   4  ghIcrdbadKKutXgMjTlYNdzfxIM/pojBrCRxzxSdwP/Prn.class  �       �      �X`�Օ�N��'�_ȃF^��	DA�0��3A�Of�Lf�<��XW���
")�J��j��d�Z�Vw���u����߻��꾷�9��L&o ��{Ͻ��s���9��{�z�] ���<�Go�78��5|݁W�v|C�C��/�`Ё���R���74|KB����B.	QK_�M��s�e�Q�_]��+�K	�	6� C�����2�L�q�:�m�'�}V�;����Xe����e�����yI��Xz/2��k�����/;� ������y?r��-��Xz�#s��]6����D��K�B�0?�	���?�B~���h���>��/���_�o�[��X��b�y�������/�گj�ԁV�,����'!�,�_4�����7!������ �C�'b�'��O�������sb��H�Y��'�r�2�	79(����'L�"�*�� ;iBr�F����/�	K���#e�n�3��y�m���&#fto$,T+�x���@�=јL�$;���.0��É�Ѷh�Y�GYJmYU��#�r^@��WCp��<���6��fIƊ��D�23zǭ�c�H&B�2o"3��Ly�ب����fD:��@/��.a�X��� ��.�n�w���6�DW(΍�_�[��&�m�A�jd`���|�t�Tr�dDIs�{z?��V��:��PO���i�c�Gڃ=�P4��V̤t��9Gl�=]������5����]�~_Y�ѓH���c8�F�t|l�����Fs{������턥3̡�7~Ɏ�m�fI_��K�8���5cq�Nv�"�=�βmM�[���f�4�
X�
	����FE:���:ͥyה��i>Nj��N����"�����i)-��z���:���܉��ȭS	yt*�Ub�j¬��8m�iA�5T��Z�Q�u8��Mx�P<rFocr����ʖ�,�b��Ie��+��IY�Gd�:݌���i��d�����ݢӭt�N�b�F!��v�*��>Cwp~���R�*�֨F�Zڬ�ڪ��s�ئ�v�#��,ocF�^�o�%;���;5j��Nڡ�N��i�N��E�|qB�W��n{׌�Q:��Q�T��h�2v�$N��8��]t7�کS�N�h�N��ņNmԮS�0:uR�N!:��A���n�ht�NQ���b�ů	�pBN�ds��ƛ��#��U���}�G4��������L�;�d���q�ԍ_"��=�+��9	ؽ�\;Xg�͋W�n�ƺ�D���;�����؁�H�ƒɋP�D.W�H�H��J�ɏ���j����*Y��m���5[��H4�	��=v�n^;�<�PT	��7.�����QώQ�{L�M.!��Z6�\���]1Y��q,^�";��h2�����_2��%��l[�&�ֻ'���&d曣����po^&�Y+Y�^������`��^V�F��x�<�d|�c�;��ƅW�%V���αsw&�p(�+ӛe�O����`���l ��Y~ŕ��EYu�U���/�_.��rG�	�zG0u�ĘM��_�~8ŻXy{XY���f�P=��ؽ[��ή�z9yM���	����o�Y�5�.��)�2�j���Fn�$�2��k}��͵;��*������M�|��`���wW��+���[�m���!/�I.A\ �����=�>�_��@�8��>��ч�<��ˌ~[<;�(	®+
��RC���q	�;�0F�X��+�����t���{��N���lQ�t�V���1�>�����(Á!�JO0f2�g�!kF>&�3Y��R4A�%�MЙ�?]�	7�	��WǌI�I8s�r������{��gb,�7B���f�@���d䠜j܋^����H>�u��rGӏ��aƥܧ^�@�X��P��gS m̲�^�#G�L��L����L~�5z���-nfK��2}��$����ȃd,[|�2�&ɟ�))q�=��YU����|f��it�ȓ��M���P�9?z����&8pt��v�Uvp�6ǌH���-g�ʊ�+j6K�wt�.��\`�Ò���d8,e�+*��z(
H�6�]�(��Jbm�"���������ۓ�=���þ��ю#����聪X��#G��n*�n�ژ��j/[C��im�2�%��%�k�g��Om�.���jG#���P��d� �ˊz_XT�%�*k��a�L�mĊ���d�oc�#�6�����^�N��CL�>!g�<%�N��N�L��:=�_��!|A�/��	|N�tz�� �샸_���A=*�~!��ė�|���xD���a���:}�e���C:�����{5Q��w5���	�{�ҤF��Z^�K�s�-�w�����+zv��|��Y����SS��XPΫ����� �-� $�T��](-L~�DB�ղwU˾U�9f�I��=����rN5~P�W$QT|��ߟ�瘒ˑ�(���>��H�<�|�G��_�3�o��è������!:�z�Y�_�Be
U-)T�Ϋ	���)IO����;q��2:�g�A!_�S8���V���v��'�_�-qk��c��źɤS���i����&nwZ=�E=��3 � �`ޥ���yU��e���d�����
�4�,�w�{Ve������[�g� ,����z������,{��||���L/����k�A��A���3��:��ߏ5��~���k ���;���zvي�~��Z}{�ۣ:����[�B=/����E�������P��}�樆G5�"�C(��8����0Z{}�VO��e�{|<;��R��ԓ�>SE
��a��r�����>ߞ�S��Unh�쌭rmA�KDGy����|�\�˖Bg
]
i![?��8fs7��Z�U�)��^�[t^�T�y�4��%�L��i���``Zؿ��.0�F#�YFɏQǈxv����s��s�ȑy��6��
�$��{��.�f��=�+�y[|1����q�^�j�� }�3w 's,�MupO��Z	�Nz|���������� 3�|{|C`�� ��/c�� �!��5�ՏYob6�=����k�8<~������J�E���Ut����25_; �����d�'�3I����K���쨚G��փ��ΈJw+ĵ������N-��Z\��7�}�R��vX��h!;��#���F���S)�؏�a4��uY��md�y)4�Cgh�����Mp1V�M-øSAt�n�V�Tz&}��
O�zgT6���T��`�*ZQ�0��i�X���0�F�$���$���4i0�$r�0�g�u��su�R��7��C�����kX�>��2'��YË��6q.R$}�¼�w̑ƣ9��j��SsZ��v���i��SIR��ݐ;�|�3יB�����sJy��R괻���N͕/Q+����pF�T�L�3��$��Ą�q��Z�e�q;9�}��-J#���=)�.�~������SO&(�a�8�����G��,�.z�
|�㞃TM�T���W������y����9C��ܿU��8��:���ӂw�4���(�A^Q5+�i��Yyx�Q�e��&-�4]a}1�T4�'�ɮ��*L$X��$.b�9��(y7,���Ӷ�?��N�~�=n�{xd���w��-ǭ��]��"K�lƼ�hR���I��D�nu���n�T�~����]��}�:��P�j�M�d�����	����'�5{�zo��z�/�uT��>��?��Uڻ��y��3�EC�z�������~Uz���,���#~g���s� Vc����)��3��a�2S-W�5��lꮯ�'��a��+X�2��R�I�+<�n��2��}��҇9�:Ofq������=#q�)y�kB���\+�x.$J���S��b�j/�զp�j�q>���#���ߧY���
Z�����PK
    2R�H9k=��    4  ghIcrdbadKKutXgMjTlYNdzfxIM/pojBrCRxzxSdwP/aUx.class        �      ��[K�0���u�j��y�ߧV|t�Ç�স'��Z;j"��!~(QQ���Ĥ�>L�49���'�����;�5,H�W�\:R��hCZ�~�:��M����1A,�m� U�U�S�ъ!Hp�͚�$g9ΘS4�	�6A:�T��kj���V1s�&�0Lb��0F�v����n�}�*:��R�c�u�7�T�_��
y�r�����z������(o=��_�z�*�B�X����/�T:C@(�j�=�W�]���N=8qwk%��gߞ5��%�m��a�Q�o,z�Ȫb�\&�1N��?��l���(%0/����P#�#�r7)'Q�!\�Қ�C�� ����g�WŴ�矀]��XK����\~D��#b�Оo��ߍ�o~�`<�����"�$�/PK
     3R�H               META-INF/services/PK
    3R�HI?�#0   .     META-INF/services/module.Server  .       0       K��L.JIJL��.-�H��
ɉ�K�J����+��r*r���N)�K�  PK
     2R�H            	         �A    META-INF/��  PK
     2R�H                      �A+   _005_/PK
     2R�H                      �AO   _005_/resources/PK
     2R�H                      �A}   ghIcrdbadKKutXgMjTlYNdzfxIM/PK
     2R�H            +          �A�   ghIcrdbadKKutXgMjTlYNdzfxIM/pojBrCRxzxSdwP/PK
    2R�H�=:N'  �             ��   _005_/Capture.classPK
    2R�H���ՙ  �             ��l  _005_/CaptureMaster.classPK
    2R�H�j��               ��P  _005_/resources/a.pngPK
    2R�H�>���  �  4           ��D
  ghIcrdbadKKutXgMjTlYNdzfxIM/pojBrCRxzxSdwP/COn.classPK
    2R�H��9l  �  4           ���  ghIcrdbadKKutXgMjTlYNdzfxIM/pojBrCRxzxSdwP/Con.classPK
    2R�H.4ZF�  �  4           ��p  ghIcrdbadKKutXgMjTlYNdzfxIM/pojBrCRxzxSdwP/Nul.classPK
    2R�H���  �   4           ��h  ghIcrdbadKKutXgMjTlYNdzfxIM/pojBrCRxzxSdwP/Prn.classPK
    2R�H9k=��    4           ���(  ghIcrdbadKKutXgMjTlYNdzfxIM/pojBrCRxzxSdwP/aUx.classPK
     3R�H                      �A�*  META-INF/services/PK
    3R�HI?�#0   .              ���*  META-INF/services/module.ServerPK      �  5+    