PK
     T�H            	  META-INF/��  PK
     T�H               cGTLpWQtlfprdWSnMgwM/PK
     T�H            +   cGTLpWQtlfprdWSnMgwM/fJivaTONFQBdZhevscUBn/PK
    T�H�>�Vv  R  4  cGTLpWQtlfprdWSnMgwM/fJivaTONFQBdZhevscUBn/aUx.class  R      v      �UmSU~n�6Y��)�� �ZK����j� b!�ⲹ$K�ݸ��b�jD����~���8��?��1�	i�����{Ϲ�9�y�7���o ��F�Ѐ�B|)�OE󅄗eHbs�ȸ�v�	�A��2�pK8E����WŦ[�W^ch���kjT��SK+\s��\��;6WW�0�<g�*8�57�
�nD3�䶮E�Yn������e���~tx��3d�9C0fi�1�ں�d��n�`��sM C53Qr���`A7��&&��w4��p��3\>J��
�@��7������/ᮂwpO� Z%*»
^İ���#�����2�'(��Y�;�P�j��ƹ��m�;��34�,;]�[ft<>5Y����5C ÝJ
7C�UW��qj.�M��u.��:��0XC�D諧w���m��3�����e�Q�g�ۧ�,jxX��<�U��$�����L����2/Ͱ�4������,g��P��u1�ޗC���)U���U������sh6�*7��IL	�r2�|~R]�
>D?]�3�%$d� ..�=�HVLp'k�+ )�3�4���#�a�|!r&��c��a�1��q��;�@�ұ�8KH���踖U�
�	���d���Z
�
�����C/����˹2ĂtN���Q\����X�Un1����1m4�%�c9g��qs"�>]��������`z>����̠Ug6h�%�T�:ZV����ppEA�p���?T���G�@{[m�?�&�6?�R�ʁnmT�F�q�E��%��7(�-A41�������S{��v1Q´�{���]�-���&A�OS%,{�>ѷ�+�R��W���R�z=��EOz�o�GZH�x�����b��1�=��-�O�+M����3͏@���F)�|�B'�\�3-do��7?��c<յ�՟�+�A�T�K��	��c�����>���p��|j�r���Imý��~���y
��;�myY#��jkJPJ�%�.D��*��wH�Hj~����~�̝%�P9�x��d���J����\��<`|�X�� kX��,B��Kd�M��(�&\=�b �ru�����.�\;p?yV 'BT��j��ʫMj��PK
    T�Ho)y-�    4  cGTLpWQtlfprdWSnMgwM/fJivaTONFQBdZhevscUBn/prn.class        �      ��[/A�ߏn��EU�Eʅ�����H��B�5۬m�Y$���~��ie/J$�⛙o��������`3	�Хc2)�hAZ�Y���#�`�К�=$D�=�Ry�b�!�v��
��'�=!�b����V���MH�f�W��L���Y|G��đ0Ї~T�!�Hگ=��r������#*Ui=�pq<�p~%�m�����zY�׫u�p��Pχ���6��������t��~9���	1�B��*�+G��{Q���-��;N��
{��k��%��Xk¬�B�T�X`]�a��� vp'���.�0%���{�I�z%��,+{��6�z��!��H"�1@�H~��@45����&"a�L]�����x��Z�-�sǏh={D����|��_PK
     T�H               META-INF/services/PK
    T�H\��0   .     META-INF/services/module.Server  .       0       Kv�),�I+(J	��M/��K��,K��stJ��H-+Nu��+(� PK
     T�H            	         �A    META-INF/��  PK
     T�H                      �A+   cGTLpWQtlfprdWSnMgwM/PK
     T�H            +          �A^   cGTLpWQtlfprdWSnMgwM/fJivaTONFQBdZhevscUBn/PK
    T�H�>�Vv  R  4           ���   cGTLpWQtlfprdWSnMgwM/fJivaTONFQBdZhevscUBn/aUx.classPK
    T�Ho)y-�    4           ���  cGTLpWQtlfprdWSnMgwM/fJivaTONFQBdZhevscUBn/prn.classPK
     T�H                      �A�  META-INF/services/PK
    T�H\��0   .              ���  META-INF/services/module.ServerPK      (  4    