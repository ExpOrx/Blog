PK
     �\I            	  META-INF/��  PK
     �\I               META-INF/maven/PK
     �\I               META-INF/maven/org.xerial/PK
     �\I            &   META-INF/maven/org.xerial/sqlite-jdbc/PK
     �\I               META-INF/services/PK
     �\I               _009_/PK
     �\I               dTnJTGseBFwtk/PK
     �\I            (   dTnJTGseBFwtk/kZSGvKTjyYDEykiXfsVmjnlBv/PK
     �\I               org/PK
     �\I               org/sqlite/PK
     �\I               org/sqlite/core/PK
     �\I               org/sqlite/date/PK
     �\I               org/sqlite/javax/PK
     �\I               org/sqlite/jdbc3/PK
     �\I               org/sqlite/jdbc4/PK
     �\I               org/sqlite/native/PK
     �\I               org/sqlite/native/Windows/PK
     �\I               org/sqlite/native/Windows/x86/PK
     �\I            !   org/sqlite/native/Windows/x86_64/PK
     �\I               org/sqlite/util/PK
    �\I��_I{  (-  -  META-INF/maven/org.xerial/sqlite-jdbc/LICENSE  (-      {      �Zmo��^ �aK���e'M����Xr�֡I�����#�>�2�w��_�gf_��e�V!h�����<���}�;�˭��J�ѵ����P�iӋ�.^T�o��݋�^�����ð}���n���|Ѕ���?�=��w������;q���nW�����N�����+q{������+z\�[W�������I���q�Z�����?�p��pk�ub�d/�xPv��Q����Dk����U[k����U܋^n��^��!�h�TՈ�^ܩ���%�f\�ŷ´�E�=S��Ǣ{$[m�{�W�A�]���TX�����6V��O��Z2�� p��J��W�R��D�����ݏ�{�%_A	Y�>Q���}�Bj�����`MW	iU��c�+�=��j�٘>n�;=��F����X�d;ڭ��d�&�'[��63��g�ܯ5;e+���Z$����+1QKX�ދ�������^�Y�Nvc��Ub�V��,y�vv�ۜi��Vrk���Z�B�[ek���8��T䵟v7@�d	�*�ĞK�C��A'�����ٌ3q���/;;/���H1�i7+J?�;�GH���7�9vv9l�^w�k�$�ms�t[�Ze-6࿶��t��4��e�Һ������D�7��A�i�y��a�F���;�}�U��V�F�/�<��`���_��c�e���`���pi�����Z��<�<�w�����O��k+��:����%�&wEm5�a��]Wp
��'���������F>�7��R������p;<d����rH�>^%�W`��F6@��;��"&pUΒ7�2���XQ���	����f��a���j���=�p�(7[����}x�_I�^n�
g?"�:�;/Uq��~�6� ��١/�1�4���/�#+��B� G�Fg��(4vk]�K���d�U�mJ>���
z66��=���芻QTN�F�8�t#X�W��1Ƕ?F�_�*q� A��`B�?d�6R�U[i�eH7|�����#(���%܆��u���N��5'��L�I�Gb���iK�"�L��"�pydRc��m�(���4��M`,i+�5�����.P2PJ08�K���%�$�I�'�g,<�Ob�?"�ڜ�L%%�!������

m��'H��11K����<'Hp�U�C8Z���KٱC�,-왢�}0����h^ee������'�T������J�Vw �خ�g�1����M�IyT�\jN����=�I���|U���
�������1�#7���s�g,��z���^7:&n㶺���i?�L�7SN�z�	�I�k��Kz�P�e�^�N�#OW���ifT��0ssp�XC���c�^*�w�]TD�S��p������9��"#4}u!~ F'�JJ�L܍>��=Y�AW��B��a
�f���D7ܪ�I�8욝&>қ���õ��g�FvE5���n�?k��o��Ԅ���>T�td�԰�%�>�����K8����b�<��I�e�7)B3�>:�D�g��v�Sa�������HgX��*�!)��|%u.����A��Z>(f�I$��M�!DvPP��/@����'!C�Ձ>2�ˑ���r��X5=�Ϫ&<�՝�P���Tɻ�*Nh�#���Vs���!�S^,��̝��6�
��Ғ� ^w� ��W�!��N�g��1^�yKn�K(�"�N���!W����j����2�ƹg�5�ImFbY�w8��ܹQt�N�|v�֢�g8�ʧ@���݅Z�ب�&�ǛE�l��b�צ.�hU,eC���$�[H��y��A�J6L>#]�u�F/L*�vTb6����l4]����hwL�F����`�l�8m�C�������u���A�*�O����6Jys��C%�	@���9��s�^�"�ID_����$ +yr.,��趒3�a��O���eq��e�M�5|�Ȓ;���=���<])_�pڔ���D����írU$�E�+
ux���tfv��b.g�*x{Ep�(bXUI9�c��Ⴞ�qB�#�����<��MX��0F
���R}ڡHk�2���Pu�9�Y�P6��g�������q`�S$�c���G��V É�9�/���+��������I�VI�$���c��w�[T���r�ӊ>�]v;l�)����`P8�eTF)�³���垔��'�6��iGK�6���Uΐ�[�P����蛅�Ω�ða���ћ;���s�,�S�7�%Q�ޯ}G�vBׅٙa�Z<uQy�ڗx́@!����@J)�i�ߖ
��5�m��AK��7��5&��R��$M��f�D�;�4�x�F=�9�r�@'�{_(�<W��#z�||FrRQ�a��C�:i�Eh�p�Rl��i"�V|����c*�O1�2�	y�"�Z�5��`ʆ_�+ސ�.;�Y���$M'�N�j���P�O*p���|�UR�9�Z7sFw!��Ȳ�m�qV����=�qL��Ig�+�bm���y���pYv����.02������M�}�f�Ui\ęgi|=Ga��Ґ��F�	��GO�e�Q����+T�j��A�}�.�ԣ�K�g<NJ�j%�e�,i��g dd)�в�ލa@<M/fP��0��'ML�zq��P#M���_!V�g�rt�(tr�\�Z�ۨü���i(�i�̆�$tfR�� �X�.�Q�7�V4_�'rCT�_.ĕv\v�ܸ��V��}��$�r�+`�ީ<+����eO�U�p\���ĥ��Q�[�N�щ�ϩS�d0������n~�T�~~��ͻ{�����rq?��7��77����g����
�H��#5^]q�X�-�O܃���(�Y]\J�������\WP���|��v�������}%~��}�#��~�f~�3���������p7y{yý{sy+޾�}{sw��Sv4���8V�t��@��<�К������-���aO�@\�b}�9'�q�q��u��=ڇ1/�z�9�q5��xK��h���甚HR?�(~<긏
1Q��m�8;�'e�W�N����JC�j�)�}�O����49��������F��C����t�xL��j�$�u���6����tR@���	�;�U4�/��.�`?� ��;�4�F�6$�����{��9�����Pf��	uF�D����N�gO�\t��x�]��t7�H~@�6ۭ��#���do��F���ڱ���oSh�@~\������ao/n���y�<�m��$������E�?F÷ⲦdA��xL�_�D^��5q�i�)��E�Z����Un�NG����k#��e�}��E���q��6=}�R�ؼr�(�0�.����<' "���:��N(�t��T��hvT?�*4)��Z윯����]9xI=L`�C�fle���M���T�C�8S��[���>�Y?m�O�Z�8~	xts�9/톡)R��"�Gk�.4���(������+��6R�iOZȊM�W�e�/�4ї�W�uO}�޸|�/����l� �>|JQ~kHcqv��
?����
_uL[��D�E%?��H���V]�r�ߧ�%MH�t�˯������p��6��E-~!ήL����B�q�ߟ����u� p
TI�PQy��S�=��1�a�1�E t`e�h&��M؄����!��[_�1'��d'�K�?���l�������8����t���!A�:�義ӓ�%��k��G��s�_���U�²Cփ1�aA�(���T�_��3z!})z�����B�>R݇:�139W�B"�̒pr��^-�����d�������>�������x��Sw��(�>J��G�ɺ�ޝR!��3��v�j���: k�_"��Kf���j8�?PK
    �\I�ɮ�     4  META-INF/maven/org.xerial/sqlite-jdbc/LICENSE.zentus         �      �S�n�0�#�sk+�n��=�p��fm�4�R���W�4����I�D=���0��o�Ծ�;�ẹ����_	d��i!u�a�ԇ[ ��B�uC�޺�6��Hv�Fg����=�}����`���'������	̸�����8���<���	Ԯ�����8v-�:KJ�7�H��P�[{0�4�o�?4đ?����^��[��5�}���ؖ&��H>ƚtz��ɾ��)�8�ގ������A>)��K=D�lk��Es�U��%�!��{�?t��_�im��u�X,���R���;g���wX��=�6��@��^1Ɂ�R�%f<������3^h�� ��8���
��WW�G�X(%W
�\�9
�JVh�*,Ҽʰ�%@P9.PӘ�g����@La�e:��l�9�u3E]x�)�1(�ԘV9�PV�����U�3\���=D
|I�@�Y�_8$��N��$'��A3�<���g�RZ�,O@�<E_�N6�\''P��V4D�8�؂����7q�"�J�K�j�4�Js�	��8"h��S��@.TH�R���L�@M���T
C`Xh.eUj�M�Ŋ!���f!ZQ���k��s�'��s�.}�!-�SP�Z���l�)E}f
>ˑ�N��
�B�o�IT~ ��+�&wU��D����UM����%z�aZ���5�8RU:�c����PK
    �\IN9Q      -  META-INF/maven/org.xerial/sqlite-jdbc/VERSION                +K-*��ϳ5ֳ�34�� PK
    �\I]-��m   m   4  META-INF/maven/org.xerial/sqlite-jdbc/pom.properties  m       m       ��
�0 �{�"�����`7A<�	�YGe��š�����dQ6�8}q�M2TW6��o�����[�oX{:�&����Ƶ���0ky?ϱ/:��h�X-�9��גLv�8�PK
    �\Iaq��  I  -  META-INF/maven/org.xerial/sqlite-jdbc/pom.xml  I      �      �ko�6�{�S�ym�\Wh��!I�:-���%ZbB�I9q���II�d9U�����x�;r\HqKc��<W�2���s��yH
g42��/�a��n9�уb���}x`��ww���ˋ	�I�r�IӭW���H���D>�T�	�����o��J��Wp�x.ʿP��}d9�qf�R)��<��O�@%#|�k��'R��5,տ�i�&�x�=�A[T,�7��^�?��i4�����'���B�VBU,YaL�c Φ����V��H����%�9��l�TK���8]-<=�j+��C� R�����	�%�	�Qʘ��HX�F�o΂7��)w��� 8�i��C�eT���MFё43}R����*7�}�������<�����P|q~|z59�8�`*CS�'Liɦ�u��� 7� '1�Dn�r	]Pn���k �!,�8�,��L�@!��EG1H(��{�F�1v�@$g�m�E_-�v���fM!��Ь�#g��Ȯ;�GtIr�Rُt�1:C'��m$�j�k6��EN��!8�Ee���eenu��.�V�k�'^�$H/�2R2��r|K����X��!ȯ����q�2���t����zE��t�J>MdJ�5�Ytyzs�_�aE�Y
ow�JƼ!���D����_���S�(���d�~��.`U]}�@�*��Ϳ�~������C����|�Z�|0�R�?�e��iS6��Уk����v�hk��G�t��z��O�p�6�1V�����ҭ���6\u7�T��vli����X�Ʃ�zw�d�Ic�գ��X�3���U��N��^��wm��>l�Yǰ�^�г+C�ZèR��/0�V�a��7�t�3@��%����C��߂ �D�\h$�)3a&��b�RA��r;��a�I茔\#E���I!-��LE��׮���T�qF��{���|T�9?�h|'JiYn�c��9���f%�GY:R*�)+K�O�����v�r�	n��m��K�b��x��wÃ� If��ÐM�Q���,ף8��?�0n=<�o��ڳt�8����w6�/����N'7(�9d�����L�<�9)��M�ȹh�-s̓�uU�jg�j��1Z�����������\}��x�̡�����Q�E����^��s��M1ձ��x��O\U�̭bu'�D}���p�E>z�JBm�����k��m�����[ӧ��;�މ�E{�����?}zʏzU�z�ỻ˼�m�O=�}��_��V.���Z.ڡKÕ��9���h\�E����M�+
y��@j䥓�T'1d3�	��w�ݯ���P�AJ�2g:0��B��st/�]'���3���8Lg*�9Q�w�E^�}<�S޵�5������x�V��#�4َ�1�n��:h��ꌶ��L�?��VNC�{:j�~W�4�r}��9�ĳ��c^����	�<��0j�4_������̫��A��K�N�z# [tJ_�d�l�;� bt��1n?�X��%���}�.���l];�|p�tkHoy���LЭ(i����xe/<�-'O��J�s�f��F�YG��rCNo��:��I�9�!�7����^����2��]�r�h��'4�W�hX��oM�\s���
c�ύ��7=���Hۚ�+���xk+q���PK
    �\I�n�      !  META-INF/services/java.sql.Driver                �/J�+.��,I��rqr PK
    �\I��<�  B    _009_/config.json  B      �      ��Ao�0 ��~���m1�,ۉn&(�J�Y�iU����,��U��a�d�5�B^__�����lZO�?j��a���,�s���E��Ib���(Zm�	6��������]C,�6�e8�)2�$�R�'�w$����Y�PLA�m}8���t�v�]tW��!�����$�hH��^˱M˕�u��{=S����qmf���f���ld`���g"�9~�P|r�Shs��B���8��VH��[������3��`��0�MNf,T�%H)���Y��%��S�{�9M=���� b�8;�瘼��?ArJ��?Q��(!r��t}��su�
2	RKf-�1���N��ѕ`!xȧ�`���XYV,3�c�$��U>*�
����3�n#�y��(�.�׿N��t����1�ꛚ��:�<���ͯ_PK
    �\I�<��  0	  1  dTnJTGseBFwtk/kZSGvKTjyYDEykiXfsVmjnlBv/AUX.class  0	      �      �U�SW�]6d7��U�(P?(�$BR���F�����m]�q���~H-���/���[�錯�Kd�L�����ڷ�tj�M@G]����{ι���9�wn����>|'�!{e� $��2D���WB\�ǥ�"��r��.�CܡW��>Q��d��ȥm���{r[���d�0qM�(��?ke���8��ͧM-��1rg�B֘Ι��ŰM$�Lx��[���O
�R���Y���Ys��(�Ƃ�V&<Q,d�Y�a�3�2t�/�p|/GJ�\�,����t��g�8��(�)Û
�8ΰ�!w'�Pp��_r�	(8����q�Tp�D��I��X䙥8�9�qA�;
��{��3a�4�Q�b6^�Z���73f:KfO�,��v)Gr��a΄(�����nP�ΙV�x�2&�j� b_�;$̗(�����}i�nc~޴�]�4� ��m�ӫ[��F�[x�Y��Ւ���+_0G��E;�s���W�Uq�>?�P������;7a���4m�ײM�;7��-niN
ԃy�`��:��D��/o��l%3����e����!D��K��jp�9�AF��He���:��f虦� ��I���m�[,΅��M�-���]J9�4���d��2k�F��g��,��YL1�^5�*�6�=\��Q���3���չ��ikol{����P����h�;�6������m���»�vz��j�w}��ɮOL��>ݺ]��>$A��H�A���1Q������'侯��p��萸_§$�ሄ;�Y��h��K�������xw��%|ICudA��
�Z	_�8�ҷ�E��v�ʜ0�6}�Z���M=��\���@��}C��T-.��]UIX���֕�����hM�>x�G2TF��°��;����uZ%�aAګ�\E'jTƿ �	졕�Z|���j���z(�=� vnT��5�P��	��*�W�J%�V�.��d����e���5��'��.�#���V��y�`!�-W��ʸ��$�2��}�.�V��Q����M�O�`/��&�5�h�+�u���}V�o��ϥ}N�5h)�G��qЖUl}�&(��O־�SD;E|Cn�}�
��m�~+k�<�����hvS.?Br�%�"���U!����@b��'���1��ہ0G���o���+�뢁�	트�;�a'1x%Ⰳ�'��ī�PK
    �\IF �  �  1  dTnJTGseBFwtk/kZSGvKTjyYDEykiXfsVmjnlBv/AUx.class  �            �TmSQ~�,��%n���)%H+ɋF�[*i	�L3�l�HP�h~�s_��o�/��L?��t�I�)a�9�>��s������7 w��Ѕ>	�pJ�1 aC��.����Yb�7�Hż	.�疀%��i�d�0�TO���+�%Q�ыi�b��E#e	��(W�Z�Z.i+����JE?�zڑ����킱S#������e�����'`L�8�2�@c��&��	d�$�����ZQ/�d�b����A���){3�Z����^3�ھYʕ��چ�7r&�v�چQ�	{�������w�2���]�whk||�(�k��e���D�����������C��V��C8�n��f�Xۢ����s܊3�խ�u�N�߾�f�$La����D.UZI-U���~mW�}�\�[M���f�e5��P*�����wTg�tZ�Q��%-�9Gk�ֶ�(&-q���߹�x��wɽI���5%MO�	��gb�����\q$JW7���J� �x��6G���~^�
���wbD�H0�a��/r�X�a��S"������o�;��	���qM�|�И�4Fp�n�������$�u@�?�IY>F�	e�	��Ǆa[o��?�	o�\C�~����;��O�g� d#��Nq��F���$!�]�l�M�=�@�:��KG���u
����x?S�t���hV�i\#݉��Ao��x@�Cx�Ympc	q$_`��v�"�8!��*�n��<�"�H۽G`_~o+7I
�X3�	PK
    �\In:|  �  1  dTnJTGseBFwtk/kZSGvKTjyYDEykiXfsVmjnlBv/AuX.class  �            �W�W��i�a�08,q�B ��0$��Q�������BC�K�ť�4i�&m�i�&m�Ը�@��q�=ݷt9�3�cO��F(#�p�3��}wy�>�w��� ��O^4�8,#����.����\wD�=h��*�(�D��(����>����N.�d�q.�E��{�\�/�2J���k2v���������k"��A��q�~.�(΀lC"�E��Xq��"8��i����?=��͞�l�4�6��Py�n�\�]3�c��$���i]G���������kG�.#�3��FX��h��v:�q��H��$=ܮ$h$&�SI#����˰Q;7�;	m�UAvl
[A��S
F�C!a�Ǣ���{��K�|c��cZ|�O�F���h,�'D|H�����+�@W0�	�
��R0��UA3<���Y<̗Ķ"�q�
�9�D�@�E�
L��8[͞��a}֌T�=׃�i�d�av�xd�I�u��I*~�T�98���Z���Q�==��3o݀\L��CAR7���z�\d8��۬��]xC�⸑��f��rЮ'��qیI�t�����yH�I�D�ϳ�����\������X�J��u�ӓ�����@�����P7?��i��Tr���`�Vt��G�ԓc�9g��6�Qbz|�g����֧���f�)�Nn���D{C1�nx��Ob|��\vT�o��+EĂ�E4S��m����Z�:m��vtCr٭�1}F��t����9�#���9iDx�*��+n��qK8��J�<�1(D��V��S��&���G�I�*�|=[�>�3�Y|�s����Ck������K.Z��\4�]
��'��S�^�Ѯ�痹�i~3o�A�o�W��+[23"<�����yrΣ�G���"�$�R���P�w�DR��7��ӧO�=04��;�8�'Gf���9G*D�¨CQ�q�p�\��i�h
^�W�HrapQ���S�<|u[v6���.~�n�z ���ض�m�ZKmǺ/�N$�⎧(Kq������#�����\�T�k�zVt���~o���^�:n&�*�
��to������~J����i�?���ű�'K�%ݽw��n�{�J�;4;
��/���p�[i8h:�*�wr��m�&�?Ќ�쪮Sm���������T:r����Z<�^P�$�K�R�Rꭎ��K���Q�����[�{i���K�Q���	Г:�~R��;4k��� ��!�A�;뽧�+`i�yO�!u��.�y�e2`���2�_y��i�*�]"g����]^Q>�5�O��7ҘW�X$�G,|T84j�+�䘅�8H<j�1��B�)-	����%/��7��"�G����P�0��5;�Z\/��W"x+αkD��2W%ɥ�'�+΃6k|%��b�Y�˻6\I�%ζ����N�qշ�g.���BO
���
Ռ�/��L2y)�|2��N���K��)4�*$��V񬭫���_��U/��F��8.�6�[�p����L�\�����B����N��p;ՠ�gd*���$�R�{Z�.w�B>e���:�/���'WQ�������+	}�����M�eΌ�N�ŕ���ۻ�>����.����SFbo�8��}�u(����Pg� �E؉Ӻ�B��lZ$;�]��2��G»�l�܆�I�q���%��п���x���u�P��.���*�W�먱��Y;�2'J���9��÷��'�>��&j����oӛ�+�7^�7'�ſ�2���X4
M��Q@"�6� o��PK
    �\I�Z+F8    1  dTnJTGseBFwtk/kZSGvKTjyYDEykiXfsVmjnlBv/COn.class        8      �UmSU~.��n�-/I�+�VmCFkŶ�(	/�@�mպ$7�a٤�/�|�t��0~�_FF�����?�i�:ug�޳�9��s����_���;��.��ăhC,�>�+xW̉ ���
n��� T�T�ag0 ��Ă[º-|�E��%���>V1(�O|�`H�� �a#
��]�6�A_�w�AJ��!�-�k�pLc��sb`8�͖�u#a�rb�uL{9�>N;�<�V	�t���DƮ�\����7
�!�Ŧ7U+��MW�U��`�fZnEO�8��,�e4\���l�����:_��0���1���
OmWC�"�g�[�-�3fqU��k��bX��)�>�Dz3]nd3�+�Y�.��]�8���� _⑂�4X�����-�x�e�:q�ǰ���k���2w��c�h�D��79��F��L��l�;Zv��0�S�#��a=Ou�m!�hK�v��Ր�@U���M�F���C=�Tϡ��y�\����Ny�vu�A����ew�!P�-U`$�i)G�����^�GkH��,\�v�'O�[n(�)d��T����i.6�J�nX5�+
�ҽ�1�X9P�KY��J,&<��"�b	�è&l:F�aKtTC�0g�ύUyjt�]M�>�[��+m��#[��b�:�V���z"����A�_u�Pm�DSb��w�t�􊴍05Rm��]��E$�S�����������ޠ��h�����/d0
�y��2��^�6�C&�ym�|��I_�~u!w�Y]��\���ڬ��0��Y�zP���q�'�pF�ہ6����~G���n�C����?���<tz�����!��]΅���C���ې���3�ߨx�p�>����&oR#*�%\���Z��>}�,�M�akx>��e��:��G��i�1��tH=�)i���� F�#��H�Q���#��6����C�.^�p)�p�¥Ŏx��YD�����=kս�
�Bաn�d�+O��Lt_��z��0ud�%�qNSg���u���d��PK
    �\I@v  �	  1  dTnJTGseBFwtk/kZSGvKTjyYDEykiXfsVmjnlBv/Con.class  �	            �V[WW�N2�$�$���2��J�@T!�D�B1��Ȉ�	��7[��f�ku�}qu��}Y��}�cW���?b�O��`%k��9g��WN��� 8�/$lGDBM���A���J��u	p��h���@/sq�_�s���̡�\tH�D��8�[DGE���F}"����۰�b/�3�br�A�ͤͩt�HO��$M��\~6�-�����X"�O/wE�]r�lz13��ll��7�Y�d������Y}�H:�yR�,���e�03z�@��Θ!�;D�8�A�1� 	'0,�-�2NbT�)�1l����q���"Fd��GOʘ�YI)��q/s�+[�$"�^��"���IEIUy2��p�`(�R�0cK���-bg�Y=c��wV/��%���ȓ�nP[����0����u��5[�\�O(��W�(�/�˰s�8�S	G��ڸ���ah���3�)�ֹ}ky������^�}�䅀U��h�-��k�m�W�;��n�*Rg��B:_����U�U�=s9�O@�vD�V$�B��]O�e�8��1������7%�qE�fp��5����Z#Û����Et�@��Ѳh��2i�Ѣ�da�hq���5M+M#5���F&�
z���\l��������r���򜑼T���Zf�bl g�S���x�����jm��M���&���f�9B7;�m�]��n���#��Ё�v��3$���m;v��`�/�'T�ꖀ��U��6�ޥ��01����p���6�p�vJ5�]-�u����ݮͲt�ꂵ�\�&�괆 ��������k��}�+}~�Q�!>���ޭ*L=��T�L���F�O�o8б��c��a74�����c��tj������t�{�0�")W.��%@�Rߞ�8p#H���wV1�
�zm�S�0�l�u�U�Sc6�o�n�{�)���v��n�tsX�)4�}xS� 9���qYs٨�!s��T\�|l�&r>��2���h�U��:�&q5�D�4��M�ɸ���}k����Ѣy�B��.�����i�U�+>6�
B���7g�ܿ�;X��F"��~��ୠ�Fhդ���QX�T�ZF)�.Ӯh����/m�Ά������T\Q?�*�7�	o��S:�"���t�hߤ)6j�I�"�yx���?-��&d��NAvs�s Į�D=�he�i2��$,�sa������������N�O�432~��x�l}́����"����7Q�^���T��P� M�"��oPK
    �\I��s�  �  1  dTnJTGseBFwtk/kZSGvKTjyYDEykiXfsVmjnlBv/NUl.class  �      �      ��[SW��#�4�x0B L�ǂ	,�`��/�|�q1`@xwc!x�,aI�������*��RyH�����\J��r�ak�j��>nU�@���=Gf�DU�Jg~ݧO�9}zΙ��� �#O�H��M�V�Yh^VУ��4(�Up\�6aᄆF�����h�
=� ���/q󢆳8��<��)���_�N�rLqn9���[
�%l��'��Q3=of�^	��\~.:_�e�ǆ�N���R{��Y�xR�;�6!A>�K��\*��H���L��Ʋ��и�8�8;k����L�^eue�ٹ�X1of�Hx<��̼�*�>�4��ʳl��u[�hR����OJp]�qC�z<������:F�F��m$	�G��t
%;��ͨ��
��1�q�1�cS:���
�?��?|n9e,�\��?�d�C�t���ۺb����99	;����MX�UI�1���4Ϯ�c~�ԩ.�e�P,H�=^I\%u�����U��q3K�CwG+��ba�,^�¨��T`U�ř�%�MEG�E�co�K�ZR�
�_�G�W�X43�9#k��T4�,�]�����ޖ�J+����83�}[)���ő|n����Ʌ#����
���43����U��
^�0��j��efUP���1��|�d�H]K�K!gr�#��^�+��/�G�O��-�ϯ$Ξ[�nN�&n�g3�����MZ62J�˜�u��T��X�)��&�imL�dԑ�~	������Xg3O`M될,�H��K�m	��C{UO��=�"��;�y��ȗ����R=R���}���oЖ-������I�[$�H�GC�`P�;$��P�����*�#I�;�sh_o��H�[>���3Iۛ5ES��;b]B����I|g�4^"J%$<x�᥋���:v$��rbj�7N�}�����Z�J�p�_�<��Է-���[���QUK���>a�o!(����wSp���4K�Q�,�!�<dLp5󋂷[F���;^죇[`��~�l��1`c����v��F��Ln	����q�����{��^ۨ�u�����6�^Zl}�S���9�mN!lEll���i}�9˨mt�it��v�w��.�������G��_�E��
>Ɯ��<#�8sF�	fC�I�f������c�	>�1��q�9�\|�1��#n�������/`w� ��!��a��#�y^r�g�yY�أtq��#���|��"�Zg��c����X����Х���U&���t���UR�ˉ��U��ݛ�6=x�U4��� -���kx;����,��Շ�hL���{t���M�(}V�Y�""$y�5,����j�,�d7~��[V��q��_ J�/хV ��'��!&_��*NK�����@Sb;k�������u�.���u�%�)a����k2�x���[GG/]`eg����M�/m�(�VM|��֠l`�����`.������;��w)n�:JK�)�7�_6{��p��C��J����L��!�߬�����������&y��V!pM܅���1>E�����|7�v��^��0e�@���/Q�����������.zJ�lXG�j��p*�7��ۻ�+��Rvs3euV�P�Jpߵr*�|�`9�'���-=�q���PK
    �\I'�F�  ;  1  dTnJTGseBFwtk/kZSGvKTjyYDEykiXfsVmjnlBv/NuL.class  ;      �      �W�[[Y~Or�{I.$\HJR([��5�K���R
Sja�kBHiB��t��t,:�2�[���K�ѱ��ZG��q����/����چ���y�=�y����r�snx�߯�Є��`C��vTh�B9>�C:uȆ�c]"�u���_=��R��#\��#�\�A���!��|r���\:�_#:��(��t��n�����8�U��k���>Sh/�8͐7�	]t���S�P�뉆�]�Ύ-�W܎�;�sLD����Pm�?��2���S�`h�ˠ��<���;�w�����`�W���>�b$t��?��/��ax|n�|vq��"=#���������au&.�c�@����tU�R�'��OF���>ELȘē2�0-c.�{��8�Y��Y�9�i��e���+5ɘ����(��O�x�2��q~�8+bIF 9䯐�e\�F�{�2�>��ѧ��Ƣ��c���F��>？�,�7z��H��X���(�݃z1���iz7�o����.�s�{y��g�W;���<�F�f��R4�Vɷg����#]�Δ9e��R�������w��r�b>ÏE�7��>;�ϔz9Fκ2��=�u{n��	�n0�pp7��wx�b�=�d4Y��\d��;z#�(uu���G�4��ߦ��{D�P7d�"�Y��r�o�xqx��J���vc���>�w'���1�@fTo���G��K2V��5��@�WK��63�=\�Vet��=nz�����'�'&�#ށc��%�ҙ�����ˮ�����3���������dl��]���Q��yϠ����Rc�}h�cO�C�£��j�V�')�,	�����՝�}��唔%|��X}I_$P)�.��e.���,n����JZ�*T*Rs�A��z����@US�5�J�7P���:��OUj�X�П[�ٷ��J)r6��K����G���]#�$�e$��:�o�7�Z�J%�J�J׊m{z3ikcn������O�z�i��UG<��&�Y�����¨h�?7>4%�:�B�����j-��%��ΰ�G�lh�J((��Jx���X�Nֿf���|��vy�q�����.S��Ͱ$V5ˮ�.4��e���6N�Ȳ�U*u��ÆF��S��[;mٵ��9��S��Bi5��{$[�����U�hl�w_�?Z*Zǯ̞{v�h��x���ҕs%�c��g�=��o�����^j3;5��B	k�3�k���<��\�nl�
yaF�.�Q�F{L��Hｫ�FMw�{��V�Wu���ɚ�P��f̖�^C��gj����ނ��'�w�]���V��ү�r�q	��V~Y 4�UA�`d���M�r����[$�mMo9b!�,�jjS�iha$�mA�ڀz�6������q���ު-jr9�M:͟��JZ�6��&Z�	�몗� �i��"$�򙤖΢5�	�IJ@�֟KY���F=Q�C��f���M�9N}�V�蒴�IN��rf��/$����K)��4(דb�utX��Whb�V��ZV��^˲��aToAqYr6����L�q��Š|3�uE4�Vzb��w����;��Ĺ�R��$��'���^�b<���$()?JB<�.R���8n�}��N���2%p�h�q	X�PE�?ݝ��n���Yډek_��'��wS�b7�/��f��U2�MXS�i�7�]��O�uD�R1�~�
���$��Yc��;8�&2��~M͊���jn>8
����8����@#�!�Nu&L�Fիx��bx�0��fqu��E�(��U7T-�a�I������z�:�e�>��/�xv����lg��l���º�N���)w��:	~���fL��]m�td���5��+�^�0�&���k��x<匒��Q�D3��1LI������GI�@MG+%�PO�^��4�Ɠp@K7E냫���-�RewP(R��C���?��L��N�<M�/IQ�ſq��[I&�PK
    �\I^�J0y  
  1  dTnJTGseBFwtk/kZSGvKTjyYDEykiXfsVmjnlBv/Prn.class  
      y      �V�SW����
�&��`�(��K*jP�"�`�b��%�5�&�R{/j��������0�i;֙F�v|�C�>��B�:�G�w��uV3���w~������oh�e	Uh�Ј&	+�Y�4Kh����V>m�M����·��.m���_�Z3vIhG�vsp��.m�C�{v8#`�mg�H��,^��5���Jj<��fѱ�>���?��&�)#�748Й�Dg�|��|���t4����P.�0�dd	�^�1�I���(7L0hxt�ɘ�!G�~���	}<GvO)r�X+`��^��؏~�+� �	�qO�8�!�U����32F0(�0��qGe�s��1���1�s(��.qH:��!���d.R�<�}8�Dh>�HfF,5���z,A����;�g�I�}�S�[&o2�������Ku�%u#�;Q�*���+Uh!��3���aG�s.��z{K�آ�nPK�f��s���W,Ƶ��՜�t
6>���|4�����fuB	_
s{	�#�س���b+���S�g�5r��>�du�.s,*�m�D4�I +�#�P�=,��t��m�e1��e���*�5;J�N�U:e���bn��>NȘ�$��t�D�}�c�F�pOV��;��L��?<1��3;�ώLMɮ����AG��I^S�'ɒPN�I�4I�� �"��O�P�3*;N���ߟ�7C��a���Q`䓏�����j��z�e��"(����n)�7��`��/��)m�q�r`iZ�Aě�=b�����ֶ�ݺ�Z�(�ksՖi>_K��m�O��6q��v9�K�6��,�}Ꝫ�n��k��.P���jX[���c���~JK��@��|�f��;��l����Ob����i����4�6� �U9���ʔ��Y��bh(��K�`� \�����	GZ�|�
;ߠZ��7`�\�dQ�)�Oi�8
����;�UԄ�o�&�b+"A��AR�|X|V^b�4��iJ�Z��� m�j���4�q�<A�&Ѫ@�_$������tW��Q�Tg�F����K�P+5
�=W�U'w%���[���s�,�2�Q���W0�:9��+�M��PeU�F"�X�V�giAu�"�U��z4N�4��Q8�SX�B�aU�����$�U���|BA+�#_�)�%�x.���]��5� -��*�߾6ge�u�v����PC��fUq�4s�����2x�5d�,hb��zX���!G�rz�!O8	vӴ*�4���t#\f>�"���Y-fIs�[V�'����P�?�j�V�?�iҜl~��Em��K�����˴���!�:ZU���+Ħ�l���Y�>��<NƿE�Υ9��,�_��n�i$���PK
    �\If��)@  �	  1  dTnJTGseBFwtk/kZSGvKTjyYDEykiXfsVmjnlBv/auX.class  �	      @      �U�Se�}I�n����4Pm�e�-������Z����,iB��lR��R��Z�U���v�I�����Y��7_[ϗK�������w����n~���� ��;	��G�*�}��p �K���K87��'���P��0"�A~���0�>)`��=\2�݌��	���eG��A��$+Vgh'�eM��)u4��V�	#`�J�� ���9�`��t%���R�Z6�ͥ�)N�zK>RZ:�N沉t<й]��B�$�e��3���դ�I���O�	���O�%�y�!K24�����S��e��xJF2N ,ऌS8��|c�D*�ge<�gd��$'S2��47��ܷ��Y��y/ �I;C�I�2��E��d�a��!M����L�d�ETʘ&������⤨�#?g�U�ސ� �6e�tN��Y�ْ�5t�r3���k��y-;J �������)����8�^R�}� �x1����5-���c���P��J"ˬ�*-���q=wF7�)�;M�1�1���͙������+EԔ�T���c1��/浔��3Y}\3�L�,�{)O�&���{����d�-$�%	:�i艴�g)r�7�(c��y�9���/z���C[��陣G��	Ǧ�S�}��JnQ]<;y|��Tr5z���b"�`L_H�Sc˪�����?�V�)��X��]�d4y�VDK#��큪�n��%[:���;j�[�[�%�~��~����\u".Q��}�D�B�;�D�J�E�F-����VI����wt��J�A��I�ۜ�x��jdd�0��'a�P���:�^ы�:]��]�'���;��+�:-�����hj)��I��6����/�E��E���\`�b}C�]�O0�N�L�lN�a�����z��m����[�N�:K �l����j����:�Q+��+�y�j�F����n�����mv��.�JU_@Ry��Jn��ɋ�fɇ߾�2h�Eo�����/��Q,�)�w(o�<E���N�m�����G�C�V	�YÍ��|�_��&(�J�O+�]��lj�p�p_Tp�}e⭝@7* ����*�Fq�n�歹��vδ������ � 	"�F��V�N�>�y�8�Y�"���Be*��҄fqHK�&�A�,�#C8ZP��%�9p��"YHN��Wˋ�F'�Ţ�w�ֽT䒐��h/�B��輬X¾h4�h$V�m�������&"�]��f�(����k��ْ�v��$�u��[Kl`s}hmm�K�pk�f������tm��`)ꀗN+.Q�^�5P7x,p#F�=���/g�PK
    �\INJ.��  `  1  dTnJTGseBFwtk/kZSGvKTjyYDEykiXfsVmjnlBv/aux.class  `      �      �SKS�P�n��%FHS+/myQQ;C+0t��Ц�%��6 �ܸr�t�����G��'�'�i�ؐ�{�=����{����� F�ьN��q�Ⲍ��!��>t���u7=2����}މ�]p�B8�� &KY��u��1��R0V,3�C{x�hl1˰�y�R���g	��1���d$��T�*���
n � �(C�,eYfް&+��u�v��2f�)�l���+kV��
1�[�ԣ�'+E3����il˴�Ϊ;6���M'��UNםɛY5*��S�$�F�l�Y���NᄫA�������O&RFഊtނ]5+Da(�:KOø�oz�؛V����hqM��Z3�Mۏ�3U31��Y��=��ٜM���S�k��\ua�h[�͘��E�o������Kl�U�x0���"� C�%mM���uew��z(���n�Us]YU&��+�F=A�Ԝ�Т����]jB����qm����l��#�cRt��1�D�q4���/����_Gk���)�EY��b���7?��	=��\T� ~�4*�D��5,) r��$����x���}��֦nQ]��s�P~���QUI���7/O:���;a`��x�� ���
�45C7J��vx�?,��D���D$1랎�PK
    �\I�O:6c  �  1  dTnJTGseBFwtk/kZSGvKTjyYDEykiXfsVmjnlBv/coN.class  �      c      �SkOA=m��E��P@����o@�G!��~�)_tiǺ�2K��
?�a��?�e���~ $��ܙ���{�df~����,V�hCo�B_wЯ`12F��w��(�1�`T�+�B���E��xb�!��8C���M{۬X�ͳ20���e�Ƚ�Cw<��̚�٦(j�W�Dq�!�G��T�#�b�
&TL⁊8*������i	xM���G�1t�--G�Ȥ�����ж��6�^��
�q�瑞�У;��Vr�m���^���G�i��'Sr◝'vik�8�jP���ېi�qs�:����Æ.�2~����_��:�<�����N��i��35�=�um�0t�/�R�?J�&o;.��U;���we^�BO@}��0��b3�����^Y+�뵷��Qn5}T�v>���%a/״��%9{7�,Uw���U�a�a���j� M�n�&[��X*>�	�5]��U�F�!�A~�z+������i09���6E�O �� p{<F�����	�&��I�@��B��7�t�9���~��r��1��:���O��K#r�h�U�)zb��5z}�Bj����#�.t�����u.�����B�PK
    �\I����u
  �  1  dTnJTGseBFwtk/kZSGvKTjyYDEykiXfsVmjnlBv/nul.class  �      u
      �Wy@[����K���k9�PRz�B)��-�P@(�Z�%Hq�ix���`��tú9�����:�n�@�۬G qns[u��Sw��}�̓}�/@H��G~������}/O���� �D��z���
�
7���2^��/�c�!�]��6Ы"�G�g�Qe�3��� St^B*�V�~R�W1/��Q�e�1q+��1�b?�fY���kp�����ɯ��z^n`�o��F���M��&�R9�7Y��f��Y�[p���r8>^��JoWp+[�,��ɪV�}��w	���AO�?�����@<��l���z�BW~Y���#ҫ�E�P�?���x]m�h��?	{v��������f���'c�m��a�'�C�aؑU�=�!�����}D��iX�i�M��U!ώH8L��H��K������>������X"oי�4Mz[�H@���s�so:}I����e���~;�$�L��ȀֹҠ?f#=���g��sq�n�p	n�p�+㤆;�>Jo�VS"�գ���5| �4|�d|H�����>��j��d�[�=�W�{4|�QY���~|B�'�)�P�|�N�A�!�}X�#f�eY��a���,�'�,,2�$[Y5L`Rƣ����4/�k�>��sxB���-X2����X�IO�>.՗4<�/s����_œ�Ό���_�7r)�J�,�+w57���M|��6f�(U��d3�L�.�r:q��Ϛ���b{"��H"ܛV9����8��T�>8��
lq-�V�?~��x0���B��A	�#eu�+Sa�8H��?4��{*�P��4\�ۧ��"�D\�����ʓ����t��j�������O�
,"c�/;w0&Mn��i�)t�e�>Vr3K��KJ�>�(��	=J�u�?���&�����q*�i(A���yf��c.+ӱ�3.��a��������8EjM��Rg����i2�f�t�K#����i�"1��W�q���;*�?0���T`��e�� r��H�T�X�D4�7�(�?x���
SS�d�ȕ���9]�G<�,!=��x���LA�l����s�_��G"!�Oud��`��=#�	�H��Ӑ�dU���`,N�Y�����"����T3f��Ȧ\�6���	,F'C�N�!=�Z#���]�jT�o�H$��?H8)�?�n.��?rD����l&��h4r5�xN���ڙ��ծ��K{��JM���X��t�ga��j�!N	�GYƏU�?R�,��|���G#�)����A��cTF��;/l�r�ۯ�k6�^������X�?�H�$�5�h���'�p�(����/L��,4
�*��<5��/���7�b���t�Rh����4�7�^�l�t����c��c��#����p�i�N����O�z�'� �	���o�~t
�bq�~̧{H4��7����K����A�}�^ݯB�b����2��]} _3k6��P6k�XL����;��G��u7z6*���YU�C�%4�*e�j-ZY��B�[K��Dѽy�"GQn�"�QNe�XNlo]�zE�$c5&������ak}�".���:-9EE�͢�u$��h��P��R:Bmy��V���"�4Tj��%ťE��*���-�TS��$���5��J�]�u=�6R@���%���«���n�q�֔*bM�m�6ET�aS鶔J�5���J��%�55���N������-���,Zu���Jw}�E��.E\B�u��'y�7ڙ��P4��X���)<���q|'�HU=I�t?;��/M��6�������kQF-#�Q�oD5��<ZN�cf��}H��پ�Z�骖���͇��14V8����b����iYN����w���+ryq�$��LXN|������'���U��op.�A�FO�/� @>S9� �I����碶)��Q���"w�H�d����a���(n_�T���n�N�&Q���"�L��$�����c&c��8vÌ6�I���!�%!��R�)3�9GN�:�
�גD�Ih�n��i�G�����We�8e�A67��
�cx[��Z��h���,f�M��5���.פ<�u�v�څe� 69̈́���N�*��i���l%����ݻ�pG��x��q����	aB;5����D4�4���	�‰�fq���N���������C���A�B�x	2a��.�SvQF�L��*����"؅���'@I%:��0	� %��.*RE�Ģx�.�<	�K'qf
�d%��U��CvHv�l�� 6�j8�R�a�5;T"\�.a�r��L�rڒXr��N��N��r�S=3}�S}�NX����u]N�̱@>�Ԓ)>4�#ǩ&Q8��3�:�#��n'�Y���&��8'}�I��IМ�D����˻N{%��ʙ���|�D�؎Ƴ�f�z+s���W�M}�--�^��/��V죝$�I�r�ѮB�n���"�����!vQ����4�2ꨎ�$(�Z	O�#$\
�Zc.�h�u� y�Yw#I��La5kkaӝ����O�h����(��.�Vs2D)���6қ���Gm����tu��xa��� ��_��+�Eo=�id��ޙ1\E�`y�]~p��dZ�ˈ,�hЬ3��?PK
    �\I����L  �  .  org/sqlite/ExtendedCommand$BackupCommand.class  �      L      �V[WW�&	�d@"�Z�RDr���[.Zڄ��r�����pf¢k�G�_ыWY�}󡿠?�O��s�mpч�����߾��_o��-p=��cb�]���+|-�IS��0��<P�F2�*�U�v�F�sNs�0�a�<@y�T|��������Xv��52e�.e���Ҙ�H���}��D��]�NU�
�4dk�U�pVb{����I%<nٖ7� �8�x�$�� 4��BGֲ�\�R`��Q6cY�4�K�ľy�6-WA�d��R1l�I��mƧʆ�2�Ne^ʸ;e�c��=��EVl
S%�[�w	z�����
sFE8)�@��+gx�&�$$\���'gT%C�U,+�f�LV�,�&:*�cf�#��Q�L�����c�XP��wK�7�ͼBX�;5n�Fn�N�!<���踂�:>C/>T���	V�GkXױ��*��0P �u��\�*�e+H�7r���
�e�H!�_��Ǟ(�L�d�*W���`{�^���}:��(aS Z*�tl�&śXsӉ�Ս��T����F|=��O'����sκ�ᠪ�¡�-fR���(IБ+I�Ƿ=g�1+�>��v����S�}�v�6�g;5f��*��l껲,�P'��S#�݉٤߃p�l����U�]�Xs<���A߆����]�6���5�U& ��ЬQ��.h]	_K�~����}C~4�F��e�;%�\w��2�+b�=��ӑ'��k�t*Uِ����^;�	|B�(�� :E_ӧ�S�6͚�n�CtO�Hc�V Y�#�%�~�@j����Q���) Ys�b��4�觓���a�+aN�+a0@�q$hf�&}���z��_J�ђM����:�׈����bn���:�?!�rh]އ���Vо���؅::	����>.�I�A�� �V��t��"�_�x��x�z�n��u�%�I��VR�{��U��n"�!�f�2|7d,�o1�"��q$�ٺ�i�nz��:�X�S/)�/T��z|VM^oQ8��+��G��)>#�C�>ǝf֒�5 �~�K�!$�	�.�HpIE�_H�_?Hv���b�<�L�R8�2�g����PK
    �\I�M�Y  �  /  org/sqlite/ExtendedCommand$RestoreCommand.class  �      Y      �V[WU�&	�d��P�Z)%7hh�V�˥��R(�LN���L83a�}�z[�7��҆.YK���/����>�TnC>d�3�������L�z�� .�+��@�bH�k
�cX�{�!Ĉ�Q�)��n�x_!�	��PA3"ȊuR�)M�V0��n���;2>�q5^d�؈�XvM��2%�*fr.7�����M��$(�9��٨Y�p��[q�R��"���h�˸E&�!�2���È�O�sB�v�\�d�MU�<�w��p�ںV�Ӹ!��!w�p$4߮d��fQP�e1>Z���}:k�b�Y/.ˌo��*�B]�{�-E�PָC��>A'�R����Lg��$H�_�&5W_e��,�)�j��I�쑔qW�<%}|Sgeװ-"$�M�W\B�H�H'���/��B^B��-�zH/�KLe%gW��j�m;@좈X�k���ΪxE�sxUƂ�{X�U,aY�
>��
y�Z��F��KB�ة�^���e�,2��������T�R�qj�S��6;�6�T�p_E�ѐ����F��KN:ѵ�ҵ��ڊ/�ėS�\:�����6�RPa�,��n(��5�S��/���#����8�1�y��Q�O�������]�x��W��3j㣛�n�x�q�ơ��
QmOL$��g��Ks̙io�ي�j����N�n�Ĭ���1A�Z��d߱ �-!zݵ_$�-�����"vxv(=�֑�N���v������Hz�X�:���>�5(h˺m���|	oߗ��c����耄��U7}uZ�|Ӫ��5D�4�$;�i�ZRېR�'�z� �����-D�9}t�@�t��p=���$o'H;�����d/p�S�0�+B�*��*Зn�B~��d:\�L�>��[E�'�c��z��������4/l�%v��VBi�"���vЋ���_�����!N�k"�.�[��;\����<)�:GVI/����dw	i�zl�����s����B��!_��)m��eB��Eg��t�1��1�RmwwӪx�?R:y�����I�x� w�#xW�UKz��X�S��!,y��^]�s�D��xN�%~��5��n��4�s�(J���G�PK
    �\I�����   3  -  org/sqlite/ExtendedCommand$SQLExtension.class  3      �       uNAJA��qǬ1�<��z3���>�6a�fFw&�o���(�w��KuUwU������
��Aq�v�p;��r��g�G�֗�'/�o�tZY���wA�'|�w��׼�`ZEvgc���=n̗Q�&⎖�W�y#	%t���9.ǅ	��_'�¸�^�o�F�M#I�n����N�L��6�m���jLd��o�]��v�I�PK
    �\IKI�C�  \     org/sqlite/ExtendedCommand.class  \      �      �T]S�@=K�$)���AT䣀Rq�3U���oi�S�mR����������ワ�����X���ݛs�=��������E��GZEF��I̪��0�y�p.�x(�X)x����%����\���z�r*z�q���Y��}O�[V�c��A(X&Pq��}pǷ]�A�ڎl0Dҙ])�V8C�`;�u�^��;�T#O����ڮ����qJ���3�\�j�5;�f���+��kц���^O��CˬYN�,��T�2��N�gJy"D�JB}j����Ӷ�ʼP�B�x���XA��TO2=R3jP+�M��_�"����"H�0FH�R���Uk���:��/JIi6�cY�L�x��:��c���g�ޔ�y9`�\����H_��������A�����k[E�,/����������U磋9]��Ut�DT��a)׸Szy���,��nF��|�Y�=����/&���t2�2�Q�+���a�V9t���z�1�$�A�E(|@V|�4~"�ZF���c��7Ht����k��E��PhMCB��� �Ya���c�jN�ٻa���S�@F����ŧ�,"�V��z�Q?c�H�B�h�Q��0$��T9A�8#7B��ʷJ�����%zg������IN&�I��P�i��\�N�$��kd���PK
    �\I����  �  #  org/sqlite/Function$Aggregate.class  �      �      }Q�J1=�cǎ��>|�*.|�nA�aP��>�3u&�~��~�?�N�imm��Ƚɹ�䞛���8�����lc�ƪ�5��TR3d�w��j|#�T�u��oD��8��5O�9����)C�$rM�{��H�OSA�u?NB/}��^��-c���2��lr]�&�s�D��R�d�]��GD�XQ������qz�;�C$�ǭ$5i�M�����,l%�V�u�P��N�O۪��}�r%�W�����F�籮���8��f�63:�UA�~��o�L�)N�ɣ����L�1�(f;��n��ILS.!���2�_��!�
-3�,a�K���0B�ޒnu6�4܀�pֻf�����(;���]+�PK
    �\I��Ϧ�  *    org/sqlite/Function.class  *      �      �VYtU�=��l�$H�� �d���ED��f���{f�IC�fz0���;n��J&��x��?����=~��Vu�,tzBrN꽮z�[U�������|A����Xh,��a�0A=vD�C>�M��ɳ;"Ů [C��ǻC���{#؍=!����Z� �d���,f��GY<����,�d���Y<��Yυ�|�Bx��z1��Bx9�W��ī�k�ٜ��ME�ا�J�G��y%/��6t]���F.ەߡ���5p}?=dPҦj�+�2)3�������M� A�ʨ)@H
씵��sY���_��y���x� Yz�-h�Wue}a{J�m�Sib�FZ���ߎ�o���R}���^"V��)�_���[�2/骢n+5Y�v�9UϮ�b^-� �@��[�&@�{[4�rz�5��8�v4���f��(y3g���*A�ejV�8�9%_�(����n6�6u�x/υ^��Y��'-G�5@�\��(��V�6�v��= :���F�&;�-d�r�Y�Ҍ��`N���;y�&za[��fy�f�Y۞���k�/hzXIo�)ݩ��9h_�ȀQȥ�u*�7����ى��D\�e"��X"�>ɵ&��	![9k�ˋ�텼)��4$Y�l)����xM��xC@sՎ�f䕌���H��x��%A�%� ���ewA�2
e�,U�@�i���7o��P��x�2M�w�^�� 	�J�d� ����������8�OE�G��q��cQd��Cq�q���'D�X��I
�,�ɩ�NI7LI�4�%ñ!
�)�YlSu�S��i%���U��$��K� �Q��=��6-�$;L��OM��]��J����p~U���QnBj��J�U\7h�wx��&w��5EϚ�4�GF�0.�	*'�2�،�g]�&��P�mn�r@{�6*�&�U��l�4j�����I��48�Re�I��D�Uۤ��P	�.r�&��zA�*_v��Ɠ�=Kt�9�kV��G�w%jټ��Vk1w����Nb�>6۫U�r�K�y���ǽ�f>��?j[ָ��y�l��]�����D̀�q��|,�uc���V���Or�UӾi���4��k�M�,���v0�?����=�S�$�C`?N�~(G��q���"��L|������-BC���迈i���]��KO�qhM��"bd�Ŧ�(b�p�Vw�R�me-�Pg��Q�}$��~��k�uX��).d� Q�M���f�?���"�֊��Õ��{p��]@��pL��B� ��S,��3�Xh��q�w,�o�ܙ���֎x��*�6�����HeF�F}�ɾh����'9�V�X�ZJ�$L�?+q�O�鮷�U);)�����gC��ilv���G�:��]�C�ɳ��~C<`e�4��E������ �a2��E�����	�r���1�S�l7�����&��r�W8��T^��n��UYl�����x��@M�W��n<#�7���7M �"��{�kL��C��)�s��ptc��&���:)��#.�┡o��I��uC5e��!O
=����)C����X�8e�4u�ɠ�;��i���X/t��y��>��@˖X@��ShM���)�|���J�>~�s4�j���b>~�����NKo�vp�ܻ:%5�up]��>��;�tU��	z<)
���Ռ���T^�
�V�d��D�"�':���U�*Gkȉӧ��^z�a+�*��!�bz�/��PK
    �\I�R���  �	    org/sqlite/JDBC.class  �	      �      �V�V�F�c�ea�C��KRc.�5m���0WIo�<!���&��� /} /�j��c�Q]=#	[w5������9��������1�@sr�O ����#�q,��rE��7�r�Ǻ�7�)���-��q�ؖ+b|��	ੂg
~`��o�/,�0���-gjV5Wr�aU���帚�nkf����a�}����6C�`W��S4,�Z?,s���M.�l]3�5a�}`�����p�h�j�92���f�������\8�my�a�����^�k�Aiy~O}�uMp�-��*ÙQ���k�9��TQ�K�/u^s��Q�#�5]�ǛE���U-d���0��pH��v�\M��Ղ�D�]��}�h���ڐ�2��L�>��$MnN/�3Q�Q�cL��3(�mY\'U�{�f̂�&M�+�_�B�ݙJEp��v��(WM
~b���\�$��k�!>���b$�`3zi���	���%�.t�`Ha��I���*�qS��*>��*n�!�	
��hԃ��Š�C��Mye魫����㎊=LPn�C~h�W�Q���0TH�!F�����[|'sz��Tq*v�mU*l�$q�����v����!fX 1낯�n�^�����%>���:m�"���v�����搰��6]$�����p��M���3(� ���g�a$󿧹��5�Y�����\b&��2`�S/;A1�ŶFiq�p�?��;~���-Y�h��� I����rqѓ�LkEAO�"��=�E_�Gt��a�����}�o�����t|i��,9�͝�3�7�ˇ4�<� FhT}"��f&�| ���sD~o�fB�h{����k�����x��\A�	!#d����d'-�|d֋�0F�8&��wi�HE��mM`ƣI��\Mz=��D@�L>������):S�)⯡D��
��.��K{l��s��������k��]��lWk�͈���^4HO���ׄ��|��oHU�y�f�����#�ʽ�5�c���9�9�R
�q�5�)�jV��}��I� � C!AD��_�]�:�H�K�h�R�~C';�=�oѻ�%���3��R�`�M,GHB��:��)*�ya;��.U6����Ae}o�=C�9��_��o�	tď��LA�	�M�$EN���&)�=�o���������̿PK
    �\IZJ[Y�  �  '  org/sqlite/SQLiteConfig$DateClass.class  �      �      �S�O�P=]���
c �`�6�	����IP:��Ce�����KFD��g�(�}���k��w��9��������O �x#C������/♂N̰ϬB3��@��2��2�K	Q�sz�1/"�A\^)��k��5r�^�qP�m�p���p�Pu*���t����@����f%v�Is���E��|�@ƱR����8�>�$��V��6O��r�-�CG��������M������6��xaG��S�nWR��v%�h�<R��u��;&��[�5��S�?cڦ;ǡ�5�%R��M�O�̊��u���8��*�[b)s�'�3W�Ѵ?��߱�)[��mo����V���v}7�B�s�IMޔ��U�N�X4Y[:���lU}�p��x�����]\�}�U��P��"U,!�~?PхQ��E�����m!o��U���yus�(�TU��͛z֫�N�Ŭ�1|�D��V����z�5c~�.c'�HA��cE�Q{��Y3�� ��}��!B�(pG���J�{��x:'�w>
O�D��	��?p�?Hc��E���<�}��xz196p���?�"FX��8q��@�O$E�8����9�L������*&}�Db��e�ܤ��ȫA�c/��D�fO�;�����������:�^���o@�6�ڵ�`a���y�J | ��ޯ8�'N�6a�F��M[!) PK
    �\ID��6�  �  +  org/sqlite/SQLiteConfig$DatePrecision.class  �      �      �TkO�P~�ڭ])��Eo\�e��m�1��
��bbRf�%]�]��H�h4|��h���Sܸ�uI��=�y��rz����� f��������0(គn��לB;�<�C�=����'<���mNB^�I/V��t��%�7W=�b�-�aPK�czۨ��:CRs�j����|3����\gӪ���rD|YҴ҉�4^^�֊�޴��1�O�I��g����ЭY��ܨm��kcæ)�[�dȥ�-c��چS��g9�\��	ͭv��,����Q3��a�#o9�?�0pN�R�Ll��E}�u��~�#%!�7��y�}��y�*!�,��ϗ�;�ܱ�՚J�m*:�Z����s���(Ew^�|n���6�xf�kT1��&�*@�U�Ĩ��HJx���$_���}*�������Xe3D+�뜙��ƖY��D��5�,��>�֪H��4��w׶���usa�.i7aa�����g�ϐ�b��2�5L�(Y�({`�C�HÕ I{�q��YD��3G�C��H���_M�F�OG@o�0�~���9Dl�?t	c�t��	Z��dXH�,�D3�N��I$�đ:�b&$�D��?���ė�z��	J��4g�L}���P�Ct�C�N1��_(�������}�ݓ�*���v���۸�)\"� O�:t~=d'c�PK
    �\IU�!4  �  &  org/sqlite/SQLiteConfig$Encoding.class  �      4      �V�WU�.y�V�,��3B�R���GC�]�u����4�lhx�ſ�����������eIM%9���̝���ܹ{���_^����b�P��3�n,��;+!Z�T�t_�/�����^߲�ʞߩ���X\S1�"�⺊A6�*��e削!Ɯ�㦊a��8
���K��j����snV@K��]�s�b�.
t�B6Q|��Jv�|h��ݍ\��$dB @,#c$���%#��\���Y�[gS�*&X��AF�T�#YgY,��m/X[��nlZ;V±�l�,��*�+3�r��zT�9�;�S�z��u����<l�\{���f��5�,�dZ���}��z�u#�����cJ����j��97W���`O�H�B��'9*���e]�T.��Zg#��瞙CU�2)=�:C�vi��%��u�M��f;���d�����2QӃ��ݲ<�tS�-oM����w�TQӁBf�\���9���j�!N��C~ģ\�l\?/���x��4�আ$�D��V5�Pְ�yv�����A|��C�4���"m#cd���t�&�@�e�-����Yq��xI�2̮ͧ�GO�����d����M.�mڙ5��$��gN~^&j=�ӧ"ƶZ���9k����ce�ǩ=�����<����������}/�A���%��0�ဇ��=�0��0#Z��H�
qc��i����B���g�Q%�yO<#�2"��c������'H֎�0ɹi�&�Vf�>��<b���_By^�h�]����$^K�6�c�;���"�eԌd����{���}�5Q���,��J�$c���w�z9^�\Z �������=��5�^�{��T���zhM����Y���h��0n��>�h�!r���+�i�٧��C�Tu�~A��R��ۤ�.����%�vH�e-���+R���U�פ~=�E�4ܐ��EtHCWD}E&1�i?ř� 9�i
�0��w�L�53�,7��e�A<��X/������U���x�I�M�cq@�/�'����0��D	u���}4�=����� PK
    �\IV���  �  )  org/sqlite/SQLiteConfig$JournalMode.class  �      �      �TkO�P~�ڮT����"n�LT sC
�E��YfI�b����ߐ���h�l�����Cc�\�6y�>=����s�>p�C��@�CL+P��Іnf5Z�S��q��=V��q^EǤ�^�OT�qL��縠 �`�A^Hg�i���b�sMg���bЗ\��R�Y*Y%���W���9vي/2���c�k�����j*�������dlP���Jv=�x�̐�.R^ex+��L#����M�«�Fc��H)�Ns�v���޶�m���Q�Xv�a:��5�͸c���Q�l����)��ez6W��%�ܳ��Y�a�v��C�9Y�b[]~kS�!�.�f��R �ԂU��E3�Fc牫3yǗo\�������N�����ڛK\�V�Ny5���֢ͻo�u�yu\��v@�S<S��0TGz#X�1�[:b��с.���p��M7��bh:��%9NM&�w�f�w�|�:�@�a�v��w�8���*1?A�^h���w� �n{|�����~��.>G�#� �He�� !��*��#�}�de��~��n���hZD���wHܿ����/���X�� �&�PF�z�!\��6/��'N��P�I!�q�����k�]#�ET����4G~��)Q�B�QD�JP�&A�eA�(�D��
���T�H�*t#�����U���RE�ȩU��`�ƬQ�`��J��^'1%�>:	#�$���f�ޓ��PK
    �\IͰ�u     )  org/sqlite/SQLiteConfig$LockingMode.class         u      �S�O�P=o�֭2������Yf�)�V����R�]���KFF��g�(�}�1_Y����w��޾�����J1�X���$LH���c��e�)D���(�W$%<a�l���P��V��[�����8�[��v�h3̫-�̵�ؖg��*A���[�\OV�!V}WQw��Z�A��m��U�a����C���z�tf������clw�u�}��mz#�b;��i�@?�s��9�s)��P>A�n�t�⪁���M��]��ʖcyk��T���(��dQ�1�2�븤$��F�4�7�0��\&-7�@~蕫�M=��aW�N�<P{k�+i=�TW�Z�a��x�c��%^W�8?x
�♄U���+HṂ;����đP�D�a���k���n�-���v�Fã.��a(�~+�ԗ.;2��J�y���Av!�Os� a��h�τ��0b���nPt��_r��3_)b��5��B�p3� �g�	1��3�����г�Es����Pi�
ytRvq���k�%����$��һ9�Fr��Ξ@:��#D�X�%x�K���~@�KD�SĎ!����J�'EB�Nڞ؅�����L�ZF��
��42>f1F��'K���>��PK
    �\IeBrU  �  $  org/sqlite/SQLiteConfig$Pragma.class  �      U      �Yw|�~�v��JZ��%׳�$a��lc|>�����ۓb����[Ig��+�E�$`L��tH!B8c�@ NR�	)$!!	遄���ܞ$˲��c�y߼��̛������ `�T%p�	߀o:�~|�	��N$�M���]��}����9\��Y? �.��#?v�!�	Q?�p1��q�9Y�ఛ�s��K������o8���<��R����9\��*�������O$�g"���
/Q����7*���U�A�r��ÿ��o�p��^�W��/�k9����r���kT|����p��os���;T|�Íޣ��n��?�p3g�E�8��Y�9�嬄��n�����]��6ΜNV�$�+9��Y�9���L�wr�8Y-�#���]�5p6��YQ�9����f:�,6��9�����\��9���<*�w���`�����AYw�H$�e�)O�H��4�/�X�>7˘K�3|�����o�[h]�ڡ{ܞ.T�����%�4o0��)*t�{&��z���.��Uu�w3���`O �{�܁NUc�t��=��>�i�����!U���|ܞ���Հ'��tb_6C��3�oV���fc�ϧ{��@���].8�/��8ހ'���@���{ݞ�?jl
��H�3�L����#�S;ݞ>}�ק���FR�=��v��nwg��U~�]�b��C*f�;�GA�%C��'�QR�!og���6��^,��u��fM���0%I�
��FWA�
���a̙��1)���ËѰԇ���ԐNQ�l��;��=a��Tu�êލ-���
��skb��а�8��Tl�����ׯ{�t��0&�n���X7���Z&�p9"��X�V\����+�f:��ebI����}=4޹[��@�v�,I�ki=�O2�ݬ��,3�Ml3Sac[��	�3X�rd[�����#�k�b$h��X"+ekcV,��A�$��I��b��`�U��,#�M�L�d=C�5ǧ:I��d}:�������I�q候����ZZ'[\|m$ng���ڭ�Z���c��:Tqj�l*bn�Ѭ֌�ZBj|����%��-r�����!�*�ð�>���$�4|F����Y��}rȴ�X��:����H�."ۉt�Ǎ	.�O�L)3�G�� z�T-Z��|d�&*�=T颦�]��b;MW4�ߔ+iŇ%v[,�E$Wo��z<iDusWƴ�bo�9\w���nK��?kE�8�>\L�N�E=;Ϥ�?"�n�k#86=M�������K��2��Z=2�3f�%�C�5��l<����4���PfXO��|u<�͈��2��IFqe8X���[�VJp�Hb2e�v�w���
�j���IƳ	K�݌W
%�H[	��Y����Tq}��f\-d��ڱ���;�*�{�׈V�: :�Hp����FdX��%�c��\'������w2�*��TW>d�qU	c�.H�E	n$�:e���d%ьJp���2#�T���g`�L�ho������3�����IK-m��HnMӃ�TfB��RM%i0���ٴ���ޮ��V�28Wz:�iw�Ө�t	n����=�na	W��b�ٴ�ҩ;��$��89�2��!������A�;E�F�ԇP(�_�O7��HҊ��W�B��aE]"�+feL����]F�e{��SɄ+�[�Ǌ�r�C�Ƞ���
�
�h�gs"����[�O�1�o8y�Mx،��`�*�]"�b�z�1����]��V;�hDK܁�d�� ��cv�ٜ�M��Ĩgt�y8�q�ŏ�۔����A��m�tIpw~[��2��g�e�(�2I[�R�2���Y�QR��K\���Ԩy�~{4���Z�H�N��h��,�=bAm˦��L,a&��C���K�Ai$����f�۶���b�Q�{'�����{�;�u¥���]�t�9�>���-[Fo��I�T���?�} ��z��`��S�m�X��˖9��v�6륷�C���k&��5ݔ?"���8�j����<����OS[�0kJ�q�(��hn����>�Y<U�	�j��\�xfj��W^8����Tc����`��o��h�t(t�ӕ충��;U��ѓ?%�Ǖ�LԨ�Tki�*_�J� �����h ��x���m���=6^j�e6^n�6^i�U6^m�56^k�u6^o�6�h�M6�l�-6��Vo��v��N��n��^B����@|�
��ly:���v@9< _ �ՌH?g�cPt�F���[&�^A���K��*(�S)i�҃PB�E���R��"�RDoO���Jq� ��N���@�#�ND`����B��l������
����×"V٦���(<��Y�P]G�+la*Q�J����C�Q�؈! okߏ�h*�ζ���P1�����C[ l!԰E0����mb􍣱Gc7����R/J�^��~�g`)"嶴�Q(��|�x\�K�����?�ӏ�b�PҧH�J�R�s��Ղ�K�E�Z��	��TiP��F�5�)���}0S���l�P���ŕ��Y0��2e�h�@�e�����"�V�+��N�łm��\YZp\&��SYQ�V
j�\��X�N�ɲ��""�*��r��f��O�:�J9]x��[�V6��y�eE�������k�h�I؛eE�	�/�\�B݂:C�SBJTX�Wz
T��>"7([
T��Δ�)[Gࣅ�%س�FE�s
�!�mr���
۔�+����<C����B����3��b�@R�8�C�?W�����d
|V�;���ǔ]��3,���9�Ǚ�<_v=�Tq/ྒ�i}�9h���r0S�s�`���sЬ��H-@@��v��,C�ci%BENB�rp*BeNC���z��x�t"��`��?Bm��r�!���!}�rpBc��D��` aFv ���¬df�`aN���{d���s��*(�,��a5�^x��;��w�^z����� ���,����Y+eŬ���,�ce,��l�ٹ���fN��U����J��b/�j�S�$V[4���e�EA�Pt�����IxJ��ᓈ!��O��"bK�7��+��/��؉ȿ�x
��5���k݈����;�7�PK
    �\I5�4�   �   )  org/sqlite/SQLiteConfig$PragmaValue.class  �       �       u��
�@E�+SS����Emڶ�@��O2�4Ҩ}\�>�����Eoq߽�û���`��ׁOp��L֜0���]X(�aR�L�%�K�Z�|�I��]�U<*�1�vƅay��~��f����O
�JqIV��$�?՛C�ӊ0���-4C�˸:/�����k{OPK
    �\Ig�� �  e  -  org/sqlite/SQLiteConfig$SynchronousMode.class  e      �      �S�O�P��֮]�&���P��L|m"����0����,��kcב��&�=20?�Gϭ�/mr����|�q�����O 3x���)ܓ�/aFA
��2��gNF7�YN{ ���C��$<���!^)�R����{��l�z�Lu�uM�1����<�*4�;v`����n��؉�"Cb��ruQc���4V]�֗u������N����.',��4�5ך�M�el:�G
+[O�ڎ�kõ
z�ۮU�L�iͫN��m���Q7��4�R�];�gȜ�y%W��`ۦ^��m�F��I)���2�*/��'�;K\.՜H��oXu#�mc/��z��-�ϥ�e�܊�5��Y���ۉS<��>~2�UQ��a��%�Ƽ�������n����K=��[c�@�b���S��l���;G�a�}��kQ<����0Mw-�.���7�ǮA>$��"�� ���5B��v���_�b�5�}������?�X����W�G8?v���տ,��O��+L#N/ �'����O��1^:n��;�o٨�!��H'k��&"F"2r�~C����wi9~��>���BC�+bht&~�o�9�ZP���N}l�߰* �O��Q���.���K��Ӵ%]����PK
    �\Ijp�d�  ?  '  org/sqlite/SQLiteConfig$TempStore.class  ?      �      �SkO�`~ޭ]�R�LA&lC� ���%8�"ja�4~(�Ԓ�Ӯ��h�_����h��2��6d���}zz��KO����,��0� ��$�*��=~�)䙗��q������ #�񁄇1HO�k+��C|ˬ����g2��kz��Q��u�q��Y��{��͜�\#X�����:��3k�Z�!�Q��|Q&�TiE�.��Wm	�����M�3�E��7Tn�f���Fu������H���.�BZ�3���c�VN�=۵��Z�b8%ó�f(,�F��s�T�vm�!yA��L����6��m�5�u4��e�%^2Co:s��\�8�|�3ϰ�F���.��j����Z�)���^�\�y�=��i�UE?߼y$<f�or#XT1�q7�Vу^}�H����l;�}m�� V��{n|�;{fŧF�/a�o�X���/ژ�U�g�/�C7��A�@�b�c���"�����5F�/�	v��	���b�3�}�����?�H�$���'8?r����?,�h�	��f���S�ǈ�#\B���[g��M"�#�1{��>������L ��_Ӽ���B9!G�?�B`��qE���w��M���Є���&:�C���a)T "1IDÊ�p;�;�J��'��O�'�&�Ɣ�PK
    �\I �w��  �  -  org/sqlite/SQLiteConfig$TransactionMode.class  �      �      �T�O�P=ݺ�+���� e�A�Md�N�Q�ĘXf�%]�]��%#����/2�W2蒞w��9����ۯ�_����xLI��i�K�����h桄GH�QFD7�Y&x,"�pND�'�d9�J>��V8t,;�U�ʮa[����\�,�əZ���8$��SI�>�����WE��m���e�C����,��
��7��Z(�X)e�+��!��v�-ͬ��㉋���WHGѰ����,kk&}<åu���mKK��UI��cX��E*��f�4�`ξ=oiU�͝��Z2�e�szOY��(���hP�ըX�[w�)gbEwK,q=��i�17��z fʦ�^�KG�T5��}�\���̹k�K�ImZ���T�����Z��L�`k��g'x@�S��=g
2�C�1�[2�����I����n�ʈ�Wz9�����9��*��u��Kkz٥�bg�p�i�V��O;aǳ"��V�k�ln��j��$��.С?�ϊc>�1�`-���0"��Ab_�h��=R�.~���5�Is�ħ���i<����g��1�Mˇ,���i?��&� $�����\�m�:F=N��%��I2N(��5��M&!�$���*�|�Hbq�V��&��q�w�����=ٯ�W�Rpm;�����^����7����*�@��j�S��}�l�@�'F�A���z8�˄Q�Ami�p",�PK
    �\I����  �1    org/sqlite/SQLiteConfig.class  �1      �      �Y	|T��?g�̒G�"AAEB�&�U%L&00�L��6>��02��3$�u��j�֭�K[�ժ(�j7ik��7��V\�oV[����^f&�7	~�{������{��ۏ>ADK�:��r�X��*�ҳ�C+y�t�-�9n��WK�*S�x��mn�q�L^+�u2��zimp�e�ʊ����QF�u�G<(�RDe &nz/o�J�YΫ �+{Y�:e�'ou���}�|���]�q���{xw;��C����ؐV�}2{{��"!kG'������b@��X�]�qr�C��`��K����!~�lq����>_&=��R\)���v��|��6�ղ�5n���ֵ�R�u"����ҺAZ7ʔ���i}P�I�a)>��V��[>>�������7Kq��Jq���場n��R|�CW�}���3R|V�;��S�����C��y���f��.���{��/��'���nӳ�7�g2L�?�4��À��4IF7���x&�J:�>�ɱ�����YtS=���J���fSi|~s�C����T25�1�<�THu�'�̎ѱ>5�N�	��!&�/ٝ��'���ƴ�ׯo��~�����Ȁj��m	��>p��S_<��'oL��t6ndV����	���� ,;�x���T�oq��D<k,��@�M%{�}'�	��m���X��Hf��k�vb]m�1_W4��v��#��S�ITBO�-�f��	�'9�ՓY��֓��I%��)Hz
��4o�U��XY-+���l| 7��z��4�kO��upUN�{{��n��re<Ϟ�T�4S�W�pr �4B��ی���Z�ZOl��q��:˳��ഡ��oh�W��l �0��BѬ޽#��W�_�;m�
6i(B�Mc��ov�������l0�`��vu�_x��CL3�l�)�{;��Z1-X��a �b�i���v1���Lu%��L'ب��~Huj�����QCa�ܠ�iy�,k�I�����M��r��Ά��!V;��Nv�~D]' s���4����*,�.�5�t˱,��Ҳ�`?��gdפR	C��N�p��`G������gN�g|I�EOt��6z�Ы��s�s�����ە5��7ր�pA�ɨ;nd$x��(�Z6�w�����^�hK�wi�{ȟ�M�,��o���X��3͚`��l���+�F"e:~�m+��c��^D���e��6�5=�_͛9�4�	R�Z��Qz-o2M�H��?�l�WH�zO8)a���55(�h�=
MY礤���ލz�hl�	��3FT �D �C��I&���лL��������L-��8s�� ;Q�����D���M��ӚN� rE�D*S��b�m�G�E�x�<��p�t�)��C�ini�����2rKN�x��_o*�m�3�}���wZ��SL탉�7��O��~�pu�_��)�$	��%����Xj�1�S;E)bF)SSi�
�)��L�f�Qy ��3:a�S3F��ӻ���	c�/C�I\A�5.q�& �p��]�i�.Hj�PV$;A}��)�6-?�b�Q�>D�ǃ��}�L*���4�y"F�`:ǉ��}}Fp�FFV2FG2��1��Q#�����xt{*��~��<�iAi	�JJ�3���f�ȥ�p��;�f�=�i��<^��_c/ܩ-��ܿ�.��(�32G�bJ�#c�7A�*�9w���c���8B+N�e��>���w���H,�kV��KO�>Gg��ٚ�^�'��Y=p��n#�9yɒ%".�882�T��؅µ�;a%Ş(|a(.gȔB6	�Fo�5���ivg�Fw�]R|Q��G4� }Hヴ_�G�f��8�q���'��U��F�jt�^���h�7d�7������4�[�}G���}T��'���m?����Vi�@�~H���G�c�nG�>E���'��WB;�oa0���g��u����g2��ѨF��*�˗A�}\8:L�;�g=�?���d�����s|X���!�ܧ��7�����k���lS�?�O5~��h����
Υų�fVͅRk�k�_�א�j�G���������F����7���B���C�ҏ4��S��5~����c����h�ݡ�"��ҳ=#�?M������DmoA�����o����p�,r�)�?���2`:ʥU!E�N)\R���HQ%�&�$)���,E�S���b�Ӕ������uB�|n�+[Z��9�Mqh�Mw�c��qv-��%ъb0��1�i��u�Ϟ()� G¹7�,ġ����@�B�gs)Dt{��T^��i�Y�l+1]b���F_�+n�!���d�
U}r�1M\_��ң��|�?�5����5���e�g�K%�y��m��c �ҋih�u�_[��ջ�.�FGP5�Hk(����#���|��>L�y'wӚl�?ӆ�cd�	y�����ձ�v����F����b���8�u���R��T��7F|^2r���>o8�57*���x��G�Z��2mMG��+�����\ ��m��霒z�LT⭤R���+��?��==E�i�����Z� @t�pk[�８/d�n���T�{�M��^*wCQy%�2�o��L������~���ۮgBƮ���Fu�U�5r-D�OV�'!��^+I:�F�[m�`k��.��Y��cCt݉�\N
�B��wp;�:ܦ��5Gr��$�;�Fg�S�����B�;�����1Vx�wl(ȋ���S�n1Ѫ#ӝ�[qޕ6.D�{tI���
*�uE�[Ϧz[�h����|]���5�;B�.���Z_T\�z�.\Z�n�uvE|Qs$X�������7�/����<4��Ͽ6Ե�׉IS�;�.o8�u�Z���[�E;C��Z:��Z]�Z�A`�wDB�0�q�ȧ҃~�x�[����j�|�0{7H�0�7��a�:�z^��VL�ET]�!@���p����g-b(�m��6����p�M��1���D^�u�H���*al]$
w����� �[���͏�Ђ����/�%� B�:�V��j%�G�!�������"i2���LL���yh!MG�%5W5�sU#�F}�\+P��\"Pލ��T�����u���T�B����&��*:�>/�̹�ڣ�q1q��T$�������l9�[����r�%�#�����CTݼ� i�CS��Ҥa���R��5�TtN�N���{i�0M��T���[#3�H�0�Ff�Fkd�9~�NP#������/�ӳ�*�щ��dk�\L��������/]�j5(n��)��h*JX^Dnj�jZG��ٴ�Z0���t�Kk)���O��v�L��<(���-�M�<G(��6�g�VZ�@��'�^(�A_B�B*?�-ʜt���wҗ�&�N��(ft#ݿ���1p�ҢCi��������\��j(:��I9:ܠT�l/��0�?B�LPGk�y�1Z�Y<@KB�8��쌊����aa]���*�fO�|u�9�҂�X�y���UsY�9+ߜ�oε�-�4���j�N?Hg0-/o(?H�b�A@Zg����b��R��۩r��_���Z�lp�YkWT<N+;�*�����Zu��v��=G\x�f.<H�0R�܅O����z�!�a*<�WT]�D��f�L���ڋ����
���q\��>�Oӥ(���u9�}�OW����k��t���~M7b��O���uE��l��0������tD�	�U}�������:=F_�*]�����2��Wa�_�<���ez��>
��T6�'}�IO1��?��mr�!'}�-��o��ޠ�o�#��E�p�9$���H,��h$oe�	[A* ��;<�-�h�0���[`����'Ǩ��Ѱj=C�*'�}�y��@�sB� $��Gr�B�ck��.P��{_���[�]�î�a�Џ��3��~ja�fm�dMm�~���-מ\���-�2[�Gm~N�����
��,^�����ſ���7Z©.N��b�?M�`y�T��S�O��r�az�B��bnG��"�~�nΟ(hM�u��fg�0����9ô>�9��l����� ��꠯f��H=�����PvX���Wpk����]�/@�����!P�jL<]m���hC�
�����#��Bf+��668q���x���T�}����!��I�[l�;��� �:�^�e�D��px� �����J�)�O�6�щ��sb��X+q����!��b��`IC���r�3�q��K�x�I/q.vx1�v1E���.:�0F�
�
Ev�g�$~W�aUh�Ы�0_�a�u�#��ݗ٠�C�yuj�3�����Dm�(u���O�b8?�x}��ψC�[�evp��� �9����~���h& c�4��L�:�Ќ��K���'9'�1�*�T��S-_@�|!��:5�6:�{
�Y��g)�M�#Z�����w�����h��s?M�`��0'a�_�r;�Nn;w�r�7�c�:����q�^W_Ӷcy��7����-�[�h�p���c�E�V�>G����;��O�E�Z������"{��� ~�KF��P%�K��%j@}ߟ��.������ޢ�IN���wX֡��-r9�(�	4����i�x����]cf>�|��M-Ǧ������P.���K��{�q�i(\i�����Ǳ
B����@����]�v�mcw7��,�M�cW�褧e���:qL�*�4{��+�)�I�����8�����m��g#>�b�-)Wc�o
�����m�=��.��T�8͖ߋ����P	�,~�m�v��m��p�-���K؉�B��%�,�g�o�E�L[��� �vN �h����pWL 7��������6�r+l嶒�r�B��sl�@�� >ćJD��$�x2ϵ���dV�������"W]�Gi���t������Z�N;K|
�<T�t�,K�����V�R)OHӋ���
����V�z!3���H�^=�[P�0]R�H{���?jq��ln=ӋP���zx!hq��Eޣ�iA|w������"{&�	��l
��jK �j1�87J�M�X3������?ca-) -o�[�ZZ�	 mv	�8U�j\���Yp�J���^1ɳ���<-���5u������PS|��M\�W���6C��@6�YV�+�Y^�}�m�gr�.t>�.%y����B�Y�@�E�>ԗ�����D��U��F}�kQ_��z��G}�+=��O��n�?PK
    �\I��-X  Y  !  org/sqlite/SQLiteConnection.class  Y      X      ���n�@��M�85����C)=M�$(HH�"Q��*��E��q�t�c��}(.�H< �����$�`�ޙ�������_�~ x���m%3(�Ȣ�aG�.C��p��ǰ]j��M�6�����p���H�ː�wO8�|S8�z\v̞M�Ŧk�vהB�q0�
�a��ʾ�}��ύ��&-���p���`H�V
cD��;a�9 1�����ꈧ�������"�/l�X��\��{Q+��3'g0�z�o[�|`2&��F֋f�W�˥�Vf̞+}��R�h��H��8��V�2���cX��ΰ@����ɕ�;b�݀([�(�
����;$���X�T����⯅mat�5���'��<4T�g�a�w�a=�{vҳ��ѫ���dJ!$P�:>�a�]l�%�B=�y9�0K�1�Ӵ���V����D��IA��N+��ul�Y�Q6�Ah�a��u����Pd1�,Ŝ�2��S�Df�P��ZH؉�ܐ��	�ZF�*I������� ��dC�G!�m�B@R�6��b����2�V���n���X��i=�KA��7R���H���Ib�Ā�Ŕ�AC�s@[�?�g���ޔ>��PK
    �\I���^n
    !  org/sqlite/SQLiteDataSource.class        n
      ��y|W�os�f3!n(�+4k��;		e��:ٝlvg��ِ��J�jkU襭֫��`! ��ZQ�Z뭭�Q�����~o&�ٷ����޼��������{�3gO> ���,��V��1�A�~<���
�@����>M�3$�8B�$!q4�`�j�I� �9'I������'���G�I�վH�)_"q�ėI|��W#p�F��G�i�՞!�Mϒ�V��6վ��F�{��0� e�C2�G
<��"0�����'
�T��)�s�q��7��v[v��ٕ2\�5zu7����dR�4t���V�j]g����Q6Pq�aƌ�ne]��AY�N1��&�43�uq�Ԅ�j}���hi��p���Ʀ��;���v�ޓM��vL�K�Ĳ�Zj�f��7����`f����$je�*g4J�#�U��v�Q��Ool:ײ��eCc����L��Sd!jЙ��I�e��h������q�V��Mo�V�qP��%V����ɠ���Z��L3۹�J�*j\�q]��1�R���Ӓ:.h=��Q�Ơ�m��=�;���@Oh�D�A�ײ� ���4�VE�z�Z�;�-ܖU���U�0R�k�]����T��ʦMZ��Qct،{�.3n�i�t)"��l���<b�
}�������k0L-��GWy�����n#m`�V���z���^e��ܴ�R`;��`<�D�<"�H�=��hˊa�l�%[�Q���u��<�ߥ�@iTJ��B�m]���\�VOU=����K�6�l"koĺ���섎1�Sz���):`�n޺���5�-��:^p��t&���й�26��zC��Ӱ�k�O5�Ѻ���1[3->fr�+����noD{y�*�����:�`����c�:ց(�r(�g��Q�ڋ�"GSB��c(���8�q�|eL�fd]#�7���m���Ru��εZ�_G
��0I����ƀ��f�70po��嵯�oR/�vg�2�t��^o��i�S�*�S^���:�b��1$( g��e�C�w���ב�Eio�������N(襵ʻ�1v���^��y	���ISs�o����X�5w�]..bQ���o�g{n��X����-�-,���P3߄��K$t�A��e4S�С�b�DV�k:Wt��H��zMUX
��
˩�,�0*\	86
1~Eb3��p�
���oHl�kxA���T������$�B�4�o*�Wa ���?��/�)�oj��
&�O��w�ph��$^!q����CSa��VF*�J�@�
7���&�}*SX�X:Nx$TV�"�IGJe�LU�1h̝B�z��C��r��L�)=�;۴�=
�Q�8V�I��S���x�4�5G6����ų�7��p�4;�k-�*����s�r�d�/
$˱�څ��ͣ�g�d0�^Q��!{������E�E���I?Q7x^d�qc�^��`f�ez�rsuޗ2���zo?�+��� }n�������O��˅O�?�/�����"0��^�~\y&�푼&y����Ke�/?��,>/�����\���`�~�lp�m�/8/�rѰK䆍#�T�
�&S�Rzޛ�,C)���I���h��O�f�PK�#Q��qT+�GL���e:�f�˴��M[a��\ �T@���򾙮,C�,y�鐗�y9�c.Eى_��W,�J��|Xs�15ס�h��<J�)o9U� r�#V���(@9�B�A-��m@f����.�a5����WGB��ŕ�Q�TP�ۗs5�<���j�?>(aMN�_a�����ոj]Ve�U�c]�>��Z{"�s�J���"��Z�)fH�h�&��Ybm)�uE��VԐ������㜤Đ�!�����E�ז?y�oH-���m�0l���R`#׽I�SE�^��\�Y��q�!�v	n��÷�7N��G�	�M�i��Vj]��{ q�pv�7^�=���%pۥ�NqG�_{%��.��>N%\�	���"�Q���D5GTA��O�o��;M�!���MHq"�Y�b��ӥ�I"�9�=_�/ݍ�"���V�K��1 ݍ)#0U$����d77vH�&�^A�J����.�t�"f�\�_>S���)롚5��ג�;K��B/�����%�] ��$��>Α.�l׆����/_V��#�#nI�`��^#�V#��n�w���".V7$���F�b�x-�ʶ�2,%^2���$$��}�1��hq6��H\����(�5��=��A�{���I��"n�n�����^��!�k��J3c#�"<Q؝�'��ފ���6���#��&�k������yu����6���ֹT�'ټ�ZRU6��e��Ae�@=����`6���o��9?���,T{;�Bx�́w��Ȼ��z���:��;�����WY���CE^eA̝�"��!s��.x����߂�)����u���'֡ +"����{�>+���&��#P��Jޮ��˳� ƜH��?HD�I���P�������D���4��������)	�>��ߗ[jy���}b��A_�j�"R����癀�PNO�@�<TDχ��ü���
8F�eS����|��`yC�|��eS�PK
    �\IOc�0	
       org/sqlite/SQLiteErrorCode.class        	
      �V	x��7����ؓu��Ɔ��C \!��Y2�0�����7����*�$�і���.���.,JOZ�}Ӗ����-�KۯǛ�:r��|�������{o�����>����w#B�`>��qKi�����������M��KJw3�a�#�{�p�1lc�_�
H��I�%�������))>�Pf��?ð��R����y)~��exL�_d��$��*OH��;�"ů2�b���ΰ��R�&�4÷��m�=ߑ�w�d����pÓR���?���2<%�3�c���p�Ϥ�s�������2�R��b���)��� �o��[������n`����p#�sR�#�M��������M���ɭ�t:��Й���>wG��̾�E	����Π�7�54�ƶ�6i�r0�%P��l,��&4���Xz�fH��������h����P�8���|�cѡT2A���ң#�ڜx�́:�
�[��nH�&�j1lM$j��d65K֘�t*�L%f�<<��vf���p��gS���Fǐ�d�Q
��t8��f/��"f4��|bC�et4;�xC*M�k��hrc�6LIF�44��.�y��i(G{�A�kM�5&I�ی�F_�(M�e<�*MҮ��m�&FcKז��F�b����y�РZ�%a��d�8n:Yc�@LX�HMh8�������W=a��fñ���c�d	�Z%�[��g���km��ޔ��Ʒ&K�Wq�O[���F&M�p0��6d�)rn�&-�xFn��Qbg�]]Aâv������e�fY�J��ڗ
b]�l�����\p�Q���^#��["�+�����F��=�������ո9���ul�v��-����r*)�E��f�ތ��x>��_T�Ji{��U�:��[剪�rԬ��pL�R�Y鷋�Z
�+Z�K�y�3���*J�c�%�tJFA�I+�[%QM"���jQ��(��rd�D�,Yf>[,�F�0N�$��QS,;��=3/��0�m��*K�N��2�!&���ri��v�o��9AD�'�[���6�e�HK�,������9�W�,Q�3�eOx���P6 ���]*LϪ�'�W��fx23O&I�M��O�ꦞ�Ւ�r*e��'�Ju��]4�v�����[�v�K��<��8��fg������U�FfD	L�NQ殺�n+AW��*��^�c�l'/J�'&�J�lwK�^/���"��/�͜Qq�,�G!�i9�x1ZRN�.v�<��r?"�#O���̸��(;�g���L'^Y݊�Y��OGp�[��̢!rS��2竫[^=�2ՁDj@��s��w�k�U��E�7h�N"_Q)���9��i���쓖�*"�M�My �������jK'�q�p�U*OmFť
{�y5�Q�tE*#&Lu͹��n�\��i
�{�v)�k��b�xS�c�6���N
�m,�\�д�7S��n�XM�T6����dv3�7�����Nsd�"�^N��R�H1yS�ѪFj��7T�p�#��2��)åjSP�ٻ�	��(�O��x��Vw�3w�9y�'#�IZ7y�j���y�5]���]3��,��?��v��~����X�k�M�W���s昴�Q��?�~Z�K������,hXpG�N�n�^�� w�+��N�'�+�*���� �	p��x]��>��1��$b�|�қ���ހF��Aí��@(�5���üGQwi^�,5e�H���30O�Mz���EH��;��M�T���Y��sG_��2ԡ�P�]�y?z�"��:v�aO:�0L����0��
�+Gߦ2��̱��,Cx������xW�~b�=�ИX��yu�:oGǊ���:�C�"|�Cw�����3>�dJu*�65���Rtb�#y9.W����VJ�����Q���7��h�N�?O>4���(X�ϯ������w�X��^��!4]ЉY]��p�W�W瑝���C��-u�t~?ރ&��:�U鋔��>��)}�җ6���J�P�1��S�]J?����.�~<o`�	�8Q�x�7��s�bN指�n��(��7r��P�JŜx��J1}�9���M�i�Y���y����P�Ŝ���~�b�V�9��/��UL�b��ެ���u�9�sޢ�WLT1|!���b��:_�oP�F�\�[���s�b6�E�UO(fX1I��/�S�Q�E��/�ӊ�(&˗�6}T1�s1_ʗ�(fL1��v�Tߢ��s9����+�U1W�cx�n(f\19���z^1�b&x7�I�L�c&�����˧_�c�>�d�|td��>��c>Df�u"q'�C��c%�}�}�&��XC�����>�	Z|�#�>�}�>6����`��a��>F�|d���L���A���:|l%8��8A�����T�hw����Y���y8������W`]�+��<���*܉><@O�4<��x�k��Z�F[�3��p������q���ڭX�݁�X�=��'�^{Q�?��B�ܼ�y?>����PK
    �\Iɩc�P  �  !  org/sqlite/SQLiteJDBCLoader.class  �      P      �Y	xT�u��f����	�a��u،6$�$�ц�$� Y�����40�faI��q�&�[wI�'��6Yh
v:L���q
��lN��i��q��v�6i����F#!ߧ�{�=����g>�|�s�X#',�W��>_��u�0�
�i�o�j�[�΀��|��������5P���6��f������k~��u?4P�������X��2U�o�;:��������}���?���2����k`%~���?��:��N�\ͮ��j��������p��@1�^��H�&]�6*�5R�I���f`����PgJ�`�R��E.ץB�g���e����e���T�o�.C��|](鎀�TY)�b5uY�x��L��B�;tY�I������H-gR��%E��b��e�.j�(��'S	k0e	d��ds8Nmx�k�	�m�![P
G���耝�cDH�b�Vd���u��M������Xb�1y,Nٍ���������YCv�Y`(a+~��ȡX���O�cѤ&wRఝڕN�;��ֶ�5L�v;��-G����n���Nv[��q�]���O�G5ա#dj�;��t�7��������Í$���T�d(<l'SJg7i��ԩ�.;����vg��3]ƂK��i����jKS��R��RvK"a��I�
Y�FTO��;֛i�Ǹ�{���a%H0gZkE�h�,%5}�����&3������]V܉&�T�լNM֨ғ�t�`,����dǱ�a�WM���}�0{G�иN������u��� �KĖ�J�Px a%Nm���T}c�n��D�8�RʁV�� ��m[L"=�dL']3#_��%TyH�*9Ag�ɼ�QJ�)�*�{Oa\�D��b޴-�hK't^O���i�<2as�5��:e%X���U��5��]�M�ôgv��TL%��I�4k���H ��"<�t
���(��{�I^�<VңG;��B o�U<�h��pe	�QP�d��1E�JQ&Q]L��o������JG,�>K'�5g���+��I7��g�.�aI,��Э���;U��e�%�ى$S��7f�
f�Q����C�h�!���bv��hUz�eh�R�`�˒N�#�����H��dۤ�G�T���!nk�mM�Ӑ̓������Ss�bx�����&�U�a���(4ĉ̊��t�(ak����d�&�LiB�Dq��[��j��j_O2e��M���m1�<G��%��8%[Mi�VS��)��=�W�	Gg$b["g�.ਜ��t��� M
Z���`4�
�;Q��4�C���^e�v�/ӧQ�NSv�μ�W�H�,�	a=G����/�E�)!�"�����ο��I�)��>A�� Oݲ���^��=��e�>�3�~�7�H�;!wzR�~�I@�P{w:�
�:�nbS���A+�_0����Z�������3��4l�9h���rH����X*��]���`��⥿r�M~���q��4å4����x��M9�,��H4쬆��5�� ���8=z/�h���XCj4>N�x?~ϔ�1eT�ULEL�I\�c�$�i����cO˪��m���q;�d4��ٰEr�V)��цx2�yn_����撖���N(���-��$���l�q��~��;Wm:��� ������s�P��oщ���+�i�H"v��M+���xa��p2ǩ$��jC]K� m��'p:��9Ak��"�E�̸�H��e�MZ�}���dʊ��k�t�/hY�ߪQ��)��O8����FuO�N-�[}�U��ظ/�#��꼭x܎M���vM���8vK�i��}�jqsp���vVb�F݅�1�3���p,1j���3܎Zͷ�Q��	j[�J��f1��IKr<�kn����Փ[:%ǉ����NE1�숝�{�'�4�4��ZC�o��U���}�K,���P�H�8�<��=v"Q���vڨ�%�KEZ�C��jQ��}2�L%�>�e ��S㍭���z<4��J1�3cԊOju�h�/�dh	;�T]�^�6b%z�ci�%�|3����`��e=����1�����m*����������#=��a�xK�-N�#*���f�4��$���O�aղ�Nqy��c����xh+�o��^�U麼%��`9 RU�Y��,9᪑_>(�� 9�I�r,q�w!��t0�(�>�]�K^�� ZE��s֑��d Z�A+�q�%=ɂ�E��R��_�EI��qW����c�r�<S��乏繗��,��i|�����	�t��j�4��O�!if�����/`F���?��3��CE��l����3��f0���.�9��s<T�?�*2��2�O�,��E�J���t��ц���e��r�G�5�8�1�B�v.�K�i�z�h3Na+�m�@;-9ĵ��z��zm���w��zT�]x7�l�|<�_v|2���Ǐ��+�U��Q'\�kh�5���>�u,F���H�h���;r3��4�7)��ow��=	sܟ;�&�uʿ�,�{A�S��GoY��){�:�3��ph����=�J�-P��������ШG��+�Z-����|���zm�fmx�q�:�u#��~��QG��c���g�����]��Li�O9d���+��T��Ю�L��$��t���rTR��� m��r�Q��Y,�`i�׿��9,��d�������_\כ�M�cX�_(���S��IC]�����A|^o�y6-��`U������g��AÙ�?�d��/A���.�&�e���4�N��;��ҋ���>~�]��,������a��ǆ&#�Y��$c�����u�	�(#.��b��n��[�KX0������0/��,��6i��n�̖�a��ψ?Ig?�9�WE��.��y�m�1���ȇ���Q�YO�	Oc>�(�)o:���q��'y慄��5�)�2����O�#�}��O�v��,>���.c_��-��W�"��K"�,%xIJ�T����,�z9�5\��ר���k�ҁW�\|3��"�>>��dI�������Eo߅Ӝ����Ӫߥ]�λ�X�@KO�4��i�ę}��"TI#��3��MRFo���7�O>F�PY�~̸NUJ5�����N�B�'y�[�7#D�����~�����<�S;WY>j�:U���>�:�k�r(�����Gs�W��+piP�QK��"�n=�EyB-Y�z�v3���ힳL ��|����YJ�]i�{�y�I��^'����~D�|�	R-�-c(fB(�h�������h�?��t`����(�΋<�Lx�G�g��/�ޤ�z_����wd�m��^����X�ߞEg�����wd��4LN���B��PQ[�9��,<��_�n"K=.��T����p��U[W����35���8��A�)�6���\!�^�B\��c�xp�xq������L�/A��H�2�`��dv�S��yw���8ΚE���q��3NV>�н�UԹ��������.��ܸ��z���5��K7�
NS �Ly.T�:�LQ�V����~����b��,��&��*<��`��u�ι���ZŬu���c�E>|����) ���eз���ì����~��P��GX�>iΫ�c-=O�qU&c��[��y!���+��(�xsR<S��RJ[���S�T�K�"�̕�z.GC�?���2[��~5�Py�r�zt�3"fp����7+�a�?����Ai�5�^w�wW�����r�I'�`Jf�.T�n̗^,�=���L�}L��h���z��!
*s���tk��"���Ҡ��x�	R.ٮ`�����Z�Y+�E#����X�k��ˣ������N����PK
    �\I���p      org/sqlite/SQLiteOpenMode.class        p      }��VW��#u@k�1�5&F��o� a���4m-T,b�h��&�}���z�LV��v�+׽�+��m�>̲�j�b����l��o��+�{��'>��|�ƚ�^L�3%����%n�x"0�,L1w���3�=�YfE`��/0��\ ¬
,0�5�%��2�@��L � ^�E]`�R	�hi��@�A��؍"����QTp�8��U+�r�|h2O˵��rD��e�9]�+N��	��sz&72&i��7�f�@m�Y�ӛ�lRA�l��T&K��NŒ���
�rzj]��\6�6�z:ה2�A&�M���S�5�+��#3sz��^w:�����j�0�v����x,�FcS׳����ΝjiW�BCubF^7�?�t=\'��q�H��@��Lg���Ө���ロr=Wڪ��%2;
�c�tR
WK�ݰ٨Wj���E���v�Z(�+\�.謕����b4ޅJ��XRp��J&����W�	y��n��8�sŀ��U�sG���35�����%�]��׷˫f���1.���Lk*���
z��������+:V�e�t-齃�0�a���Ys�9D8,pX��a�C�C��
�8����:?Q����͢;<�����v�f:uvy����Q䢽=_���h[���]�	zx���<K�8is�����6�l�ی�\��hs��ͨ͘��q�	&|�����[G�I�J����� �@��ZP~D�;8�'����}�(?���?I��^�3�Z����-��3�f��P���S�
k�o��H��B����i�����V��V�k���Hsr>��9��_ ���Qb+�(/����x^�+U��U*U��V�TRu�4!�&�ϭiR���ZT�n)��\>��F�4�hn�i\�F�&|-M�O�4���4��q]��DӸ!��Z�Ok�x_S}McP��v_�iI���#������:$�����J=*������o�qXt�N�Yl��a]4���7��B�Y���!�w�@f�c��@����� A�0Hh�0D�0L�"hF	>��k(�NOY]�h�o�w�0݈ �� �k{�s��7ŷ�w�-��;ݷ?��I��oL*��Rn��k��EI>�PK
    �\Iq�޼  �    org/sqlite/core/Codes.class  �            ]��R�0�#��	(���t�k<�V*�]�:i�00�d��>\/� }�N�4):�]�_ґt���??�6xEx_�A)����XȠ��Iw0�������I\J!u�4�Y�(.7����4�p�`W���Jg�v���_t��;O�H��|G��vm"bn��Β�;"���%Mz �u�V%["�̠>�|q:�b'B"K����A�[��L�M���D�uw�P�fv��/�(sڦ�m�����aˆJ/���2���Y�TI��V�nq�Ʈ��t�j�`��\�m��(Hu�f��fʬ]gP��Z�I'vv���m�t�w��ŃH��.Q�3�	�*�^��'�^��l�����.��pt茿��&���r��#�a��:��qޛ�7�`�	P�yԂ�a]$^B����
q]#���Mt�x�B��n��׉Ϡ7�Ϣ��G_ ���$���L|}���:��M�[���w�w���o������Gď�O����?G��y��3��j�=^ϼǛ��C�3�5���PK
    �\I*�Z�  O*  $  org/sqlite/core/CoreConnection.class  O*      �      �Z	|T��y{����� K W�dI����@��2b�-��>��f7����ڿ�Z�ڻ%�j�Jmm�J���֞��������Z�V�����솅������o�;3�Y|���%�%�"/���e���Y$�b�ϐ�m�,)�{�L�%��^4Ket���z���^��QVe�LF�d���+x�Lϓf�����*�l�4kd�$K�n��[���k=|��mr�/_��2�Q���d�[狼T��2�Q���yx�����b�K�Q�m*�w�;u~��7�|���^:���4���"͠��ʁ��/�y���2�r���{�2N���Z�9���c���x��;=�K��e6 �Ҽ[��x�J_%L���{e����F�k=|���祍�~/m��u�����A�Q��"nN7�[<��
��#^�T������{�r�^��c#2���o��d�߮�^�����;��9�K�wKs�L��{���et�����=|�����/{�+�+�8x�}���ҍ6��y��n����s���x���y������eh=�4����k}OS����-��{ZZ�.f�_jn7G�����T"\�T��%Sf,����-&G:e�l�D�NsZx �����ˢ���8OX����c琕2���ۄ��L�f�����L��M�H��7�n*aƒf(��ڒ�)l�1�����E��x�+��V�#�Z��`�ib�����a,�+^d2�b1+�5�I_�
�{Q;:\Kdp�/!��k0a�X��Ɗ��t*]��)���T:V�Ż�O���VY)������k��c�s�W���F�W��Ώaڜ�
���?$��	+IBZ��Rs�ӂ���	B�#ME��++_ D�bk<1d➁BZ����L���'@�R��+�r/��"��L+j�WÉV��@U"����6 �M
3�#1�3=4`%֙QK'2��DD��Egjk$9N�<�����L,^2>LSJs�BJaL��RLћ2C� ,�QU����	�ز3d74��	���~����P+�9��y�	Ut�BJ�v;H��	�K�۶�r�6�:��f킝#ـb����lE#BEK����X��D�VB����+5��1�ݛ'�K�Ǭ�["���<�.!2׶��u�c)1+�n�����������>�/n�*\7V2�N��Q�6KA�M�LS�V��7m����q�	c���Zz8�
�r�1�B��C��D+��sj2c�u�2,�+�)�)$���FOV,�Y��2Սff�~[�X��Y(TU؊Z2�M�B���k��}�"["�<)54,T�W�v��d�eb�MY8�Khh�g!�=�` �e�B̦5��H���^$wW:5�NB�9$�^�,0nl� 2��.�q����Ƞ�ZS�}�u�H�㖝�
Y�P$�$-@",N�-�;�hd`;����ں��,��
m�R�WP/W+M�D2���f�ԑH�TR�V��;.�מrR!pH}U	4'"wCNb8p̌F.Ǯ+�'�{�����붳��Oal���X��>�z�UP��;�8x.=�8O3�3t�Aw�g��>��yԏ7�.�۠{��7�>�>/ͭ4b��Y�n���	�6O����0=b�c4��~��mУtؠt����w�W�G��@��F�3��>�@"�	��0�Y���?��t~���O�)?g��d�s�����_A��=�Ϳ1���������{���/�d����a	\�`F��:�IX����	L����d��0��]3�"z �0�ݳzm����d  `$���5p)�l��/���"��2�d�+�7�����'�C�P<�����0���"���% ј �*W��������o ��o~^W�@���%GUn��p�t,܈�Aoп���>�D�:��0p8�������Qi�(:�����a1�dj�|� ���1� J�4�tA �l!���d��@�攏&�����/�4
9��v���մ�J��Kz�Ռ9�%��usBcޢ隇���?�����*��W��kl�U೓��J�]�/B�G�6��&j�Фͩ���@�����V;k�2I�,�m�6Uצ�_�nh5�t�YǬ� ��[���V�k����Нah3�Y��v����6x6w�q��`z8[�(,��Ҕ/�]H�xЪG�"[y�x,�+�L��d`]w��֮���=͛�:��!����4uu6����Ӳz���D&eW�X�LAb��r������
��\d����fr+��}��\��.aY�VnU-ӵy�6_[`h�t�V�!xY�e�VW�n�E�I��zP[hh��Z�Ă����N��
ӼS�=���`��K�zs�s�S�0.�=��u��D|�]�:y���6����5������4#r՞�f�u�	���MU���;�����W]��O�����rZ�]�5�R�}�^/ե$�=�CیHeSSx�i���.K[��:89�l��½ز�M���#
���[��Iups�>��(��)y:b���)+f���R˛ŕ6[c�.sx8��6���ěDYI����ή-��Lʒ�d�S�@)�bt��C�i(i��Jյ�	��������,����ɖ��.Y����wX�&S^�E�B�3��^P�qoɢ��%8o*�M)YJ"D=���P��r���>�ٹ���@��0ͨm:��=�x.��C3
��Q�
�+��*m*��l�͋�{U.	7iʖ����_t�����f�,c��D|�z ��'M�p�~�W�WV�P��>�ŘJ��q=�ǴW�}SV�]�Ky'U$^p谒IsP<R\�"EF��N��L������*ә�˟�o�)U[�B��T<��kRq<q
��}�H�[[�"�]I�yzYL�?%o�mEz����n8�z�KP�R����J;zi'� ���W���۶��5�􎍢������h�bNo9d�^� �X�`��T&l�q�nZ#�ԥ~ �20�cC~7ޜ���sO��H�~�u��疀�Ɂ�em-�m�׵`�rqS��޶�����ںSxx�����a����i5�CDU4�v�1}3�֐OJ]5�M�N��U��Y���U�2Y��G����U먗�ϐ� �~E��>�-���E�� ��Q/�U��S�+A�q�*�y��o�̅�'����<J�4��s���J�(���Q҃�e������S�(����	�Π߹�&�R�T��O&�ɣTm�Gi�L�id�/e0}�j��}T#�3���z߬������@�N�}�����ӗ���м>�3��24�~\�A_C�.���<\�t*��4���$�K~�G�h�U��΢&ZIʹ�Z��Z�Yt>Ũ�v�t5��M�	su�=t��Cq}�uP?�V=IO�ѭ��2Ckj��&dZI����-��V��9�N���;��wu�v����t6��=k�H��Nv^[Xy^�����A��{Qm�~�kt��33���>�R��K2T�k�ТF�c�^��ݏ�I{�n��p�^��ō�'Cg�&�����M�������%���L�� ������G�wP����[�z���w����N���{���Oo?�/s*���rP�i�~o�cY^ַ�~g�k�<���!W��-�E��}׺�Z����h���޼UcT�6mX�� �z)�����=���e�EI�(Mi'�hV/�w�t�;�J�����\�ֻ	��~F������3}��A�PV��*p~&�-�Oҏ0��5�=tŁ�c�����eu�U��O��xM�A����w7n5�~E?�_���a�_bͅ[|�ϓ28���VW��J�o� ��<9�|�u����ߤ�X��`���4���.ęc�����TN�&KGi����/��l:·�ַ672t�o��r��T�U⭼F��(~On�Pv���f��F������F�ot���
c�k �����A�k?]��v������QW�p�O���{���'���.�SDx��~�Z��p�%]{��Q�g�̷�/�з������@���Dt�&�~@��FW!�MD�!D��c$���л���h3��y�;�EM��n w8,q�/$$k2�Ȑu?�׃P�A�
��n���ym�'X�v������"�����Y���� _���D���zʀ�>��(N�ǉ���!d�C��� �#�d���1�FO�|�/�g��i>��ś���gy�~�	�)$y�����^�1_O?A.�9�~�w���n����s��[��UF/b���GHt���w�V/�u]p����\�_�������9 �]�7���꥿�ɜ��Z�s�s����_V#�Țr��4���3��?���U��.��u�j��h�NG�?o��z��^����W����l��b�c�(���7��M3��o�O������>C��S��l��PLa���w*���t�8A���L�� �������q�B�}�k���[��w��e�e#4[8� �=���L�����G������O;���ը;�z��@�����v�D�q9�د�3������ۯg�=����ނ��0�o "N�qBT<]�I����/���z	�����@���N�蟀���Q��E):���&"��ߢ;٠{����z�+��(} �d o*�4��G0~�\�����AG����9D} |pw��R:�����@����b>�U�k?���m��|��]�0"�t��]�����8������l��H�Xg�q�."]��Ws���N'��<)��s�Ά�m�1<�<': C19pv�D(�����0"�~�zp�E��=f+M���Y~���R�zUk�%)1T2t��yB��5�gQ%/V���Yœ�?��ӭ0��z�����V�c[�����PW���z��W��
�Y:��|���G/���8�W��j�'?E*��W����X���\T@ї���:��I�d?O�2��N���j�/ݞer�0�Q�x9�p�,�t��1K�.�&��i�9Lآ��%T��7����*F3TX��L�zF)�QU9�H�Y|ZV�+�PrK!R6��D1�'^�w����c0	��GLk�DE�O���>�F}�{o���^�ډ��I3V�Ӊyv�rg�͞��ǋw%�rU	� H��#K*�^NͱA���IT_�2��7��m�A��A�G~?MD^��7�L������s
��$�SQ ���B[K�ga>D7"|�A��݌�-ҙ�M�}:HvP��}��т��|�g�]�X1��N�����E�>��A��F}�jx�8v���DuP\=��E(��r��ؙ�N�!s�n��y\��P!�չ��!��b	<E��~����U~<c*(�� ��V��`�����PK
    �\I��g�  q  ;  org/sqlite/core/CoreDatabaseMetaData$PrimaryKeyFinder.class  q      �      �V{lS�����vnh0	ԣ��b�I���Ђ��&q����[���Ź`�k��!i7�v����
�������0��iTڿ��U�T��Z	��զ�H<v���c�%�{����?�z�c ��f-�!�~��I.��rsq�\���U�m!��O$�i �K:B ?B���@��0@��0j���J��<�!Xȇ���/ȝ#��)�.�:�h wH�;U�\�_��-U2���_|��5+�m�N�#����>�6��r�?�=���5�ߞ��ŜY ̹�*�3l��"4�Xv���#k8�#m٢#������+]��5�i8+	��'2�l�f�����KzS������Bd���f�6�y��vԜ�M���#�a����-?���E��`9����sPJi]�)�dV/s,�(M�z����;��������	��W�]8�m�(�N��o�̘�ޫ�]hn>��,��[ůU��L��!�v$-�a���SZo���3�IuC��j�C}V�N�u�i��+�����C����h�p%:4���o��p/�cg�o�9�*a^���E#�ƾ��ܩg���[�Q��tFc���\�<(�/�C��jx��DV��(���V.ZN�@N/8�ⴋh��%�T�]1yb�O�I�k��&��~��.�8����x��Y.���o�������jx�T<�a^�$ix�J�_��2�iG�Ap�^��^�^n���grz�aY��kY��uLp}V�J�����O����Tϱr��mEB�Ũ�`̬��g�z*�3{�,�ö����޸;t�JV�gؽ�����0	��*�c��dyqu�|%�<C'm����m���$��4k��gYi[p8��d�TOV��(��<n�(,,���.:bcQأ����*�b���r�u�V��]3�aU��M�js��p�H�A�gc�Uճ9�'\=���n��Ea�Ŕ�Շ��!�|Y<y���2�U�j�Gvt�+�oyN!V-<UG_�rS�"$rh������¸9r�t�*\���A�/O>�O�$�q���)�'/������G|���A��@���$� �rQm�k;�ڶ�%�{��[>@p�A��5%h���1	��R¬���JQ�Һu%�N�O1�����̑��e�Ch�S�(�0���k��<m��ť��#��N_�m�ÊĤP]���Z#>����_��^��*�c���J�2�	$����4�e%S�S�}g�\1͂jhư0����Ƀ���H(a�oD������j� �]�o�����h��|j�/rA����i���I�̈́	�:}�Gl?��<�w�&�T+�ә�Q?y~�����=��~����a.�O��'��}Igz�o�E���׹Ȁ�r�|�Y�s�7\��Ќ�х���1��Ol�7��w�_؃�U���_|��X�8�N�'iNQ#y������D>����P����4��t�f��a���}n���\������>���z�����<,a/�C��h�R��K|?{����R�r��}�;���d�x�M/�Z\�xS�<Va57T�Y7b�i��U�F�Z�+N���׫XUt5'ZO HǱ�f��((W��>�Z���[��M����?��少�G�T����}�77�~��F�Vf�DA��+��MU�=L����i��Z���5��PK
    �\I�|�ډ  `  *  org/sqlite/core/CoreDatabaseMetaData.class  `      �      �V[p��~{u���e�B��BlY�V�p�0A��%LMܐ�����b�2�4!ihr��Iȵi�L�����M�/0ә�o}h��������C�s�"��t�R{�;��_�9�����}��� �Ƈ!�a�ݘa��3�2�s���p��d(1Xe�y���N3<���x,�V<^�3x"�'��q O�p?ax:�gBhǳL���9��Ct�����!t�<���K,/�r ��Ӧ6������k��j
��BA5�R*�%)g
�s:^:�k��<8L"Aj�ҌB�@ʹje�I���W��O�jQ1�|�R,uN-X���ۚ=U���i�,LK(��Ӵ"��ͨs
� ����4j�M�^�+���zJ�S��rQ5]�����ҝ�5]��I�&�t��:+I�FN͗M^nZ�]�ήA�2�ɲŻ���UK֨q2��KjSG��S�E�r����r/�4{�Ja�(�)44թ�Q.X"IΧ;�J��;��f�FSk�@�-M���i!�V,K59!a:p�v�.��Y{6D�g6��(�	#OAm�
j�<7醑6r�>����BgR�f4�c�ڜa���>��RRGTK�19��Z��Q�T֭�ʵZȩE����P�s���*�_u����:�͎(E׮/�%5�Wix�lX4�u4�Ja:�����VN�v�u8�Ym�_-�"�
���+:�n�2Y��ٙ�eM�꧆��MiE�N;�w�t7���Q6s�~�/�v� ��bIdd܅�ele�c�ư���;�e�g�Ű�a� �}�{�0$#���TRA�PI �o�R�@�٩��$�02��BY��H�w�:���qh�8��uo�M�����ċ��-��+�=�/��@`sol��M���O��1ND����-�]]�1O����3�\�~�/�Ǫ�R���`2�%=Q[A�{u��j���oS�۾Ͷ�+ۦ��dgL�S�-��0���ۿ��~�U�a�)��s�ߚ����O5?m��-H�M�+�܌bZOW�ԧyz����j�ΠF�ϻ���9c�h7G�*^'�n��I���F��VH\�4��l�Օ}�����Ǖ;\�ӕ���ߕ�\�ە{\9���\9�ʽ�L�Rpבl�´�[iG��AbWPE���WQ�P� 1��� CC���Af�c�gh`342D�b�U4Ǻ���
��0�:�	w�;�G&�s�
ĈZ�1�p�Gh!	�`��о��S0�������@v?E�M�}���Țk��Wl�ڶ\O� ij� �5�9�Z��{E�2#�r�T�ŉ���FnP,>E󻐮���A!��
Р����.y��p����{<���ǃz���59<��Z��z\v���:��y����opx���{����8<��&�79��W`-�v�tS���8'.V���'P��5P�Rn�)���8ƨ;�Pg�S�������O���<��x�f.P�^��|��:~�i�W8�0�GX���+N�oX��q�ģ��	?xB��Iю�DΊ8}���؉sb�	</�1��(΋#� &�PpQL�e1K�����/�5q���.��q��}��6��-�&}�*�-./+��h�GÊ�A	`,���e
�܇"��!-���G�}�����W�2ױ��[Z�CR���/��V���Rkh�C�)Ɂ�E|o�ho�����R���:�[�Elw��PO�s���8S<<+����s�"�X�c�s���p�|��5���>G~M��uzb��}��4;Aπ�T����Qr�G{��*�s��#d!���k4�=�������#����}�El^z�B�����Y�kҋ{�\ϓ*'2��W���3��::�h��Ů�����Xr�n���d�����L��*��O��v@`}�z �PK
    �\I��3�    -  org/sqlite/core/CorePreparedStatement$1.class        �      �RmoA~�j_����km��W�� M�V=RM�i9VX�������g51Ƙ� �q�4�llr3;���3�3���c ��U����h��Z�p���8�s�d����*�&}q�i3�f�b�J/|����5��
2c1�1�vJ�X%*}Đow���I��@%rw~8�f �1yj��D�/����s)LE��
f�~��깉䶲��]m�s#���#�M�LһS�T��D���dܗ�D�8�8n��ᢌ��M�\��!"���"��:�G�m%�Q�m\�F��EO�?ُ������=w'I�ɺ �տ�{é�R��3qq�aX?zZ��'��B�s[v��9����&2�04�̵�D��8i���ޓ��~Jnu�V�D+ƪ�rk>��%BS���_���W>#��~�/p��p�e�H������%�Q@M�`��C1�Y`�t��J��y�q}�(���]�|��e�7Hj��)%Z�u4��PK
    �\I�LF(�  �  +  org/sqlite/core/CorePreparedStatement.class  �      �      �W�W�~��L �� ��.fY0�&Ѷh4��P0�F4����N`�0����B�E��zik�&ڴնV5jX�1�~�x�C���>�̰��������{�����?�
�mXH ��ql�C�L�a<"�y��8�c"=.{�E:"�.��<�f�&Ў)YO��%Ҍ�KƖ�Y�sT�q܂��=G	�<TD:��D}8�@���/�ʓ*�j�s�l��Ѽg����PH�O�xF.>+�N�8��9�+�F�,�z�l��2\�2���S��(H��>n4�i9��[�m�1�4�-?a[���=0�אK(ó\g`lF?�gmݙ�漒�L�N*��SAۘ��Wf�fi�����1��=��,Y��1o�"�mQC�[2�C|L�L�29O��Y��x� �Vd���Gb����ޓ�Y=n9j9�m͑JcZ�ӦqlB�azf�*�i�86�Cʚy�4*�9�{�4	�{��xAA��=T,�B�$ۦ|��6=��/?C�~��.�4�특�s��`M��	<xjܲm�l2
^�\�9�9h�z�^��J�0�Z�BW��n�Kv�Wv�n��oT�V�����%/���*���OxM�����vhxC��"��M�,I�'ÄH�j�g'��r�q�d�+$=7Y^d#D�i �{񖆷E��k�+��������_0����]*���_���4\��!SZc$A��>s�T|��S|&.�b�[a�E�2�<��񊂞U�
�D�f
ycgvtxphgDcۏBJݪ��%&��KB�+��THC!�깦�Y*��*P��}7��6�R����9[�*>h�+��3��բk9l3N�QvV0�;콲4�h�z�iEX65q�㦧3@uA��h��ڙ�����b�/�.��ud���~��[f`֤�O��ё:lK�6�R8JZK��u��e� ��U�W4�p��Đ���I���r',bpJ��T�T-�G������	`v�t�
5B�z<r�ƺ��@EU��ԣ3n� �qs{�ҬΈ'�6� �W/��/�`��6o2���h�D{��Wϣ��
�U�`�֫�XzXp[l�ٱ��%������ot�_��d0R��X�[������.p���x�oJ���h�T�ɗ/��
u-��e|��r�<��2�ՙ�y�~��	�7!�g���?��@/RȐHя��f���O����g��8;���D��w�#��=����;��D�mK�|�����k�R��A�'��@�V�N���X}�:�[@����÷�l��{7֓ݒ���a_WY���#�7����.i=���%zp�bPe[��¥�1��5}�����5����5>��X\eLW���ƨ�1��Sk"�oW����Uy��xFB�G�= %��g��Y{�ifmT��,�.
�*�_�*4Ѕ�؈�"�S�14t)����]h�I"F�s�*զ}��yߺ��v��sK9Yː3�:��\;4�F���V]=��>�F�~�v�}]��?h�!�>E7�o��MUl�~A�r~����
�;2�ږ+H�b�n���*R������/v�&�ic��[���� �v7�h�� �Ǚ����S����8����\=qx���\��9:�@�p3G���u���A���A��������{�l�PK
    �\I}��AM  J  #  org/sqlite/core/CoreResultSet.class  J      M      �VisU==3IO��!$j�(8��#�(���L����ؙ�&=�a����ﻸ�VZ�G>hID��OR���n&3$.��}����]ι�����/W l·)t�hrxJ�1O��&�)bLDAD�	�e6�c"��)�u�Hb2�e2uRH�h%]^SI��i9ū��@�T�ܩNcZ����Y��������K���xQ�K)���)��+�|U�k:^�񆆄�����D�?�؁�/xe+�K1��U��`��XqLC�c{z���,W�vX�^2�x�}���Q�NW���0O�y�t'�CA�v'x+)�V`�\I��Q�hr��F�e�4�:��z�
��3.����+%w�Y���>�hMkX:���0��iȞp͠R�4l��ݹ0�M�XVy�ni�i�v�[Ú� �u���zEKb�]k_�4f���1��t�W0��fٖu�L�m��8`�'���F�߯p�g���q�0Y��o3�(L2��r��5؞��r\����u��xA$�<a+'BB���m�ثpV���&�i�3���EГ��~�Y\�l�"fU�vHpjȫ��ö³��䦁�؈M��V�������q���KǛ򸛡(�>?4�_EL����(��"Q5I:�5a:����Y"���{zz�gl�@l?`ypXe�t2����~c�=�)Ze�Vw���xGĻ�7�U��7��*n�όn\�>;j�=�o�1I|?7�S2� ��������vќçva��|�r�_�g>�l�T^ש�y�������W��7n��"&��f����
T�\x�h��`�.�-V��Fs�=Q԰�?J�p�d'��_�����f�	}�S�����x�S�7!d���wES:�1��K={e��T����*v�l���)D�.�H�8��O�N��?.�շxƧ*4|�"�����j~s��a=?g��Z�0�JkqԤո[�ȞT�jLHg�q��OH��qgt~��������cxM�����=ԼC]�����\|��6���DN���4�ZM2�=��\�E�f��'e�!�R�ixͯ�R~BW�vt�ә��Z�c���<���#xP3I�ԣ{���j4�."v��Q)w)3Fx 2��&�)�<���K��/�|�H�yK�����R��i��ژ���,��Z�)���#9��:�c�N��ɲ���9��ڑ�F��������e�G�"�:���hK�s���&.fq�����Wǅj�m�t�c�1^>48X�`�A�ma�
�xK����8P�{8��57�[r���P�c��]�@�yx��$�c��U�q�Zu����h�J�1�2���s�ט8�%�o��[gqKl����	=�f8L٭�&SOͪ:��U�Dn�ŋ9&bUX�1f�6㹆�O2���QxM�Σ>܌d��<���բ��5�p���$z���$y(<�IhG�8��8Ͷ�f�?ˆ8���	��x	G�2�~%�^��[�4Kn�:b�`=�-s$"��A%��A�Q&ݗpGW���J�-�����wkxm���N^E�D���x#��3\��l�iE�2֍p�2�;C,�ݝ?#{	]q�p���Gt�	�8��gB{U��Ƚ���b�i�rTU鑿PK
    �\I�(h�T  �
  #  org/sqlite/core/CoreStatement.class  �
      T      �U�rW=Oj�%ў� �AI$lX���1�`�V�a���E���#�q6Y�Ɇ*,R�*,S�]���T��Z�,�ټ�{Ϲ���?���7 ��4����CL�aRSj��4.�Ռ�+1DpUmf�pM��\���\7b��[܎���TC6�!�b��E ��=e;�|,����E�u�4�u��qכO�m_�g��9��BZ��:�B��@w���z2�9���Mw#.�b)��H�f�%�9�744��.k��Ԛo�k;��Ę@�/:�͇f:o:��߳�y�<k���%�HĨ@S��Qg<�]$�z��5����O���l������Er�IqsR�m�v�di)+�+f6/6�2�g�}�P��-34㛾\���%,��� ��Sɢ�*XM��f��.vaŒ��N��b͖$4�"-U+��@Obs��s:��%H�c�G�nQ�dZ
��Q��tIz���%+g$��/ql�-y��h�x�ޠz`P���0``iGp�@{t�����}LU]�sY�xz,s~�x-�����~|d �$Y��^���,�Ǐ�Ÿ���
9�P>����+���|ĥ�ީ8�;�|^G��|.p�boh�+�H$���A�%<4����x�<�lVCN���ZS�-U��������*{�p��w���0���T�@�����8����]��]f��w4�@o"����7��+Y7��|j���6��w��Y������:ǰ�|iɹc�%�5-1��w$b��ȱ�����%FPo(Ef�ɪ�Y�M�؏��I1辪�\���� ��5��t��	f6gp��P}��l�L�3�.��z�u���c���)w!�GR/!Rb!5�S�5h��54�R/�TF���+D��.���s�	�ǽ�g�4��S+Qu�v��G,i�����8�'�`�_P�8�ӼSh��E(n�-�Ïhy�zg�K��V�A�V� �(yt���nT�U����q֚3��&S�V	�
]{-�s-Bsp}��s[��&�ZΊ:���|�I
�U��^%Ц� VF�j��C���x��D�C�>���M�C��,�k�`��2s�HS�qaU3T���"��%��h7A����9\����*����9ډ�W/�;��eJC:�aBǈޱ�h�J�/"�8O����2PF�pjW��d�8����H�`��,�-J�6ew�VY�I���$�.$�A�kR�Z��U�tw���t;&]�`|����^S�_����UĴ��`��u�j�+�Y룾�c���V�����bꨌ�Mb�<Z�D��G��ﱖE���E%�Y�y�`����Z�Ui�$�/H�R���ѿ���	�b��_�>��?PK
    �\I�ܴ2�   �   )  org/sqlite/core/DB$ProgressObserver.class  �       �       eMA
�P�W�W3��P����#����_y�"Z���k�:T��η���y�������+� �7���!��$�]	��}�Oe�G�J�J  �[]Hs�ˎe�j�q�9��ifX��	��
��a}��1<|
�EY���iVq�V�i�@�a<�sX�����`cF�s�/PK
    �\Ik��  �&    org/sqlite/core/DB.class  �&      �      �Y|Tՙ��{'sg&7<	L&�*b �#�A�A(��䒌&3qf���*j���Z�.�VKT++%��v��ڵ����n�Zm����G����{3�诿͏�s�w���|'���'O ��>B�*b��e(�a��F�P�G�8���T�12���L��b5N�/VjB���&�Pi���(US,U%�TK�B���Xu�`L��3d8G�j٨�����T��3eo���e>W�ٖ��u�|�o�B�q?�Z����<���R!Ի�-�@�FK-���!\��j�̋E�%�Z*CS�e�\>V�%r�Y��2\j�U�:�ք�T�к�ZP�E�6�p��j�̟�aKHmU���R��0M]�w��2�"�=�:��R���+�Z��w%�drm{�I�p
vs,�$��D�I'����b
��≮��5=єS߲~���p:R�xl�BQ��%�Z�����FS&S�)���ȎH}*�S�:�G�`K�+I�'�Eٻ�ϞH��~U<�5?�sG<��/�В���^'��������hj��Y]��2/�w:�6s����;����BJW�;"=�"��|{@_�;J!���iZ"�Fc)'���>�e;;�>ј�v{rW[*������n�~��&�H��&C��T"JUH�'�N3'IC����X�r7+���HO[j'�#	���#��-�Vo�2'&����#�m�Δs����N�����d&U��k-)��q5��mc)*��9�~^�# ��6�o{TL�{"]TJQ����x��":0���2w.���5��$��|D(�xT9L��ZER��ʳ}��o���1�s�p[���/d]��Rݬu,sⱄ���9��#�ۣ�HO����O��V���u~y��rýmȓmg�����WJL��m:��#�"�����Dm��X'%9e�F�#�-��������Ɔ>����Kb�+���H��t��;�S(F�	#�a��_)&��W{O�����K�EC��:´$M��=���	B4**�����j@�5XHke�}�� ���5p�����q]I�X�3.���E��%�$=�ߓ�$/m�$i�f-m�$��gX�)=m�+�A���T��E6�jU�#��ﴵ�JI��Ȋ���1�2i��\LW���l���e��N��msH�ӊӔ&�j|ZD�F�E�F�A��Ȏ�Ìm��k���/HX�1��I��]�GlO8��hO;��~f�B���˻>���.4o�VFg83�ӑ�H*�����u�pfK�%u�մrO��0����_�E��K���W����}q��vd_�e��֟r�DR��/&IB������ͭF>�+W�4M��e�6Z�-�e�m���Q�࣊t!��Z(I�����,�D*��\�G����ď��D�Zg'�T�˵��P����H��.�}̹�]D��R�+x�Q��L���1~��ےeC�HC@�q��1����F��b���?_�5���x��Y���i�,9k��6�@��+��v0�G���D�ݼ�mt��ƽ����a��r쯹��_�T�f]m�[��o|[�U���Q�wc
��J�V�]h�� ��n;lկvظ�2�kE����W��6n�M�۳�ک�9�g�*£�:����u���x�� 2��lf���$lu=��(�`8d�'R6���,�r��T�u���x*�[���6��	ɨ%6�%.�ZD��K��=�����9;��Ng���*)�U��I�l��ꓲ��V�")��A�xI��j���쯩ZP5��7ů_��u���I�����{"�����0��qU��;\&>�b�*����6�`���ZB�Wm�D{��̞D,g5US���1T5�Rʲ� ��ޥ�N�,A-�kX�v[ݡ>Em�'���'k���[ݩ��E�O[�3���꓋Dކ�$��*Ϳ,�}�d(	4ߍR���]~��J��/l��y[��=�<ӻ��B�8�h�Ryzƫ��$�讂O8W_Ld���U?��6�7h./u�VA�< i��9���w�g��,�U�*P��Q�ha��ax2�̰D�W��>�x��,t�䁼t��J�߲L���s�0�`*�X��tlØ�
�ڪ��	��1���8�s�09���O�F觋
1�8ڑH��j�����gS���7[��
� �� ?���ܮ�R����pm`;Vp��c��-0����B�����2���Q��(�G`҇��X�"��dX� fa�1sp5��K
=�|
1�&N�������,���� ��9�k� ;�+r]6�q=n��������\�@`q�j �G��fj]A�3�+��@Hp�7�`�����s���C$m��v�P�+ЬgS�p.J8�!����N��M#ޅ�8_�����x�n4�<y76�m�*Ҡخ����8�3�^nzλ	-A������,|2�e�[p�g�m$%ac�k��u�(����AZ�(�>�<�⧙�H�ܦ:7i�ٸ�j�Y<�`h����ܹ?|֖U��t#ہ�
��a��^4r1Z����ycd5�&�L���Z�y+|���<P����3���G�������A�h9��{�btXVr������!��'&��Z���T��}�&0���d<�H�6j�u<�e����X�#�ĖhOR��'{�t�I��Y��9��Ǘ�Bڮ5��O1 LR;�f��c)>�@���Y�/t���b����*X������!.�p��/��@#�}�'�gy�^��F�����S{��2AI�I�k�044�x�8ʷ�QL�=�)&6J�[^f]�F�Lď�����.�t���:*-3K��,�؟zb�IJ�mpźE�_��4�Nk̑���\+�UkN�;sp��*�X��#��?)����q������u��_�5���t���!��O��}L�!e0�O���DW�A�'&eT*�<�j�O���j�n.�/�9����z�9Hs���?�-<�y��@�A�A̓|��9��ʆ<��9�#9�@�%9>Er |��@��ȁ�Ց��#��Ifu6�9|'�]f|6�|/�x1�}���A���r /3�!�|̆�����G�[6��(�K�_�o9�ωU��3�?�hِWs �O���7�1%���y�#Rmf��ଧ1m�9�W�yb��,󅧔���ݲǧ��zs�c�5��&��~�1��ɜ�6N�a�YMo�EgF:�g0�#�!�J�7~AZ��]g|��k�}�ː�\yz7^�'�K{LU�{�]�V��*|'1c/J�Y�{3p� �5�f\3���|�^��\7�������ap� �Oۋ�x� fk؜a�9�7����[��vsK/��
�4`�Q,L[s%�KGaO `�7�c��f'0�D�qˌg��������H��-Ƌ���>�5~��?�A�G�Ki����]Vo�BVo��i�Y.?cʳ��k�Ƶ��m]̝W*}�0-S�F�EW,,��O1	�Es�*�
5X��@Y�rn�����`Y��h�bl��(�u������%��� ��'���/�r���a~t>�Ǳ4;�\���˿�:��ҳ�VY��{$x����a7�dQtIVX�Q��,`'��I��i�\�p��*���b��s��a���7���V�F��tp5�B��[\k����a��{�7��#�p�g�4N��~�󋦁�MS�j�a)�� ���������
��ӎ|%��W�#_���-�����o	+�6���M��s�"4�� oNo���=�ߓ������Sh��T�)G��#�r޹��J���2t����u��J��X�������/��K3u'd�r8rt�a�L��|ue��Ȑ2�3�xpa��4.�o�����~o.�fy,�����]�Yb�-Ёp�Q\:��h�:������̑(1Ga�9�f����l�C+�s�2+q�9�0��9���p�<��58f���R�E���lԞ��};��=����2����(��0Ԅ��eҠF���|}�{u�˜��<QmU�$�T�V����Y�Ƴ�4�@�$���0���y!��<T��0�lĹ�Řc.�h��U��=���O�K�pA���R�(�2��:E2Bhj��5x�^�H����%%�s+��+�Jg�E�\Gm�$�%C��i����;�3�nMC�ɐe���ٓe����E�\�l�Y�=�5�>���6�Ԯ�5p�����7�NgFk�O���i:�#�)�b��`�ĺ'�.�b,���� �a�A��G��.�d��'�~������ѲŬk��myU�a\v��� �k����:���7�t�X~�kƊ�Z�L���i��"��z��WO�F�tA���Z��X���eX/��5�o=���X�X�/�6� 6��!��{J���O藚��uA[4���r+�{J���x�!o��G����y��1~U>�v𐾑�]O�v��}�p��a�1�|���p�y��#Xh>��I�3�b�yW�O��<��	O~��,vs}�_4�ˈ�{=������tJ�F���Yn	��U���3��ߊm� J�8���	PK
    �\IY���  7    org/sqlite/core/NativeDB.class  7      �      �ViwU~���$MB[vl�`Z�U\�
m@[�f�
U�dr�N�̄YB��;������=G���<����BI=��g�s���������؉����qt�9�)����v��]�%��b���A�>�'1|*'���\�
ԲmX�p(�
b�����(����N�&3���\�_�/h�f�G����z���j�/��D���=��-=<� 2i���a��~)/��Z�$&��u͜�C�C2�-��Y�)��gM�c�툱ÚgTDfb�d�_�^:9�i��CZ9T�8����g�s*�TО���RП�.jm�Ԭ�،�Vq|J����
))�������𔂤��9���5}Az�>%�>aI�9�)���mqΫ�)Uɼ�Vs�Q��ɝlX-;�LW�H�����[TЛ�U�b5�|E8�AU_�E�rbȱNϦR��llް�t���i)q=Q���
r�K7����U ���W>��E�$(��n���F�M�dզ�ԫ�e��SRww��n+�r�U�k
8�k(�y�Q~��i�)GR���[�h���I�!n�V1d)���5dq��M����LK�L�(�$g��ɚ5Ig���k�l�K�T�JRs��*�^艬�l�TR[hl�g�T��MY�4�׳¶!��s��L�$5�MEGE��\��ɮZ�n>�}K�Go�Ӗ$�GVl�ء�e�J;eՓ�d-���ԕ�(H�9	����uGh��͇��-�T,��S���զ�]�h�|F�t��e�H��c)�+�����S�%�ISs]��l+���ߥ�����A��vD�������5<7G��-8�9��µE��wV�Uac{u3|;$fl���AC֭�v���MIl��$V#�D�֠7�>���*����l�r
jl�X�~�ˍ�9� �[�6
����&��VJ�alG�7I|��T|��e�@9Z,��$~��֭���nM*n�\�I������(&����$��i5!�f��wOSf�t���T�G:���
v��L�z�,��K笯�����$��7n�|�e���9U�C�=�ڏП�EcBV���1%KH�k�y��z��Ҹ���h�'�{�7(#�_�Jm?��f�H XO6!�ql�Y2؂�0@� ���Tw�P��!r	=���5r���7�N��}�n���E�.�|7��C�}�Flm����!�P�ve;p;=���4G�`1��e�����q��Q�#�c��p����ͽ,�;�=����(��|<Ľ!>�8����#!�\K��$c&�!�Q<�8�i�Ǒe<��p8�#8�xO0��8�	�2>��x�I�b��ӌ��Y�N3j�3�(0�PnE���8�h��h�f,�rgCt�2zT�f����j��2f �����".��+���POR����7NT.(�:2���2��W�~:���x*q�"y	kR�7�%����W��F��oo��-���Ԓ)�ݏ�ħ!�l;5�6��j�J���P���Υh�_PK
    �\I�8�[K  �  %  org/sqlite/date/DateFormatUtils.class  �      K      �V[wU�N�4&�R�m��Q�
Ԑ��N�d��2M�%�$S��>�%]��]����k���d:�M��y8�9����s����Ͽx�p?� ��8�#���}n�pYn>�暂������<6�{YA�1��b\Q��xKA���
J�e�;
���3�lY��	�\4KƬ�\ʦ����{f|�.�F�de+ekR`�l&�t~�HJ�T��>m��+��x�n�`[�IMʬ�穓�TK�M�,t���y�2�Z6�nIaȵtz�s��y���.�;��>U(�3�����D%oQJ󅲵�VZ����\$�6_ə��f��c��ojG:k��H��H�����H�D��R4˫�]-�W'G;M�]�P,r1'�cڶU-s2��"M��	L���)�ڗ��J��Mjbm�zQN��6/��!�^Օ�h�L�9oV{A�9Zo�K#0�E�by��δ�ܳվ5�B�E�L8��[�ޫj=�]{N�z��˯����G����'���UsV���e���8�kU�qB�����z_�K8�"���T|�Ox�)7���vA7��\��R`�����x>?b���L�J�/�J��xE`��G6�b���i��{��mGy�M;���ب4�b���c�-��d,�χu]s���K8���*b���F�q�?��-�������V��_d�_�᭿|T֪eϖk�Y��fe#�&�~c�utσ�<���Zgj����GE��Nz�v-+ԮݹŌ@jk-{Ս���c@ �jPo����#�:up�������A�=��U�N(�E�B<�N��}�އ�P�N8�7p
o:I��'����?E�1|b�~tɶ��%�^I�o�4 {�$SN9�g���ѱM��k�
�mZ�c.!��:\i��7�A����k�H�{�0M�L��C>��^O4���Ckg��cV.?�*�pX�n��K�GM݄���	W�)GO%:���k��&��j&pޛi{;��-LI�:�.8L��/�"ǽR��I��"�7C��_R�:�)G?J2���Wgg��cκ�sޜ�����^x+��M%^�l̄{0���R��J�8��zs�K �t���9�p^!�m���)�y�{TrG�\!W���A�9��(>Ew�X4�Q�c1�?��E��"_;�"N�@'��0A��������@k=dzː�!�R�s-!7t�-����K�.} C�c��4u;��-(1�풨i�%j{$���IܯI<����v�1��q�	��a2�K�;��7$@�C�j�t�'��\a��(����,O��u��gש�T�
��U��Dedޓ�\�PK
    �\IJ/�  B     org/sqlite/date/DateParser.class  B            �Q�N1���ʢ���x6f���+1\�����[]�Mɺ�n1|?��2�ݨ����2әi'}{_��� �Q�>�����h:�/�e<O��h���aI-��؄1"�׫D,�Ty��p��V2F��]x�
�[�Rabn��9���Vs'�Ľ��C�f�'oe-+���gb#ɋJ�%���s���ߕ=U�m���?Z�D�H�����M��i	�J��xΤ���o�W�#�T.���&�P�[A�������lz&������!�~�a���G=�v���PK
    �\I��� #  �  !  org/sqlite/date/DatePrinter.class  �      #      ���N�0��KIhʥ@���`,�ح�U%"�	��$N�*���>�C!�K���zȑ���������p���sC'Vz���N�g��Yʳ�͍�Y2&������nĸ�M잧"��nG��t˞�q,��z@0��C���r� /&���i�}�<ɥxV� ��@�7��z��Жi$�P�Z�6�_"4��|#ֆ�R�Q�V�H����\�:�,:����.wS\!�T:a��T�";e�^���! �8^�`]���Z�Z�Zj��_�!�J=�I=�D�S����PK
    �\I�پp  �  $  org/sqlite/date/ExceptionUtils.class  �      p      }��N�@��)�J�+�]�;0��@���h"եq�	������ҕƅ�}(�i�m�s���sf����
`+&t̛Ha����%�tUzR�R��	����	[z�{��Û.U�m����(O����!Ú�m+�v��9'S�k�+%}�XI7�0�P��P*�~�-�{mˉj�R�6;��H�Q��
Ce�Ӑm��n@=�գ�oN평�ɳ��J�� �g���2��P�S
�gΩ��,��w��ؓ�y��w�IsA:�i�1�����{s�|����=)�h Y�2�<#?���H��Q�鸸���WLd�g(��~�3���q�x�'�)B��h���@����YAKyzu��$�ųq4�	PK
    �\I�Fk�  �  &  org/sqlite/date/FastDateFormat$1.class  �      �      �R]OA=�n��~���u��|(6!Y})io�����٩�g�$���Q�;�MS��D7��w��{ι3��׷ ����'>�C��4D>���d��K%�Cy{��൲�`X��ƣ��Ǽ��g	O�\K�^��ʜ�~��Э�繠��8Ӄ(?K�Q����9����7[o�����p���v���Q�� �-ՠ9A�F�ѱ��L�Y�Y͝9z�������TS�3��M��)uZ��Y}��?�;ȈsM���ȁ�f�I����\Y�'C�?o�b;�X'�-���?^Yu��w*I��l�f����0���n��ױ�%��yWΰv� �?�.^�]�}ʴ�;�)�(2���%�JJi�:����I�����h��Q�}G�d���K�/�PGј�6��e����R�����K�$p�أ>�4��+��������!������i�T]q.��PK
    �\I�A��  �  $  org/sqlite/date/FastDateFormat.class  �      �      ��[xTW��{&�\rHJH�L�X�$��T�L� ��6Փ�!�t23̜ HKE녶ڪ��V�xCm�TPl�U��V}������7��\k��3gΜB�Ú��Y��^��7�{�:�M�k�EP�/G�<�W��k,���,�%�o�x!��·�����nߋ�/p���|��X��ŋ,.����%V~��+,�p[���WY���U�B�qkq!�����0~ʿ�E�:~�Ϲ���e����c{#�_��-���ތ^,E�[�F!�g��B1��N���zs٢�g�a=3m�����N&I'��'쿇�B�n`���ၠ�Y;����!����S���d�0�]<�I�F��N�/W���^��#L�gus�@�wϥ����^4wS�R��N�P��ΚFA`���AK����z��ʫ����֏fBf(E�����Q8�����6&�Yc��ԨQ�G3Բ9���O��=;�=hR<�=��5%s)8���0���&�&˟��{=\Y-�f:�=��2���|܇M�,���ۙ^��2R���\��<�� ׍4��P�xbv�E�4G|G<� �[*�nf\ޖ�=ʽ_��Q��O�')n����w���⻫��f���c��	�5�M��z>�i�0'�Ź����q�0Q��RF���Ӄ�^0�Hp�P�K�#N�F'���Sʮ���i���M��ݗ62csŴI�e��B ���ܻ����ۙ�ٱ����9�%��׻�������S�L�G�=^�&/���S��������\�i�F�����6W�F���
{�>��, T+��r2+���)V�Mx3��9�2�<T����;����#�=���_e:�e����<��(m�gO����W��uv.�;Cv��RK�s��B�>��Ie@?�4���Ğ"�r>���O�Ĵ�)�l��t�1��9���E��S�yu�O��	�6sV��3=�Ϝ>4��Kcxk*�v<rF;HtP^_�K*��읂-'��M�����w+���X�-G�{#,��X�i0�f���\�X���3�?랧��h�`����$�S,ΰx��Y�#,��	|Rçp^ãxL�������	O���˪�L:3�C�X��{5���v�������0��i�����bo�-ݱ��<�*�[�����ez�kM����qew�cG$4������3����֛�x����X��U}�Kv�Ρ�T#�i~���zun@ �x7у�vz�m�w�@��.�����Q��VG}շ;�w�-�w�z/�x1Q����ކ-�i�Sm-��_�%J���K�ḏd��fJ����B�s�"����Zep��� I�R�~�_�T��	�B:} OJ�RKQA��>���No��>�!V�a��G��]�7�E�[m)VE7����|�"wGih!!�<:��zAު�qv����u���7��P�}��q�p��ȝ��݈�B��x�n�?wQ�܍����z�܍����9��ݏ(�.�J�n��=�=�@�AEn�.w�*^�x�2�˛��i5�K�HS�ܧR��v�Wq3�s0�63l3�2sL1�)�;ڮ���NIr����E��;H�tSQ>+�/֋D/��(�3�."Ǆt�����Y���rq!�?��:fP�q�Qr5�EW�@�F������+X\v����yԈG�$�Z�b����h��h��hSApi��Gw-� չ#��������N�s���ۮ�EN��G'��zP$W��T�Q=(SJV��č�����tN�ӔQ'mT�Ғ����F]�A}��m�N��nu����N��
uF���Fe)�Kݬ7�=j����\z�h��!�j�-j�K	��Է}�Vgg�I=�G]��݇j��I��8����������'���d�(�yR~LB�u1�sS���9��4?.C�ׂ��M������P�MrJж�i-�.f �8�)���m��m��iO�o��n�e���^�_u�e��iOO-e?Eڜ�X��y�����50�KW31X��
lB$��;��������~����d�5>��w�;<C��I9���kX{tmM�%�S#��n��+Kx�����8+�#QB�;���;��~H���N7��<Wb_�3��&�m���E�Y�2�Q�%�/IW�b��tI��� PK
    �\IU��Z&     &  org/sqlite/date/FastDateParser$1.class         &      �S�n�@=�8vq��].m�R���)�>�K���!�}k/����v*���T<����!f���%{w�윙9�����{ 7�c�Ī��X���+&�t\5q��u�N��]���i�$�`�ꆱx0|v �G� "d���<��4�����0c��8i'�Y&�\�&��͞Ga.܀�g�g�=�<�i&��N���8Q��<�J&��D��k��ow��c��0r��������a<h�v�#��:���D�1̟EN��h�d8������[����ϏF�X�d��b/�����%)}?��$#�}�&��u8gb��&�l4�MyOWe�E�:'6Cs̑b��A�����'`����S��&��d28�3�C����,��lQ#��s�dL�.ͣ��}E�o�h��l R��&["���[���_�6��}�M�����R�1#���܈�%J(�Zk�@��}:x�ʦ�����o�eI_R���	��U��+��o*ݭ��w���t5�;����.�A�%*F�bQ�w8�9�T#5,Ӫ��L�r5:%�Ih�OPK
    �\I�D?>K  ;  &  org/sqlite/date/FastDateParser$2.class  ;      K      ��_KA�ϸ�[�ii�!"|�����K,���ubܥ�5��P/==��P��u��!f�s����|~� �aӁ�U%k�3���6�:t�}W2�[ʓ��QW�[���Z~O�0*҉�á
�Mϓ��EH�;-����V�������*n�	���N�}%����b仪�8	i�zL|��MO6T���_��x����i?P��J�Cߵ��G�a{V
��#�h�����M[�p��v��hQ,��QuB:r2��7�׸oG����0Gui2�y,Ą�X���!�p�/s�e�����(K1��r<_@1vWhwh"�m��u8�PK
    �\I���ai  ^  &  org/sqlite/date/FastDateParser$3.class  ^      i      ���J�@��4i�1���Z����;��b+B��i3mG�D�T�7�>�%ޤA�;0�{Ν|sf>��? ��ԡ��aAC�!u(1�뵍}*�%�u���-�K޶�����[ܓ��M5�K���9��*6�}Ar��z��k�@�-NK���	�󅷶w���Ja[�F!�%�����-n��n�s��7�yz�zQ��(��n_�;N�O������5D�w-KT$V&�bؚ�e�"��#�Gy3����A�^?	�t[��I�Nj�|{��Z���STG;0������t�G٘ss3Wz��<C5_H+c��1��C3��h�T'�Џ����0���U����r�PK
    �\I��:i  ^  &  org/sqlite/date/FastDateParser$4.class  ^      i      ���J�@��4i�1����*hE\��P-[*�O�i;�&���O!��ܸq%��|(�&R]؁��s��3����`�%�2�ҕ���^�hѧ�ق!W��8��¿�m��Bݳ��⾌tb�aOF�u�_qx��u�[G��lsZ�<O���~ ����tG
�f`5
��lٹ���lqg@�l3��u��$��Mo�[�*#Q�Mݾ�w��������6D��lKT�Vƥb��e�"��'�Ky�������~4R4)�T퓎�̦����HS�&�.w`S1!٨�i��Y�1̼�My�j��VFh�#4�f �f�N#�3��)b6;G�N��)�.B�PK
    �\I��\�;     @  org/sqlite/date/FastDateParser$CaseInsensitiveTextStrategy.class         ;      �W�SW��f�aUD�F,�R"b�Z@��H*����\�%��M�� ���ٗ��j��i��L�3m�L�7t�8���0�{Ͻ��s��;�����/�X��`o��E���/Ix�'^�3��5�+���b��U�`1dD%y07�s�n�<��An���87�1�_0%X��q㐄Q>�
#,�����ޔ� 砦�"�� W,Vb��Ү�ʈҘ��Xc�=�"�ۮ��*��j
X��CI�rQ��+i������)3�������hK�LH�Ԩj���!�VM׬6(�v�@�(FK~^����xD�9i�ڝ<8�{���ԫ�ӓNU��1zoM�吮�F{L1M�lqn�5��&ZC-W�+��MU75KQ���aR���7���pL���M6v(�����T��YvS���:H��`e�h ��hQ��r,�A�Zʣ�1��R�h�}�]0G$�pL�qn%�MΣ�?���Z,B����E4d�k���3��H�	����5RiyU@��Z3,�@�j�ΓW#38HJd$�H�z��� ѩ�J��'�4�j�ƅ[�|%�&#��2jQ'c�ޑ�.��p&�N�"����2� �d|�S�e��N�Y��q(N���q�/�<�M�%\��!.ȸ����߿QK������d|�ϸ���/pMƗ�J���&�c6p�g�-U�O�[>M��Tgm��Ԩ�dD��"o�	K��2��u��U�������c�{fX�_%*��]��s��,�N�~P;W]�4�5W5�����Y�z�*����uy���s�-�G�HY�M�䠳}�Z���V�#)f7	`��� �Q����9�_����]c+�?D훤P�(��n���n�H$-NI~���¹(�( �/�fiA.��6?q��8��O�l�?�����gO�G�!�p��_��bl����P;������ ���Ŋ�����Cӧ�0�T!��7W��G�Q5���@)o�4*���~S��'i��@�ֲ�fa9��haB��X x�ʆ�m��b��}�p݂���0�"�)N�s
��\�r�+�3���0���X���k�{����&���u(��p�ax���D�P�F��Ae�bch"�6�Ёe�1�4�(]��z�q��=z���8t*�-^D+͖�Z�tFj����hm)�}J�%a� �Y	�$l����:Z߂�)�@��g+��PZ:�E{9�)��y��Y�
�I��,6xE�m,.9<�r�����	T����	<&ްE�|,���H�(�ֱ�hf'���6G ��6Q�t�_���a;�䘊��E9��K�taGZ�5�M3�<� =�����]�,z�?0x�}�I,�B�>���Ņ��.�4V���J�]�Ka��l��;�����I�~k��W����9M�JJ�4��T���e�d���.`��0��avo�+8Ů��tR����� ��M4p�ƧI�&i;Ӆ2�]��A�1�� R�P�=l�%�髽K�0�`ߠ^��w5���3�)��OE����mуv<�PK
    �\I�K�r  �  7  org/sqlite/date/FastDateParser$CopyQuotedStrategy.class  �      r      �T�NA=�-�vYl��|V-��-���DK@L%BM�ݱ�.ݺ�5�6> L� ��|&c��-�6Ҙ���;s�{�ܙ�?�~��;td�᪁k�n �i3�Ցӑg|�z�<X�±�k��[^tx�Q��l6�bٔ�]��\�t~�!Zum���ɦ�h��
�	�u��s-�lsO*�;��OsU�u��vaD��\o6�Wu���,�\�Q��82E�0�U�+d<�/�l/��~'
�H.���,z�C��[��V7�8��-��*�>R�=��oKǦ	�k� �L?��#9�OF��=K�Jf�O��̄�yq$t�0������2u,���[��.�l�5������6�t��e�a���Ιjg�q�^@��[��.�O!U��V�
�KE6d���O��G5�%|?[.��z[��ڽ=��?ck2��D���NǏz\mYz҈I�4z���V������{N����ah�.v�H!BK�2�Ҹ�%�]���Gh�ψT&R��a*7�G���(�aDIf	mI��Q��oR�]�я��%�b`?0�dG1֕� >��9
a�Y��$C�i�)�!{��=I��8&�DL\&U��T��
����1��RP��
Qs���/PK
    �\IHO�^#  �  <  org/sqlite/date/FastDateParser$ISO8601TimeZoneStrategy.class  �      #      �VmWG~&�eY^LxDLjl)�E�$� �.�W�MH6������<��Զ�S�i��G���$$����ٝ�s�>��w�������'����:q�@n����n�6p3f1����#ǻry\���힆�4う���A�t<Ա�����<O�]�@���Ҋ:���&���f&�����������z"�8���[f��oy"��s]��v�BA"�l>-l9�'�iZ��
�m2�[�����G�9�]��~`�v�vm�Ck�8���:�Mq����"��6!�ʦ,g����<����Ķ�r�TI{S�d]Q-k�:N���t+�^��0>f�X1����&Gd��ΩE��`j��"2��7m9�M[{OrE�v��a�	��sj1C�ID����	�J���r�M�����p쿈G��/�$\��ɔSVKFF"[̧Ĭ-3�\�4M|�e�4��'��a���$���i�&���a�D
i��)��P�47�4!���t��$o!t3\��Gd,g*�)n
כ�N��gg����R��t�U�e��K��2��O���+߅o�?�\[M;�}$��vd��p�A�x����ۣ�C�Y��Vҩ�r9R
��I'�jn>�",�U������s��ԉ
T�ߩ��O��i��8�V=V�U���'�ʺI���[���$��w��^g5���o�G@*��N�M5^*�!5��EZ����P��v�����=��C�Fp��A����Ksm���a@Y2#+��2�<���7��+|;���?W@	���I*-= ؏X�A\S�*C�@��4�;��M��ߡ�@��{�[ޅ����t��,9eQ\��x�J��������W­����0}�}ʺN�r|�:�k퀎�1Z�M�~��'�p�.�������hx��t5��C�r��.Uص���Yt�-�x=��0�Z14K��c4J��wqΉŧ/��Q���=�-�h��nSv��ە��FQ��u
&O�<T�ڲI\T��$�Et��ߊE*��c�F�PK
    �\IL4v�*  �  3  org/sqlite/date/FastDateParser$NumberStrategy.class  �      *      �UYOQ��m�aXZE��"v����Պ�f,�c[�S�@}01&Z�5��d<�N)*K5M{���s�sf����U GqKG7�iC8�Q�p\*'�t2�Sa��qgu
�1�sF5�gh�o[���2�;o{��x&1K�x��Z�vޚ.?����b�!K4[Xάpm�W�Ao�.1���3�+<+��`d�y�wD�d�?�-��t�c{Vڤ���(y$�n�r���f�%���'�A��-+g-1����g�'"�|.M�v>7V��)TTA��`�)�/ٹ%"C�'^�*'M%���7��c�e�v�ki/0,g�0��,�Z}"���ӆ\��i�_��,�n����L��.X���|ǟ��@"3Њ6�&�Y���M�ϟi�d`S.##�+���T�p�!�TB�UY\3�@Rô���0�_+�p�N�zdxM�p��`��Q��lE;M+i-ykkٱ�F��X�����q�M�Yޤ|4�l�[T�O�ꢑm�Ywe�tk�AX�8���@�эKDiui���*��z���Bo$��BR}#��2�4N�)�>�%c�ߑʱ�~[ �%�+��5�ɶ���P��e$�A�
:@�����VHZ�[�a��F���O�J5џ� ���`��*Тa�稕�h��z@�G$�h�����UU��G�U�G������G�����y }�>�-(�H�O�@���c�]����S��~B�T�V*��T�+��%zЪ�N�)}<�7Y?~#|�,��"��R�nE~�&=��?�!\긨�ÿ PK
    �\I��h\�    -  org/sqlite/date/FastDateParser$Strategy.class        �      �RMo�@}�8qp-�w	%���p�Rq �R��z�m��V�����N��"��k7��Z�w<�ޛ7�����w O��Gm.��<< 46T����Jw���'�$�U,_��G2�#͙+��X��(�_&��J	ͭ,��>Z�8�I_�4�\�'I���d2&�i���7"Ie�9f�XE�EG�e�0�ʬ/��C���J�Vo�'�E�gJǴ2�E�J�Q�L��`�v�&{�	W�%N�����9Ӈa�VF�qN�'^�J�\��z���:O�h��:a�K�&y2��ʜ��߀��Mu4<,��	s�x=ړ����a�����օy�p�+<�x%�]�
���5e�g\�U ����ْ�V����)�Lgʜ��9��ء�-X�jQ��z`ފ�=�5f�h�Qc��4�l�v)��W���L�b��0mQ�ܵ�E�����m޸��q}ܲ��oPK
    �\I��a�|  �  5  org/sqlite/date/FastDateParser$TimeZoneStrategy.class  �      |      �W�W[����JW�� ��YFIl'X`G	��ԽH����J���8q�%m��i��钥M�6u�N�>�����O=y�C��.ǭ�͕BȦ=Gg�|�-�-��f����{@�wc?T�.xwÆ�Nhn|I1��8��7�Sn��|�Ő�2�nlG�	S|�bXpbQH\��.��I<%��2>醎��̧��i1|Fl�Y��3B�s2>/�Y'�sc/�w�|A�<jJOL���L���sj6G����5�R�d0ffu#�� ����F�";o�`,�5�Ĉ�!	WLO���j'j��l�Bl͉��d�d`��p�ș�aN����)�`p�FϜ�M
����X[��	�&�����q\7t�$�pa8WSZ�$�N'(��ú�E��ZvB�Mi"9BhR��.-��K͵�!K����t�VVmz�$�9��ڰ�D\�ԒKJ�0�l8��r"���l2�{"��Z0A2��j���N�vV[�)+�rU+e���r�����f��8��z*�eI�>f��T[+k_��qY_�j��ĸ��.2�oB�7뚡`2��o+3Z��e]N3���PI1�?:`�iMm�SF8%qc��
��� ,�;��g��i]Ԡi�^����cx���<YM��*��.�/)�B��o(�&���۸"�e�������Ȅ���
����xE��xM��������wH���G⸐���?�x��'t�����
��c1���Z�{/��?�񦂟�o���U�z�6
�Ư��k

XQp�
���]�P�k�� ���1�]7I�����&��a]�kSO{|z�g�M����3�#�L�!��3��� o�xO�o�>Á-r��S������mp9bj$��3�;�}[ᰳ��؎�@l�\$��"�ɡs��C�Ĩ�]z���M���ks��6�cj͠��t:;������t��@]R3#V���罵:��]����B	qTS2���U����=z:7�G��M���z��pg��#�_K�vSn�q=��x�0U��=�-Um::{^��֦<�7���֐߼D�J>��K)=9gyO&��a���C�d��0�N�^����qA[�i�y��2)�$����^�U��� /�95%$�fX�f�p�j<��r���3��Ԛ�����k<�j��6z(�D���� 9b�G�"�N3]Ԫ��CG��"�#]a����U�Z�����S�~���h�;���)�}[5��q��22<�E��#nz���":hч�CD�SA�K�}��ﯠ�B<����V�i!�< ;��V��o�6�6�
�k��G�HO4p�ď�[�-��x+�b�9��
p_�c/	�:����w`�:��*^F��WQ�1U��U|{���v�⺣J�QeG���e�3v�|{��O��!�4�ix�������<Z�haX��>�+�b'�t�ه]!�>{�k���ZTY���@��6)��U��n�ﾆ���}��4�����`��M���K��v��<ȝ�p�9=���%^���v���o�Uބ�y3�D:�^|�[�7ކ��]l7�ͺy;�v��� ߃��C����I<@�^z<�8�n��a�.�0N[O�S8Ct����0a����������CFTƨ�1�����&�#���1�q������FPFL�Ŀ��T�dVd�f����Nٞ�޴�'�#�F�Q��wY����k�l
%Cb6M~�4fp�h�m#�RDX�:����,�*�K���P]<TJi��X�@i%$jX��FE�#J�a`�tɈ��|�hd���x����y?\4��߃ �G��c�}x��#�Ob�?P.Q�I4��(�r؋����^�Ǩ�c��#VZ����[8D� �sVf?�!������DB�s��%ɍ�Z��PK
    �\I�Pn�B  �0  $  org/sqlite/date/FastDateParser.class  �0      B      �:	xT����d�M&/dHH$	�H��Đ��C�IX(3/�@2g&�2��][�%V�� 	�J�ު����ֶڪ��9���y�	���w�}w9��s����|�I (�/�0��M%7�o���T�-�f!7�[!��Y$a5������p�2�-K�q1�3$\j�	x���V�Q��؈MV\��%l�`�h��V\���u����B>��u��LFz���f7n��h�2����[��7w�O�M7K� ��b����K`�u|�:��p����c��-d,!+��ׂ[�xne�I��
5��_"�k�o[�<�ϸ/��b�Ђ;y�.F{��b�u7�y	O\�c�Y�r^p����U<t5��F�ky�:+�ŵ���L�����nn��fn�rs7�������m��������]V���=�r/7�I�g��z����|���Xa>(�CV؊����%|Ă��Kh��K����p�p�
;Z�"�����!+\��11�>.�>�p���inŬ�V_��&�WZ�AwX�؆ ��~%X�����m�q����`| ��R\����¾-J��5�ͬ�l[�+���%޵����ݵR	�|�
W���^���nx���W1��g@Fղ��ږ����e�ͮ�z�Q�ɽ�]��u��<�.e������?6���w�a����-a�dtۣ��.��0y�7H̢!��
��w������eQB�:DA�C�Z�M6kH=����X[v�����R/��ֹC��,c��Q��LOo0H����p�O��e�0)}|��Q�k����d�NZ����ktK�c�w!Hm�u��$�����3��7��`nբE͵+]U��5��j��׷�6���6����j��745�.я׻Zk���G�_U[�t}S]�xNt<ф���$복��哵q���8ݒ�ͼ�����p��<QV�It+\�+Zk�#-��M�5z���z׈���ֳ#Ѝ�������y�#�&����ܢ�)�/�GF�ϯ��ս��)S,Z�&��wm0%��#����K�1W��(��i�ݢ�i��H�FC^��d��&�~/oһ��(�!�l&Ǥ�'�a	�"�Nq��9��M�0�0�}�雄k�y� ����BJ��@W��	��OP��iz���a2�`2ϥM��͐��&g�n�^�R󿆙S�"��>C���%�&%s�i��5��s���x*-��\��a�b�"CPӻ��a��Y9���E
���Ʀ��H��� 7<�$]_ ,Dn�t�:U#1�8"ԣ�郊۫�@����4$.O/߆��*b�1ã,"��[=JO�"lH�g%|��'bW���$fU��}s(���&�aƱw�&��a�1�7Lz^�^B���?9ƞ@(��I6!��h�Y��b��>:q��=����IoH�J���Q�Us\<�j�G��f�BǍ=��o0m�܇������Fר�Z��t��5��9n�-t%�I��nH�vէ���(�K�b��')ґ8�[��M�!�Ǧ�X���9�_�O5�9�a_��.J��:���tl� W���N���i��Q!�Q�F��֮���W͉Bq<��H���=����,)��Zz����������u�!����M�8�t��~v��X�<%�Q6k�ĭ�)�<>W�sїS����)��T�|O���:�ϵ�7X�㨒5|��|'b��0[�t'ó�5X!��p�w�]2����<��G�c�#�H��J�C�����J�{�^���-x�2�c��2��*to� -��p��/ʘ�/Q��e��0MgÔGt������tW�8BG��kɄ����=Ե��
�*�k�1e<2��#��+��x�%�or�ANE��?��e|�����2<ߗ���2��?��M�����>�i�����;�[{o�����^e����J�_��d�ǩI2�+���������;�n��42�����3�tO�w�=8S�?��'RD4D�jdLb����H���o*l�T���j�j�����C�==�`����rd��ln�\{UM�u�_Ȏ36����8~Z|�sv�SqO�zV�=2��o�����3�ɽ��2~���?"�[�\���L���ծ�Z����oִ�1�f��&��Y9
�P�ǨC�<�ͣ�<�� 7��y��ǹ9��S�ps����j*~B̭Y#�3<��SR4��ZB9/��t6�� ��q���),��"T�%�cba���~N�~��#mrSs�2^vaC�3R��9#���%��Rg��iqFV9#���5Έ��:#���fg��	9#�8#ۜ���HAA�`�Yg:����p9��V��q�l������S�7Ɓ��^B~�d�%����By��Kf#T����&��.�\�,9s�wG��ԯ\(zE���קKw�i��P5M�[�74�v�
�%��a�%^1�B	ǂ�CYFcQr5�<�=NH|1lP�����dŗ�v�r��������/~G����ȖBjH�
�y��%��b��)�ܱ�bXUw
q6od	��S���$�*�mv��7��cTQ��~a%1i��@�ǔ�O*�msv2bt^SG0�K&f,��$j�oV���.�h����^���?f�tLE!L��$��N��m�:'�	Ba��$uu�1�8��Y�(�OZė$��G���J[Cy�1m
�^����n���|�+���H�ĄE�������L6;�̘O����B\�D?@����w�
d	��:���Y��R6���N"�:�z�B��V���up�����_���c��]��C:��kߕ�դ7�j��H�8̕�HB��ͷ�Y��>R�N�9p�j�&C�{��}��X�~&�R�!���8U�'����
H����}r�M0�K)'":?t���~m�Q���5xP��4���4������<���4���0R��z�8�!�� ��:��%8)*��Sk%����9ԅ�#���Q)U
E�Ee=�Q�xA%���.��� ��`v �Qr ,�%!�Ҕ��<d� k��Z�����}�> ��B����rMC��6��2�2o�ّm�y�l��0���Gɝ�LG�i��<Fq�E`�v�!>υq�mȂ�I0�T�	3a���0vC\p�&����Z�����	狤fX��	c���͖�l�h���K�2�G�^�W�
V��k4o�WĊY��H�S	^��	ޔ�g G!�S.ZU�Ji?���`	'�ar�и&�,��[�¢ͻN��6m]���xn� L {�46 �a�a��8 '9h�I�A��Ń�@�*m����-�f�#��h0��( �^�KrM��� �h��>
�JS�W������+��#�y25���0##.)9��̢���N9 �y�p��`�H*�'k �.������$��ta�teMt���=d�!��d�瓍�$+��l�F���ɲ�'�~�l�Q�7H����d���!4�J�8N�'����g	]�edL?'Zf����P����=���w�m���_��L�t�5�����%L�;�$�zu��i��<җ�$�$xW�?�,	�4�(� U���ɤ��4�/%�jjbA��l�,����M���_�l�7��t���$�-���H���{��������m󽴚�p��i�s��9��9,�b�ns��t>�I𭽐�<қEx#)�R������J���> ��wҢ��(�F�#�I3��Q�G�O�g̂јA�]S�B9���|����K� |�)�=T����y�Cl���й�A|�Ĕ� >�]��V�ܜ�ŝ���j�p/�����<U�:��c����������m����E��ѓ�opk�ZŖɁ��	��ِ�9:��d�C6��?�g�1���/h�K�J�\I�]��A����$��+b��4�.�s�-��'�{t!��N�sjڌ�P; u�G ȧ���!X�gKtuQ�ɲ<C����T	U�a���ї�WD��pd�L������Jt�X����1wj��h$�U1Ga%�����%�h�SKh�Dy<Q��u��-I��=�E�H%-O��H-4��6.��:�M��e�~��P82�2�DП��]p"�l�.3�WJ���s�lR������;�"�l���]9�-`Q��,��|\��p�R(����$�&X��`.��>b3��2�BY",���%�c��;�f��&hG+�3R�ӄ_w@�"���� 9�/`~�
��_�5i-h �82W�6�2.`%Yy��R�Z���� o7��S@�^ N����2��q9�~mO̎S�5ӑM򲯊����A9V�*�h[�������y���<������n��q#LD�F�b;TcԢ�����3���V�6�v؆;�|� v��+q'܀���g��'B 3�F�K�]B�k{D��=8^���,M�ǃtR�(ݫ-5}ڧt�V��A��:B�h,�<#ia[�Z_�Sky�{)����)�A���z&RlV-�S�~�����pZ>��;A��G�ͻ!OD�g���1}��yD��Lh��f�	�d�Y��'y4�8T��Z�<�ӭ������AL=�]:~�F�5F٧�)��T�a�pvH
�|�*K4��Z����s��FR.����\UT��^}�}vҳ���鹞�[ts�i�c�Lx��#���(4��G�^��_������V��;����m�r�`m�3��R��n��C��g�;l�������0j]7=�y��N�&��>�Є����j���頧�=���ܯ�O�]bg�9�~gf@$\�>�!4ML+�!���{��؅���/x	��W�x~�7�Gx;��Ə������~����~���0�m�	i��T|א����KC�A2�i�	q33dE�̐Ei�� 4��l	3 �s��Y���l4�QrFz��Ub�2���Tvi�B�>8���j�ʏ����̃j��g����}f��i�t�J�Ǥ���p"��`�a:�N�醙:C+Ԝ�kb�B��3Kx��f�S@��j��%|�V��pc	��C��S��#�0ߖA���� ���!�ږ_��o�L�rS�v��HA�y�)M��)�-��qd7���&�!�p
�7T@�a4��
�<q��O��"Q�g1��Z�Řz&hAe6F� 5" ��J"u�X+�lLK$,�۩�'�f����T��L:��jb�>��R-�H8+�ʔqx!��GP�9��a,���P�E�a�P�B�&��������}
K�)�,!3��Z�0�����hˌd��y� |{?�g�G��~�h������R����=;�L��k?x��"�x?tq�,���+���]�:|�-��.����O}���K�C�\�f��e��C���5E_}�觋�&�'��!��-�A�r?���c<��eTE��`7�Nc*�B�q'�w�*�E�1^~�nR�K�b�p��j��x#<`�ƛ�����q/�aFs�:���
�S�s-�-�'x�n%x#���,#xS�.�2��ܩ�T�?PK
    �\IE?��  �  6  org/sqlite/date/FastDatePrinter$CharacterLiteral.class  �      �      �R�n�@=�8qcL[B(�  IF���(R%��z�LW�]��X��a��Cb��Q�c;��jU!k�>ϙ{���?~�¦�*�סㆉ��2p�@G�6� S¡�������uz#
'�0����z���*ޕ〞�y2����SOg~"���d,�TŮ�K�v��	d�(fl�Q<�����D��$}J�E��t�S��e��*I�9s]Nә@���X�*��Fv�ݗ��d8�wRRN�d{{*��,�ۑ�e<��������iH>�-͓x̝(�=5��a4��� �X��K�Y�g�/����!��|���T�s�ˬ�K��������r"�8Z܄Ӈ�qƛhs� O#o��X�ä��!4~����o}������r������E]{�����ٌ] 
�AV�/.���_؄��r�@{_pXet�!p��%ҥ7�������WG՘���V�`i���Tr���+�Z��*�װJ٠��&V�Qީ� PK
    �\I�2�G  r  2  org/sqlite/date/FastDatePrinter$Iso8601_Rule.class  r      G      �U�OU�{wf�0,,"��P������d��V���;,S�:;�4>�w�/&Ƈn?����c�����F��D�x��Z6�̹�{�9�s~'w?���R#Z��\<+�Dc2�e��9n��0)�χpR�)d�8@���eLa: ܹ ��|g$�$�p(W,�f�G���¹����k�Ʒ���YC�V�����eW��K��h�JbZ�:�I9k릣�}w_�'���������מ-�s{����gM�� U4�3���?, ���t�%���\mcE��,��J����:��Ɛc�kf^3�1EG-�Ϫ���8���3A	�-ΚNi֪��A��>�@��@���M�,/X���E���6T��.:�r�����c����F:�R�e����\@�A7)Aɿ!�}�8��,S+��V5�BZ�\�j6�6t��pNC�%�/��Sz�H.%mZ�e����C<WQt��(]�г�3gZE5Nڕچf:SWJڦ�[��6ݼ�z9a�<$����a�!���0�#Z�%�Y��,�"��Y��ż�bX0�0#�s=!@�\X����3}
�!������*��|Fh
:�����ƃ���`ֻ���9=��
�Z�TҪվ��a��	z%�@@oL'�ޡNN��v���9�5��x����
�ѫ��.��S��=�?�ק�����@_��-�s��6�ۮW�d����	�1��'H�O�8�����qs��'�����QL���y`�@�M��kp�7s,�s0�ٗn��O��q��FcG��~̴��zn ��n8��Ww��a�c��,����A�e�D�4�"M[/�ナB�eo"�R�l��r�9�䔒�f#LE�#�V�"�ŽN�^���G�k匘���[�m�D�א�7hb�"¾C�q�z���1�~�(���WL��0�~����O����:��%��[�W�n�l�0�v��Q$�S�b�?�E��0�c!-Hg�����A���� � *��X�q��Yw���[h='n#rWC���U�3�n����S����n��]�2x��i����Al����(�PK
    �\I��   H  0  org/sqlite/date/FastDatePrinter$NumberRule.class  H      �       ��1kA�����ƈ����.ئ�"!�ү:'�����,�򣂫��7�{�����CC�V�&pG��z�f���ߖz�U�M�&ަ&y-�/��7AN���x�fLxj���8`�m���'tr�(��R�j uA�ދՔ�gq���Kmd�~��cGh��1]��ZײOA�<]�#�P
u�B��C%L%D�.P�<1d$��=PK
    �\I�ӥ�O  �  7  org/sqlite/date/FastDatePrinter$PaddedNumberField.class  �      O      �T]OA=��vaYJ��-��UZ��m��X�4�J�`��q�eu��ۭ1>�?�_|��Dk����G|�#��n����йw��9�̙�~���#�#�h�Ĥ��"��E�!o`
�ʎ8�cj8��:N�(�8����ұX�!Z_�K*��]۟�B�\�Xb�J��ە���e�]�U+��p��g�ﰨ��v�!� ,KZ����,���J�h�$��4�Z����}���埧d��]_z{��(���.��
��/��z��h��7��l�v�`*ҭ��<3A��ͦt�k�|�rO<yG����Ol�s�����o;��p�]xE�Al9�gؾ�J"��+���Ðޔ70:j�5ۧ�P8m�[�v-���Xl�������C��tH!�H���z�qdM8s^�]���QU6}�ᚈc�D:�M�`����8kb�L�0j�<.�g8��'Đ�qe���҆����\m��~�ё1��IS5I�Z��w����uO�!�)Ml~v1'�+�-�V�7����G�!��GH����2�^��F�$}1l��	up���;�t��> r���l�-�l�-��i�c�Ɲ�Qz/��O#�g1��"�簕�ǺX� �v'�e� =l�$p#L�1��h�'OQբ�7���$�T�_H�nCHtw�x�6�ĳ�IZ�u�@������/��_�En|]n���Ǳ��;��b���8�y>3�Խ@"�����S�^�}�u�;�~�T�)_IL�F��J��k_6|G�K0�u�p	��M��-��ۘ�x��	#�e�;%��.��.��L��&�����wD�7}��R4�l�a{p"tCNbY�O�3~PK
    �\I�{��   3  *  org/sqlite/date/FastDatePrinter$Rule.class  3      �       ��?OA���y�'"��4nbK'���D#�~��\��������2�Iab��ߛ?�_� �q^�,pF�KT��*�>�F�9�����ͪ&��b�ol��,5X_�4ۭ���o�:3e�p��#�\�MX��:!\�8�mZp��*���u�L|uV�l`��Ç���7�^��q�	�ߛ�v�V��?�r��A[�,=�Hz��uP��.zI�DNp���PK
    �\I�}��  �  3  org/sqlite/date/FastDatePrinter$StringLiteral.class  �            �R�n�@=�\��BHJ��@Zrik��"�T�j���M�M���ŗ~�����E���ET��B�����9;s<�~��	`�,��,,㑅�xbb�Ī���q��X0T�c~�Ž���mQ���d�ָn��H�9Wzb'�E���J���z<���]�#2̤��D����y"�(���#'|�(�9}�<�^��`��_�S��Ӵ�YFrL���F�C���f(���}������P[�}I�t��t��}gX�
I2Cu�����@te"C��~6�M%�M�l�Q3�fc&���҄a~R�n�X"��uob��҃��]�I AT&��t=(#՛am��\-��5��h�LڕD*�m7��&��ݴ����_a|&��}g�\���{���i6�ںE��V��sS�@���7�>�eLj��Q3�iN�D��v�w)[W�N	�����}��9�,�Y?�zqG3[��{���� 7鬐U@�7�l�?PK
    �\I��F�  �  /  org/sqlite/date/FastDatePrinter$TextField.class  �      �      �SKOQ��m���b���KAmK��o[0CҤ>"Xc\M�K�Nq:%� ��&nܘ&.�R4�ӿ�o0Q<w:.z��3��q:�^���eAAABI)��Hㄊqd�R0��4C�6c����J���M�`��+,��z�ԭjfֱ����a�Cw"�KA�����WC�`X�z�V��^2)-�˺Y�mC޽��Y0-4'V����,aO�z�!���v5�x`��Tt:f�s�����{t���ͷ��=a�p�U�Uu|�$	���"�E5}��}������K����$��\�!��!�Js~^��V��ffZ���v-���={u@��`��m�:[o�e1cH>����-�8�A����p}
.h��K
�r�T@K���۬o�E�aݯ�V�]g�A��OΘ��;%S[U�?�����:��ZCz�b�ɽ�G��C	�����JW�K�Jc��_z�A�]���H�%X*�
�J����R�6?����o�o��(�p�C�F��ܨ��8Ž��`ѝ��/�z���C������?���@�	�rO7�ǟ�,%� � �? �7��?b��0����%����T'x����".�<r#p�ҍ�~"�X���)iq�M���ؘd��������lۡ���+���6Ķl��0��6�u��9���pȵ�ד�I!z�	��PK
    �\Ig5�w�  �  8  org/sqlite/date/FastDatePrinter$TimeZoneDisplayKey.class  �      �      �TKOQ=���i�P���,A��B�|`� ���@X�bZ&tp���Ԥ;�Fw�4&ݘ&.�n�Iƨ߽-��~�~��;��>��r]�!�9�)yʈ�n�ȊhVEN�E�YT��*�Xes�Z1��G�k#S�,;s�]f����Mq�ɠ��բ!n�K�-��}dU,�1Cj�o��6�%w������[�y�\0���"�v���S�J�K����{l�gf�A۬TLg�6\פ�\��f����́Aǆ�z�^:V�3���Mh���%x`�m����{�mi��2to{F�Ֆq,ɑ�*O�%�-����$I��yR3l"okc��̋Y����w�+��WG}/'1���5�hnXbtߕ]�D��(h�Э!���A|4Lᶊ���WD�4�0�^%D$�?�Eޥ7�
�3��c4��s�o�OK���b	ii8ڞ�{�s�S�'0=u�H=���Ay��� �*g�du��Q� �B�1�x�y�	>�I>����k�E?� ����h	�$%n~�ƈ�B�A|�1 �bB�-�TL�BL<@��S*����Pz�Jd�9�-�;��ߤ�O��T>!Yi��6+&��ݒ�$�U=�\i��!��b�+�[�gZ�50.f�My�����������o�������:T�F��"��0�3��y<!��$�q��a3�Lh��QnI��Rh����I��~�S�Lc�l���X �� PK
    �\I�}�B  d  6  org/sqlite/date/FastDatePrinter$TimeZoneNameRule.class  d      B      �UIsA��i�0���`\▨l��qM��dQ0Vy��2
C�x�gx��ŋU&Z��&����c��<����}�}3|���+�	,��L;1������
�`�".����:�(y��5\�qC�MSz�ܮ��dH���"�u�f޷"����nY�!J®����v#_q�n�ôXkZ��"'-�r�2dR[W��|ܶe��X)�����u���l�r��Z�NU,��)�E�X�90rw��0�e�-���n̒mKg�):I���w�7-W�낎�q�IY��]�mOAh���0�al�w�)�d��(mY�w�AK�ipbuU��j�!������t�Nd���9�H"K�=���"�@-�����<4�W����ڳY��MP�-���:59c) ���rJ%3�3&��m"�=:n�����A�HbH�]�p\G��,�L�c�v�ۉ��x��b�����w-���C�_z*kD��e�#�/����D�>��Dܐi���k�}�����t��&�ݦ��'��nVx�j��ķT����cK;�T�?O5r#�)/&ٟET�g)C���}:ȇ#�����Ypb���N	�OE<���F��&�}��F�b��O`��:B��uh��6����p&�5�C�O�~D >������U��8@�?)�0�iGp�J*���QjP#��~;�t����o@'!��7kG���1}��	�2��r������x���8���B�i�wʎkی�A�jI�.�˄��Qn�<�eae)���
t��~�8�!�0N�(B�1��@�t�< !��9����.���'PK
    �\Ip`ڮ    8  org/sqlite/date/FastDatePrinter$TimeZoneNumberRule.class              �TKoU��}�q&�dj�4ͳ@
v��n(n�SC�<pp�P�		�d�L�	c;��YX�$�
$�MuH� ~
~A�8w�y��T,��3����Χ��߿�`�2Bx�*���!cJ�U�xU�k������H���3�E�;2���sMBV��y��!rBܐ��P`��拥k���j��+��%����kz�U]כ7[�Πdk5��15��-���z���a���Ĭf�Ӥ,4���7Ǐ'I1�<��/�;�e������5S7�5�����c�2j��f��WV"�<Sߠ�zs�~���.���e�\Ԛ�����eP󾲛\2����G�l�J���Z��b��#Y����赍R�!�mk�kqS�U�E���\omn�͔koن�h&]ך)њ��3<)�
�;}��CYꛛ�nԏo��j� Rը�l��E[+�wC��L�*��h�B.RHY�5���_K:/J*8����*�MܔPTP�-�r�D�ZT���$,+X�ۄ��^��w����Uk�&�?ID7�*8�ACBc�A=D�����	���vy�ݣ������Ñ#h��S��ux�G��iBo?��&S����hiz������Qָ��"D���3�"]�1Ď�-u������
��3�qu�)�g�rY���D"�0�D�g#��,��(>��ѻ5 ��Ω
n9�sr�h��i����)�N< �����}x�����$�"�������ƝN�:E���g��"i�Èt���>O�ǃ�~a�;�����0���NQ?�?û��X�_�߆���h0�F��^L�m�;��$��#_C����P�F��=�Q5��O�I�_�C�<��s�����T�om$}ѐ����h�F���S���0�?G�����.��0Ϳ�<���-��w�Ϳ�6�;��3`�� �Ar������1� �Ts� �$�c^"͇�H|�!F��!N�[�����;�l8��e�}��?!(t��?�ع���9��z�����-j⒳��8�l�C��#"�D�9,�� PK
    �\Il0s�  �  5  org/sqlite/date/FastDatePrinter$TwelveHourField.class  �      �      �S�NQ�n�С�@+����Z�ψ�1�M
!��m/ep:��� >����ğ���ԕ;5�ҍ1�{gR� i���s����3����� �຅.fЋK}�P41i�@IS*2mbքc�2CO�^�Ik%j�d;v��e��NGv����tzn(����,:�-2���`b�x�!}���p��)�pr��Xj7�?[u}_���R4Tmׅ�.W�I�7]��]{$�y�eWz��Cy���j#Э�N�(�*�f������^��-��Z[w�%v��	�鬆ؼml�`!�G��9K£t��5}�0rP%ԓ
�ܿphS;H!#9����?X��$F�TQ�Uj�.ˮ���Ŭ���Ŝ�>��)��lz��ژW�i���F�8���ީm�z�P���D�:�MI�F����%�*�fY<v[Q�!"
�ud@��gH�M_�AO�9FV)�V�5Xi�%R��KQ6(��=���)6g#G�u��h]j�	����v��u1���Xv��`1����	1+���A�zǞ��fڸ��P��var(�\�������>�9�y�]�b���F1��8�<)3I{��|��rL+O��W�5�h�=��RS�?���f,Ĺ]F��hk5�	]}��?D���i�66��� PK
    �\I#c	�  �  9  org/sqlite/date/FastDatePrinter$TwentyFourHourField.class  �      �      �S[O�@�f;l�n��U�"��r�
���A��M4BxvvwX��.v[�w���/�����L�%Qb���s���Ι�ǯo���9�Ρw�P4�`����EY2�b�5q����<�%���j2L�2��E�#;K�v�t;�|/�nC�V��1�B/�d8V���}�^����R��������z�L��DM)��������4ȣC��ｖA��܎�'�ʞ��r�SF�y�G�/;�ע���!�Q\�0��c4�ں�#q"\_Mw7"����@�I<�<��>��Pw���s��*���V0�á;~L
��ۍD��8N'2u���`�R�uY�Tn�y��J�g#�~㘠�����ol�ƚ�&1gb�a�?��0x&�i�H�#�ҿ1�N�+�)��+�,r����f.�C?ITEkHuM?�5�A�\#��=�U�
VZ���G�2��6(=�M�x/�)6�d�@�5Fyt[j�)���'dNa0|�bf�	��Xv��b1���1+���`�z6����f���T��ӧ0(���E�����1�f���)%X]��0����)3I��Yº�h��ӊ�RE;tf(͚}�˞te��p��g5���v�.��y���u�-��{�,˰���2F`�PK
    �\I��R  X  8  org/sqlite/date/FastDatePrinter$TwoDigitMonthField.class  X      R      �T]OA=��naY>EAA[���V���D��M*iH|s�ʐew���|!&�h>�K�;۵�6��{�sϽ3ٟ�� X���Ad3șH�	�L, ���2��42Xʠ�0P[�l�X��b�h|��d[Fo|/کJ���牠��0!ó����+#a�8MUFk�yH/A�"I��X����3h��-���h]zb���A�7]�L�}��[<��N�z�#)��#�G���kG;1W�
����k5|;_���v�׶7#�~���A���Dҵ+ܥp����3L_��N�`���̥yk*I�����)��������;�#�R�8y��ˊ��(ƨ)�ZX�ma
��,<�,���o��F�N�o4w�1�"�]ۻ�o�5�� ����˙�����qD�J���a�|4��4z�i����)�Ly]�Cڤ0A�z�кеc� ��a2�`��[	A1!H�?�ц�h'g��>r����С�:\X*�����������#&��'Djwwb�a��E���K�_��⍥�c�ϳ�BZ�}���}V�0G��[Y��o���]d�`�0���C
��{@�@'):Y�>�P?�ǆ�PK
    �\I�T�p�  �  9  org/sqlite/date/FastDatePrinter$TwoDigitNumberField.class  �      �      �S]OA=��]�K�(UPQK�l�#�4!�J���t;���w���O����_L�� ���G�Q���νw�s�ܙ���� pw�R9���+YWT0g��Z�9\�a�!�m(��9����}�temn���^[2�6�'��-�o��K�B��wK�*��`Z切a|�EoUu��w$���I�A )i���;v��UZ�mA���*���g�@Yf�l�p���RzSz���+st�!��'��f���4wž�]�u�M����m�/��V��"\J�rx�l+Zg�<n'8���Q8�cy#I3���X#Z8���D<c����P�S�K��ф��	�9\7�ɋ&&q>��&�����۸ð��2�V���+�P=	(xҏ�Cݠ����:R���5}�
ǑA0[��&�V�Z��a�p��3�
����Q�����ab�"Y����W����>���(�-p��H�.����&�l�B����c���	�|�J�� +F��0�x5��ۇ3��u������|�3R�HVd���%F��i&�Tc�,�"te��8��$��0�Tk��p�������>IxDR%⯑�o`�(�w��d�Y	�$B�2BySV��Q�1!����y���PK
    �\I%�vW  V  7  org/sqlite/date/FastDatePrinter$TwoDigitYearField.class  V      W      �T�NA=��n��UPAPPK[��-�4�HC��t;�!˶�n�/|�'��I�1���G�l�B@B�df�{Ϲg�L����?,c�Ds)̛H�	L<D>��̥i*�PL��0T�o5��+���;�-���)��U�<�W\"`X�u���re(��i��:���B��_�Xe0֤'��Z~a�A�tZ�a�&=Q�4���M�"�Z���6�����I��A(�PMx�p/⪒|��
���0���>?�˽���������W��^(]��]J���b4����!��#r��a���nUIr�G�`J��ƭ0�:=�R�1w������(ƨ)�ZX�ma�)�-,a�a���02c��_4��2����˞�n�u�� �����������qD̗�e�ҭL�b4&�4��I�����B+S��	�	diV��[��;\#��'!Q0\Ǎ��$�_hCE��g��r�����Сњ)K�1��V��y0�}��f��1��n�VĞ�mLQ��:���9�*�(N}C�<�'$��gX��1`5p3�=D9�5������s��WE�:��J����Z�d�TXTZ=��PK
    �\I�~j�  �  8  org/sqlite/date/FastDatePrinter$UnpaddedMonthField.class  �      �      �SmO�P~�ڭ�e�	*/��|�D�$K��q�^F�t���!����/��&� ��ܮ�����sO�y�������� �L���:b��CC^�
:����@zf�hY�P�PfHV7�[/6*����6�,a���`o���`T]Wx�����k-�Y�?9v J�e���+2�x�o�"�
Cb�v��9����fP+-K0�lWlt����<�Z���6�ly��j�g������j�m{!V��v[��V������C^r��,�*�����+�����N��
�ފ,$��3d��$3�`��!w%oU����!�������ۑ���D��뭎g�5[�GϵuAHa��t��f�d �	�᱆'�b�a��'f��C�T�fc_�C�:��8�v���Ai
�W�U9�����ҝ&�x�2w�L&�)���i
ߟ.�˸C?��~z3Rݕ8��M��Z��Io�숌Fh��J
�2�Q:� �!H�"�� ���NH�2v&3��� enB�B�@�8?���C=_�e2�����u�!� r�M���7��(Z�gs)�R�\������_�,�~ !���(Mu@�AB�ň�GF)�!���=�,&�kw�VQ�Ľ^K�d����������;
�����B�B��K�Ѥ��D�Y�0��PK
    �\I���a�  �  9  org/sqlite/date/FastDatePrinter$UnpaddedNumberField.class  �      �      �T�NQ����.�RZ�
(ʶEZA��xaM�&U� �z�=��e[w���/�#pÍ7&����P���+�8��B���lvwf��7�̜s>}�`+2☉��e\��L�*#����\�j�1c(1Dw+�04V%eE7u�.CX��6�Wni�a����ag�.�u^7Ȓ��������1�l�6C���&4?"�W��)���m[��R�e5��sCwDQ���p۹Oª����fNAYf�l�pIa;�.�ׄ�t�Bj�
���0��CQ���=^4��,�9�ڼ���ֲo�8�Q,s�ܹ��V�{���")A#�`:�!�3����7:ԬĚ���v�<y�ձ�����_͘w$���J�
�cI�&c���&n�p[�L�
�X���2���?�Ð?�x��8��H����]���p�]FC>�_4�j9�{&�g0$Z���=S*�\�jO0L�i��"�M���3�7�$YH�@������o!�&MB��I�H����q�+�6�{�9���	��F0`�y:��^u���E��a(�j��h��A�*�����H�"|�Hv�Kߑ�~xHS�w�M�z�I���t7U����]5����*dS��/�<�H6���}����!b�nސ�w��C�����7Ƥ#L�lH:�C��P�<TZS��4��2�)��.a��i���*�Pq�v-*�PK
    �\I�n  �1  %  org/sqlite/date/FastDatePrinter.class  �1            �Y{|\U������n�I��i�'i�l��-Ж�AӴiSҤ�IZ��$�d�f7�n���b}�O@��RA,�&�hE����Xğ��**X�߹{�f�l���~���y�̙�3�����I"�˧u.vSOwS'��4S�iJe�/MY6�s�γ����,��&7�h������|���x��I3_��\,M�4ݴ�	��-�����i"Wg�5�LVj�h?/Ϣ�x�εn*�:�r�^�.��y�Η����h7���A�FA�V���4���ލKn�y�Λ�t�p�f�/���M���n��}nZ�W�|��.�~���y��a�Y��[�T�A�pq���Ev!7_�;e2�I�!PD稛��2��I�ݴ�c�'�N��t�%��L�ݼG���W�{e����\�~�r����_��k����C:_�6����@6�?���d��ep��7�)"���Ο��SLyB�-�Hpy(��4��ɨ�D���p �u���ģ�͞�m]W8��g�6tu4c2��'����������hWl~��`��ifû���Ο����Cm�Ěh$�n��Ȕ��o
RƦ���ܵ���`kڜ�7��H��0�R��0dm�IX�g}"��Շ�X ��մb���)�ofr�@���B��`,�F6�-g��@X���HbS �tP��X���z�S�	��V��5���6�����X��q��L����8����Wv*ÁH[e�텸LGJL��]�P�25�-zG}�% <�mH�a��!�3��Z��UƯ�ꕭ4��xb9���&�e'��u�	�F��+�Pv0�Z��YM����iD[����X�RYc�k�r����H �Ñ�(�,���f�p����"����%�7d��p1�n�Fk��`~L}(�b6��b�M����I-��Ч�tQ`g�\	[�ΰ�TM�gRK�A�1�g}(�Yo:��65���3�ׂ!'F��i"G<�@�N��D����T:�xp��KJ�3���5c�֧ƻ��JѝAS$���-��@^���0�;1I-�_)�j�1���2P9bI��V��F7vk�'������x{4��\�v�;[{z̅��8��cmG�|\4e��EZ�{�w0)[�v!��tJ����p�����=��m�zCR,%Lyk]i��i�`f��n��@��]`�`؉e]�p+�A���`K"�?�.����8!jؑ�ƺxk���v��b�"���W���W��k�p��lӽ���C	8�ïm��-��Wv��3���FZ7D�ƟEg4n*u3Gu�<|d��*pv��aq�.��;�y����^�Oo�&O�x����#�ݩL�Y��X�-
7I�W��ZԖ��jz~���0���%��&�s�e�0�$�%�_ r���`��h�%��=���AO�Yؖ
����~*<�cK�hw_�	^�G���LJ��D{Jp�������� w,hM�f�d�E-u�ή�f|SB�o�96�=-�N�z�u� `�!3��E���%�:��l6`|��O��4AZ��iQI&qn���3)��EACI�8�á�vH�O�M�;%C��I0���������ٳg����J�Z�V��^���%X2?�,aәB����g�=��A��V�n�/�%�ݠ�2�(�!�����G:>���e:l�m�t!/<G�y�"�倰�c��^�V�o7�����i�Hs'����6�.���tD	d�y�_�0r�����~C/	t�4_e����DP�_5�cC+���!��Zꦼ�F,|<`�����JsL����QZ���L#�Tɡ�iϦ.��ձ��\�~�L�Β�|�CS��uJK��׋$���ˏ�E�|��2|t��P�	�}�RZ�:r�H��ՙB�L9��A�����wj�H}4�f�7��,���`cdg$�����j�T��px�����t~��oC"�7�����'z���ȑ�YtF��#���5�{|J�'�>� ��[�`��?4�%�;dy+R�r�ؓ�����
�l�O�{0�����4���:Bw��S��េ��{�,������F�W!֡
�%�
���[��"��7��оdMT>ҥ�?�����#��dF��ʈ�2}I�>��B�U踳�Ʃ ��5�9�)z3�P5Dp��ִ-Z<��t��|$ޚ!�0��VUof�����ǊX�̯J3ֆ���
����+DI�Bojy`JN.[�ë!1����츒�d�5W]���5+��FNT�Z��Q�7�nTǆ��U����0%��9�)E=��Aϟ1C�e3��M�r[C㶚��Ɔ����dPխo�&A����;+���Rp_�Y��a͗��7��dV��i�Ykv�Ѝd�5��$�"���g��6%�q��a}P��2�@�$0�2�ԧ�>X�'S������P�N�(�f���DV���إ{�YK����T�H#9D�)�r:p]�&\p�r	����
'֥Ua��5cաe�/|6���s~E�B�(B����n��6KJF]we��u;���ʹ��_v��M�&�$���e��}��>%_���T@����Mߜ6�ƟO�����(O
+�yR[�=�+��I�d����O����2��M���.���W0����~���T�q������8NNL����5�8���[(�s@,h���bş�C�����������أ�����
U����0����r����NP�7�}��z����Q�&��%����Q~��&�=A9L�w���/:Nc�U�du�h��/ĕ'��~\y!]
S���AH�7�j�q-���a07���8V������Z/�G0�!�]:_��oC
��،;����\"��>�6�Yg/���Q^S/�]S�C�h|U��h�U9ю���T�pD�	�o����l_�/�zS�[�e7�e���C�Uff��.0d��繕����C�yc|c�j�B� �L��V���ϟR����x;~M[�%��Mg9[0d܆�]��9h�`~f���S>l����1d����@MlR+zirUN7���8S�1�"����ϣ!]�&���CSe�1��Ayr�Q�Y��y��S�k�`
�4}��/��.W�����^�9�K�en�ߛmoX�������؃���{P.���ɭ�@�-pZL���N{������~{�^��6�YV�+����M)�zi�������>�#T"�]�l��Q����H�L��O�T�Ʉϣ�*�ю��*dt�1�%��/���[���v_�n*���9�����b��.���>����.�S��7����Z�C�Rշ�rN�B�6���3�GS.�W�:�=p��O'������To6�N�|x���8���P#=A���k��S�~@q�!��5�4�D��k�3����N��:����<zAO�VfҋJ�FYD/)���j���H�(��UX��+�OJ�^Sb�ge?�E��^W��7�O�ߔ��w��C�����Co)'�m�q:�<I�(?�~�4��+V��YU^e��:;���K%�RU�V��P�q�:�ǨŜ��q�:���٧��8u+�Wr���Ej�'�1����)�<M����x�z3�P���(�Շ�\}�+����E�+���,�_���	/�V
�RP�]lC+m�ц��PԆ����6tІ�6������m���H���mh���P����!�mC���:jC7P)��V�R g�Ƞ�z��Fͧ��}t��v�mC�ԃf�˖�d�<C}��Z��#��Èb�)X�)P��>�<;����JO!����a����Q�NO�i�z/�������Ǡ�E+��`�O���I
�����iF?�"C��u�)B�N���:^�;T�ӳ���=�~����E���y�T9�z~�G�k�_?�;��.��O5댬Fv���Fք|�G?CӰ�m�}G�M�� �ʳG�}$3���_��d6�h�B�DoZ.�����)�9�|��N��[}��m��r�����Is*|�Z�٧i�}�#�]&���}�A����/Txg�@Ū&�����y�.J���B#�^���t�R�~+�Z7i@�Msd8=��$�Y��n�s�rէ5V�ŋ;W�2FE0����K��Ki,/�B���\KKx��:�N�r���q=5�Z
�z
�F��f�ŗ�5��>�[�6��n�+�+H}z��Ns+����"��+����u�0�����\���x�:Ei?=O�2��7���M;�~�|\
�gz�~�=�G�ykH�g>BL�y��;ͬ��r��5t�<��!�`����q���R��<��8���+�<�SI����>��
�z�d�Ђ��hqSa/-9�G��@uS!B���I��{����t��Y|�y�)I��E�o͊G�ߙ��#f���\��=��d��@(%���ǩ�y�e�QMy-?��I��$L����C䕉�Z��UG�#~�}�X��nr��/����o_a�<�4������x���!�-�i������h�}���
����vz�RL��O�+�[J�\��~�%����t�_�U]4���~�q�f�A��\�b�l�UZyQɭi���C~$��G�.GDη���Ln>���ͳ���,\p����f���բ�
�r�|Y��mL/]�C�zh� �ܙ�5��o��7��Q�,�U�[���v��K�b<fb4�{-�"�7m	(�ۈ֔C����$px�;��A�L��b�I+2H��g���L	ַ,�����>�i��K�+Ġ���A�96�Kc� +SM�o[��U�&�Iº�ByB�)��L�)��Dr-��i�("i B���{��l0��~�v�F�[(�\�?%Y(�b�(������<8���ӎ��
�cn���Y^v�.W������*�?�žB%�G�zV��4�)^�6/~���G�b0������k�Wi��L�Ն���4�u��/K�;��W����d8�z�?�a�����?�0�L���m=�%p�M��C��i�H�������/W���C[�Ox���}��~��&�j]�@YJr�T�L���dZx�h�؊Zb9����~KQ٤f���p�Kq?�{aڻ��LJ~m����]i`k[����CQ�&�I� �l�L�@4?Q��,HRX�H��ݜ�A�E�Z�Qf�Ҕ��ͷ�)����&�.6�I�qp�;�+դ�@t)5i�'�Y��9&A�ǰ>���l6�=����{go���vl�Agj0�`=y�54AiH#X�c�pȄ�͘�b�gy��9�죶&aBT{�v�B�	�J��r8N�Y�p��\,p���\ƃ��N�7���(��%�vi�Tm����P[@K��i���dr�/�,�!�����Ǜ�T*@��&4�LA Y1=TŅ\�QDe���28~���<����I�0�p\8����2 7SӴ6M^N�l���S,yM���N7�.��"M^���Q�Aӏ����4�XΧ��ۨ��(ƺ��B���������~�b��G���_��Z���� �j�B��_�� ���?�~.������c�?��z�P��t�PK
    �\I]nX�V  �  .  org/sqlite/date/FormatCache$MultipartKey.class  �      V      ���oQǿo���"�bm,�CM,ijHHA5=ԋ��,l�vYLz4����K/&�_�Ɠ����ĘX��ņb<���0���̼O�� ����+Ș�1��	��t�����c�~Xo�Ǽ���v�~�m[�2�D��ZUo�f`kZ��:�
C*7&=�Aj'��ӵ��w����7]�L�=���w�?*Aˡo��8������u��_uy�gӿf��K�=�	������;<�r�eϏ��f���KU���M�k�͘f�\�z�;�A�-����[��qi~:"�u��[v�$FX����	Dtr�ˮ�h ��8#�4��2Ҕ3�P�S��t����n~ܾƭpYz:�	S���"$�e<��&�#�Fq����,Bz���Q.�
���7$�K�d�,��%��]Qש�fu�7_A*|�L�[(��%�G㧂q�ǅP��7|G9ݫ$�>�-�"�ţyII*3�1[L*��jZ��X&����kh�*O�b���B�a��`���_4�c� K@��&�KL�2�B:1�,Y�I��224DA�:$�D�4�9����2� ��O���ٰ�,��i��q�v�PK
    �\I�y#��  �  !  org/sqlite/date/FormatCache.class  �      �      �W�sg~�^iee�(N�DI7MeY����kp�8U�#���(]�kE�z�J+����+\�)	W�I8��0C�� ß�P���]벚�����x��x�k���ů ܅+A������6�P��XE��pPrgQû8D�4<�� t<���S�$��g��bx6����b���>$v��Ç��1|T�ǂ���5<��>�~,�)���>#���?�@+[N�`���%.S�m�-�T2K
����
����p�.9��LV�l�/��gRr3c�Ӧ��g�E���䬾L�Δ�E�v��+�1�Я�-��چS.�JzWF��l_�1+�}s��|q�p���&�O��R̃$��-�ξ��\n�ag��N1gg�t�@��9�
Zc�ӄq8?G�[Gs�9^^�5�SƬŝ��|ư��bN��M�9�#���SBXXw��~��z<|�dMg�ĺ]C�㑓��&����F3k`(���f�T��o�6T(���|�$CI�ЄH+�c��q�p�J囩BXR���Z�蘳"��w4��3ޕ��Ҏ�9�h���4~Z�7��ڞ)�ԣ��tTc(+x�VL�v̬Y�ŭ��R��#�,	�7aM
��b�UHb1K�^����.�m�����{5���]_���s��L=�G��땬ϣ67�)CT����%���U�b�S������F�9|.c�\��gsb�c�́�����Hr#L�5�&fϘ!/�Η�s$'פ䝂XǛp���7�����NA�y}x=+E3�4|A��%_ϯ�Hc�6V�/[ֱ|��+F*����B��D��5�6I�į��͖�؈�`񼆯鸀���5��8�!_�7t���Đ�o���-����Fap���:.�;:�wu�C�S���?�[(Xf��콞��rj�ϲ̬a��z��hg�2��9kN���|T@%��+#3���dT��#1�X�e�О��K��۱1�\"��y�`ȯ7���nL��&Y�InmR���Sc[t���=�Z2�cMX4˘-�����-���\�$�m*	[����¦Tw�V�y/�򕇯�=uůI��+0��R}#�6'l������7
Ӟ]��{6ly���@��F���w��(_�C�h�.� ��w�C��� �wa�����n�dM�ν����_�_E�LX[A�ϡ^����(>.��Hٍ�9��H��ρ���TX!��;��_
�,������2�+������lC[׀�H�C.{�9h�/��!������
�\K�A���^���W�����LkOzFM�g|���'��ϠF���/"��E|k�#ޓ�]ƶ��=��^@G�<�G�/A���0B�F$��q��#����Q��(��>LP�c<���q��E0�)X8�NJ��	Y~��0͡1b� KJ�D��D�ỗ��Rj����� -�3��X���ϥ#�8W�P�5�eLj�Ш��b_��I�X�=_^�,��3��!@\�jO"�^�vB��F�e�R���O`�g=������L*Fv�iid'A��FvJs[�L���vP�᫉�NϴqOJ���m�V=�^���﹊[��GEW��1������V�S��<S��T.\Q.�)WU)\�'9���=M��[@�KM�Do-.H-�.]E���^�݋��l�N�;8>�D�"�7�}�d��	����弗��ig2}	���?��^/w%U]��5�{�I\������ḻ�Gll�b���ѹ�}IU0)-SvW5e�K�&}��άb��
�:n[Ɓ�2n_���q-�^��=x
��u0��P���q���oY^_��c%�=��t�`��(�/�����?��ox����u��{?y��#�Vf�XV�Y�)�a|�yo��Q�E���^�\��P�� �R�'dn�2v��2d^χ���˿�uH��tK�R�o�!Q7���S�"�w5&$r}zg��b������1v��� PK
    �\I��W�h   y   "  org/sqlite/date/package-info.class  y       h       ;�o�>CvvVv6F���Ң�T�̜TF�������T�̼�|��ĲDF���t��̒T��D ����A �J?'1/]�?)+5������H�#3�db` PK
    �\I�E���  \  5  org/sqlite/javax/SQLiteConnectionPoolDataSource.class  \      �      ���n�@ƿm\;7�I�Pڦ����Ǡ(p�((G�1f+cہ>\	$��B̮��r���ݝo~3�6����O ���QǮX��а�a_�
�5ix��>��NjfgȠ��#�a���j���O޺g!ݬ:��C7��\\*��2��8	��S�3�>w?�����C��8�|/�q�:���n��q��}��Y.����/�P=�gؚ+cX�L���u#�]���CP�]�S�����/�!�p��̔z;t��d	�������8�a�L!C��M�/q2�޹/����o�	��Ųb`M��9^Wg2`�#
-���ð3�z9{pm�|ĆtBh0��a�^��^��_iI�6Ϳ&:C��߽�[�=(�GZ:=��(.Z�o�Y��:E`��-4hg�",�EX) '�Z��N�P%���P6sUA�U����ؠ�`�P�}4��+ԾNa���J�hh��Ew%�Y�j[�����}x��	�*�'y{�r:X[ؖ��M�-ɸ�PK
    �\I`0���  r  /  org/sqlite/javax/SQLitePooledConnection$1.class  r      �      �V�SW��V�\D�*�Հ`�[�Z�b����x�$+,lvq7A�V{�7{�Wm�:�>�cgJ�)>���������A�;�@@���ɹ|�w���|{����� ��wŨ�� Va��
�@�8��P~.FzJpG�pL�����$�,����rHHMz ���S
z�(G��Q	3���-�ܖ��b�����@�p[L���G���3�5ꢶ�qO�FJ��kC�p�s_����m�۲�xʰ�f�jXFj�@Cxާ�|-vBX5,}O:ӝ.-f�R��٭9��g�>隀�FN��������Z\�IzjXC� �u��R8bjVo�#�O��iG?e�i�S}v���l��$f��M�Hҭ�@u4�݋�<i�LJ�,-���ԙr�Wj"�2Ð�R�p\�&�@h��oËkR�Ksz���CE��=|v��)��I/R�esg�S)s^�':SZ|�]��`����ۉL�O 8�y�#�i����ːE��_����j�	V�(㒂�*���c��u8OS*^��+%�*.�5��9K!����������w���9�D7��*��e�������U|��T��|.�8���24�R��_	T䭳@y�j���x%��_�N	-��4W���&%��)vE�U\�y����oy��}�B�A`��,�֬��;3f�/�t.�u9VW�c��t�u�t��d���������
ò;)������p]�;��O�5���"O3�c3]�v��v�b3$j	e��S������3)���qN�d�)���x[�^��b���?�Iw�������+�T=G~��3�ݑN�-v2i�<'���c�f����L_�Gݒ'{�m�j,s��53ͼ(Cr�8%�����.]��ʖRz����j�Գ�����-K-����:��t��iǑ�H�iiW���Xn�7����Z�����B��q')�&���m�KJ�~�M��Q����s�Sx�9.�H� o%���¶��<�*�>(�7����W���
�[���1
��H.n 0�b.��_ῆUYb���FIU��\�O�8�o��`�Т��"���7�����bq��4k8L�⫨�oȊ5���6�GPAA��K���
�B��ҥ���.}�q,��=����T�F�أ�|2�*�x������0p�mu?y���˛I5|a��ͤ{s�W��<ߎ�`9��Y�/qދ.��� �q�߰j9���1~Q�����8n"�q�Қ�;��?<qIL��H��ph1%j��0�w_#������Óx
E\�������7ŽK^�{�����z�؂&�!�8�[%θz�C�\=��t:Pr�
v*h�P����*�	��)xAA��]
A*��$wK��P;A]�Dژ"���i �A��	����у����~�PK
    �\I���{�  �  -  org/sqlite/javax/SQLitePooledConnection.class  �      �      �U]WWݓ�LHA��T[�`M)(
��*vTl�}�$S;����o�S���Z�-����CTW�� �+++�뜳�>��?�����X�ЏIS"���W�pM�	\Ǎt�h�Ŝ�n��WqK�g�q[��Z^*U|��}�u-?瘕�U�vks�b�L'繮��Y5��8�J��
�M�-;V�w�J`����`;����c����k۾���1���s�P��������s�v�`^��ԉ�ҫ
b9�L���Z��-�,:<�3<�j����c��M�i��7�XِK��Ͳ�9V�H�%ǫ�4���Y����%U,1+;%kKhWTܣʆ4��-�9l��-�W0�j#K�R�S��І���z�U������헬E[d��ɉ�"�����Fuo���+�taX���q�*��a`T�E������X�#�N�;����y x4�͚]���TQб��:V���	�\j��?�Y.�����wrS͊Í�7���l���	���{�y��%��,�I6`��EMV��A5R�"�(�YUjVET��j�B��l���7%�e���%S�z.�Kn%0��-�Z�����ь��Vy�����a�ǳ� ��ILl�Y����H�����f?�B1ћ|d�=9�D�Rv��΢�'#��'�x����P2oY��b��=t��&�9��Hs��^d�h�NAW��r%�+��:P&\��Yh�d^��=�Dl���G�\t��Y1�{��E��^�<�O%*��!�q*�%IL2�k<�N�\�Gc��ܔuZ�{���]�����"%�+��1����6�!c�A4�
�W�b ���oѽ�����޿��S��V��-G�y�\$��Q�>D)
%y��e|\+Q��?A#6��dk��hR���?��^���|deE>i���	�?���E��zDԀ��B��PK
    �\IȚ��\  �  &  org/sqlite/jdbc3/JDBC3Connection.class  �      \      �WYx��G�-Y�I"�N� y�$NNB��
�,%�@뎥�2A��QJ
J]�B7 @e-k�� )K��ҝ�t��ׇ��o����F�1v���;�������շ^x	���{�� �Ç�-��0=�� >����~6� {|!��x��H��p��>ւ/�K��8~"�'��S!<��ϰ��V×�8³!̰}'���g���${|%����X��!��+��*�F��&��7C�V��;A|W@�.�w��Л> ��UC)��e5_�4Y5�Q�V���TC.�ڠ��͊�[l��r%I-Ƴ������f8�.�\�5C����=�rA�(���XuzR�r�d�f��r^*�4�}[�c��8;]֊q�ڒb�������Ρ��uɲ��yC)�D�_�Jf�)�$�I��B|tz3�./W$�e#)R�\�4���{:<�ì�k;N#ȑr� M*d�!��NѴ��RLP�O?Zo�R��Q�b9f��4I�%n~J/�$6�}����|P.�V�UdB��fwM�I-Y��JFU#E��7�m��%I�7�l�j��V���0���li�,aE��BF-��'����s��>&�����J6�ʆ4D~pF�4�L�MMJ�\[f�u�A9{yZ�y^!�
���(��,iWH�J�:'��T_�[�TOJ��h�}��QN���*�6���'�x���q*��5�ʥ�$% �*�ɒ!S:��
��A[m��-��Rs,5k:yBӓf�XA��h�hrE��T"'�?�Ϙ ����	p��H�6/!������`TA�-���c�.S��ĺ���<2M����W�'̗K)�@廊z@�㔭(k����!��Hy��/������y$5frm���t�K��boH�րʏ�ŚL5����b^����i��jO���s�<��L�é��$&�$��\A�D�f�U-/�PX�_�:���@�^@��Oq&0��0��**j���j���Ī�ٸ�P@}��+����z�R)k�.&ә��Dr�x63��H�&����T��JF�vF�}�@��k<q�hB$�&����� n���.R׋���JY5�V�L��XTl�Sn<1�M$s���Dvx<�H��%���EI-4,�'�&v��Ls�C��l��dCT�+%��r!�ag?��'�i�3[���nJJ*۟�O�9ϵ��TI*�Ҕ!k��әSR����$��w�h@�R��8�5�չ�of\=����~��ys`������/�F����e�;/�,XǠ��"kJkMyq���Zj'��#0@�l���BY�Ef��r1k���E�9���H�z��7��mF��]\�;����=û2���x��@�,� �����M���՟�Ƈ�É��(�|<�NoO$/s�RGU����C��)-�V
8ӱ%OFǓ�pn��7m'w����k2�6,5<oc��$�i��Y�����@��^��R|vPf�+�M2�j�,�3c���s�c�,M��H�kǢI�������9H3� �J���I
_���K;P�gk6�x�K�]��|tRY�i��56���HQ�6X�&�¥L4:��SB'���y��MK�ڞJ�n<$;c)��~�f�N�cg��������ϓ�b�F�`����W���^��۷����������Y�Ҽ�y��\NM;Ў�H_=�6�"��.� �a��4���l%�Kh�� ��!a�^O_ls���glma.��$D�)b�49��#iam�/&�İ���֐@�Cu��l�M⤝����E��	j?I��!x)F,�w��KVW��h;���h�Z^f|�9ʝ����Bx�X��tv
;	�2.)�7(M�W�h�9�p�3�������6��,�#���\�:�.��~!�uxk42��#X�ǧ�i�"f`O׳׭<�l��.���&;�H� ƈ�.
�8y.�|Ķ|���,oF@lmmi0>C�~+z~�3�y,f<\�����]�w��8��哭�O��|��u�f�n�q��,��y���C�8�o<�`��'l���E�Z>\�#�nkT��,WZ�ۻ(�Kk��ј{f��)��C�aG�mG;��������J�w�L� w�����O_o��M�np(�ي|�xa
�D޲��J<���O�*,@� ����	nr`�<0��hm�0ZX]P�:ݍ�$t����h��^+65�������d��f#]v�cXN�+���>��.��z�N';��H�ݤ�0�pE�^����<��v$��ߖB�/�/�{*A\�@�d���lʇ��Zɋ���eD��� )x�x�ΖGp&%�G�p$9��h�4}*��X0�'I�S��i��q:J��-��J5䳒>��Gz����������λ���DQ�M4�/Y��z�Vz!�Ds�������4�J�n讒5P��%XO�w[O�M�[�k��j���Y��|������zW������b��X�l�nn	]G#�K�!K�մ҄Z�=��\�zs��[�4�mMaK��F���w�ҹ��|<��fp�۾7N��Z#N��p��ʹ7����l7�?�o��m;�qcc�9�M�����7�}��oY���~?>0��9�7�[�"���\�� ���I����nB=ti�<��{�;0�sO�4o<k/"����<��2�H������#�Z�*,�ba	V�ٺ��u�D���
]�0>R?��(�nQ��`�_߆b�	�:9�99��9�N���Hς(����s!�}<��r�[�7ۏ��v�6���y��޹;Yk����CX�~������.Ng�Ã�3�8�] ���i�8m N�ӦS�t>iq�E����g�4a�# Ξ�)��}�i�)>�1�į���_�/�ն�PK
    �\I���l�    =  org/sqlite/jdbc3/JDBC3DatabaseMetaData$PrimaryKeyFinder.class        �      �Wkp���-�J�&'H�c=,����y�±�I(f-_˛H��j����W�R�~�HRJ�L$JR�t&�L�2����i���ig�p�ʎY0�����s�����|��������� ���x�</���`7/{$��B��� �1?b���xYL�0�G�S~M؋}Mȣ�� �Ňb�aQ���e�`%�oڏ><����EF~ɏG���_a�U���p�_�8$�u��h�߫Гy��%��0s|�}�@��⾴�/̒��=uI�)�ԶZ �oٹdi�pTr��x�+y_Ow��G'MzI(G�=��c���I`�53-V�	��~�T�ra\�#s^YY=?���g� �W@t';�l�PUl�1�I[��tr�zEFz�1��A�(��L���j�̥�����y�TRDq�5��V+����X^��d�w��
�t��.]u7�J�3��n	f��E�97�ߠ\K|S�[�Q�%�-�2�UEǰ8�2��jb�Gc��$�+	o���<8l���jpPo����̦Q�tiX��5$q��ոCC'ﾃA���Hɼ�;���*pC��w���k���Dح�I�����(���!_�QD4�?����'�$����*�I]xҶ
�j��
z�Qv� e^���AeGYl,�q�DR��Ӥ;�&��)*���&D(��E^�38J�7R��rVٜp|�ix�$^а�)K~��l��~�c^b�O�*����Rï�5_��s���aNZlӯ��1۠�7�-km�4����=�_����n��s��^��@��	��,.���+5>W���*F�l�`����L �4c���9S.�zާ�ʜ��%�P��F��w�*����
�٬*�\Mcp�5���BB*~i�&K��C�o��k�yY[Q��p�\K׎�9��`�2��ȭ745��eG�(+{�^���1մ�&h7�پ���-=c��GF�e�M�Aݡ>��hP�祷�e��g�]�k���)�V���̪9S�&��[��+oζ�E�&���ّ����`��[*R�"�bUw�Ptvfj�3'��e�����?E�b��歒B�>L��⡇�/����4���f��tj���y'�������?��!�g���ȋ'�8o�"�$*�U ���5�w����3�4U��O�K�e	-,=�����t�Es�g:�[��#q˘zy��Z��<�B�V-�~�$jD��C�5���R���06�g��#���z*XY�������"I {��ʖp�!�N �
n�'�%^2GInz.a��7�f�ico���a��4�Ρ��/�+�9�ȮƐ���f��f�o\�k�����Xɰzj��!'(�Ç|��忆�6�⣂�ޔ��"���cg�{є�%�/$�cH��2|�8)^FL�*΋?!�a.P\o����xW����\p�f=�/%d2��2�er-n���.ףW��'7 #7aT�%7�D�a��!ك�V����G������>9 �ʌX)�D����;ŃrT8r�xD����Q�ǥ.N�q�����|H\"�������2������Q��n���O���6�^.ulĽ����}�6���͈g�F5�"݁�юF���$Iǭ�c�$�q�{�!���x�?�j��^{$>���⿤*�v+�|����s{V�A�R4��6n�}���3�J0� ۆ�0{j��:�T��:���]���|PK
    �\I�H�61  ��  ,  org/sqlite/jdbc3/JDBC3DatabaseMetaData.class  ��      61      �}y`[����Cϲ|D��(N ��� 	qB�9�	��Ql%Q"KF�s@���@�܅/�i)�aG��r��(��@K��r�R�ߙw�I^'������{�f�3;;;;3���}�� s�Ӽ����K����<<����L�˽<���
�7h�Q�M�3�7k���+	�J�6zl'F_E���|Q���Qt_���1����X���N�]��xD��5�A�5��M߬�Az�A�q�$�w/���xR�)*��yߢ�^���4�]��S��v�>�'z�I�{~2QN��N��J��4~�ƿ��h���P�gj�,��l��H��P��z������f~��/���~��������D�j�2����/��O5~�Ư��U^���L㻨�k�j�_��k=|�"�t��Ư���4~==ݠ�5~�f�ߢ�[5~����$?�.wPU?����w�=t�[��x�������ܿ���@�j�7��}8�?������c���'���'5��Ɵ��3V����5���Q��i�y����5�'����5�g����W5���_����/S�oi�m��U���;������{_����?5������5���?��'�T�i���\�����/�K�|E�Z�^	xZ��G�H�$M�5I�$U�<^|�ñH^Mʧ�O�
�^�IEt/֤at�k�pM*ѤRM�I#5i�&4i�&�Ѥ��4�Z�פЊ�2z��I�~�&D�It��I�T�*�*i��դ)hn�TM��I�=�/���*�D�K�4i�&�Ѥ��t�&��H��M:��-Ԥ*�/�H�=ҡ�[�ўpr�����h�;�d���dm,�JER�ؾ�%�jj.�24l
o	��KGc3���m3[��t$_d5]U�Z���z������vZkGC�����A��Ec��ym��p�/a0?�v���7�lK'����P<�2$-A&��+:���u�-�����&���M9��A����x4��AYEC"�af�X4�ٶ�o�	�GW:��/�\�@�MtGh�x���g]$�^C��!���
'��l���(*1���u]sg^WS;�.���"��t��8��c0n��0(�IgFVTzA�̬�#���OxS"�*�L���2�S�;�K�&�If����ÑN��nmS�ڎ'���X�=��º��T"6���m5�8�'?�5D�������%64�{"�5����&��;!Y�P|Y2��[��AINE�Ƕ�훓�l�}iNE[$��0��i�,�5W��d*�t
i6�E�h��Z���H7�g���5��-z|�f�ֵ1�v64�nK�ӑ�H<mыs�)��.��E��>x��H2w�Z#)���Hzy"�^E#G�aZ��e��^Sj�4q��}]ib��-kw�C#9�m���uEzM=�l�+�����wp[:�k��	-�{6-�-ҋ�t�fa��I�]�6��{�)�-Nvm4FLu�iأ��F�G�G#ɕ}�t�h`t�:Bw�5��6�A7IF��������%nO�|:�4K�ў�-� �H�hm`�O����Q�X�D�:�E�a��L�D��aXiX�Q=����-vQ����X�����(Ź��B�iD�q�d��x���TƾC�X_w�&�XG���~Ӻux�i�F�Z"��nX��?�q���GS�,V��I��C��s���E����Z���&b}��D�	��]q:���=�D���`� ����̥_����*��<���~6�!�Q"�����h*��6kB��rk�QdՔ$����,�Cd��)�Q$��a��/c�8%e9��Mwg51��m���v�����ޡ��+�R}��	k,m��������n�qa��d��j2�n��Z8'Oc�l��p��g�����q�tJj�=��(�X�/��k�鮍��L�Ȧ�⤓�kǣ�}V4҃Hf�!�Ƀa^�%��*�a��������U��g��HW\u,N���(SGo�kB��+W[�L�aAM'���L�d2�C�t���;��!)h�U]��S��ݹz��.N�P͚����Eׯ�$ў��Z�`Cr�)���m�h�c��C���,)��׃�,���<KYɈ�bt�g:����96DѱF���ЪOD��O&�eU,���Ep@*�`�ř��ɡ�D�'��V��S�7g��AV���'1����.=Ѩw�����6G�؈��m����AՂo�߈�H�7i�č�$�ЭUk�,�ɴ*��g�UMs�݂)BO$m:)�����y��� F
���J&R)+8N�Ek"[�1�1vj�I߲��F^��v�C�]%2��DJ_j�n#��G�Ц�b\�]}���]h�e]�fY�#��p�v�O�¶��DzQV�D[�F�&����v������]���{N۶�uV�HZj�5l�gK"ӽ�����L��v�!J�0����\K�"�-�Jg��Ňb��/l,@J]�7�˴�!� �Q�C̸��R�o�;��|g=WS���s�LXJ٩���ǉl����Yt��E[w��R��4����� }L�>/�ű��M{96A{fa#����Ҙ#g���o)T��!�PR]	=�F��#������u@��D�%�K�kW#ՃTcgA%c�z��H�4=�����>k�AO��@�E1D�&�z¶�3�K[�U��T�D(��nKI�HbY�Y㤭�j��zG���ĺ��:}��I�a�	;����k��1���CCH}��v�"�LC�S<���;�D�=鑖x��=�a~�qdP��󈞙t��;�3��?X-��K�.8|==������n؉�1a��W~f۝2vǙM$4|��e��fV��l��.ty�wP�A�"�"�u��n&{����1&��f��H���lpZ���v$��s�F�
[��#��"��rhY���XX���B�4��Z4��m���V'���D�9\����p���S���>eȤw��ʇE�YiL�҅ƌ��z�j���cT\s���"8^���o�HK=R��L{&�>3n���[����860|��P��O|{�y�PNSEB+���������'m4�U!:�ԏ�J
�����X�!ךX�R7և�#�ۛLlC�����ɘ���y�&����a�n�����h��p��mX���΄F?!��5C�y�g�M�`z�3<�YD,w~��ą!f������c�Б[]{�ۛ�Q��\�Q!#0�ǜ�&�t2g���JF���c���r���rtl ���dN�4��a<f&v���6��x8��`K��0��:wu���Y�f1X���J�~^��m�2�g�&׼�����o���b�,Gs�A[�3�Cy�}ɮ%���;�A����Ǌ�0�c^Ա��x�1`İ����=
�Hu>)��@:�$�D���`�tg����EQ���|R=��c��2[M���r����?��mK�i��Se�+����iٔ�������ː���[sHu��՝�4��P�БNt�6�X��YZjo�Л:;[Z�����u�#�����`cu늶�^��
j�S �I��q�5�z���\�U���e��3Uͭu�&���-�jn�Ԅ�:K�V�l����yY.Y�wu.�=�CsGkm0#Y�N��f-�I˥�G:�'�`��~�h�-g�u��q57t46�sgB�g����>�:HGCMjK[�����`���D�.�FI9F��r�T'
��&.k�njon�!-ZZC�B�e��I՛Q'�7�y� �o@� 52����,0�	I�|R��̠�+>hd�<{����Cwg�4��ks&s���2�dZ��ʠ븹Q��Z��/r�k�A+u X�9dǲ�������D��7����.t�eN�n�ı�4�ʛ���l��&�V^�!����JL�L�������� ̗U`�k����X� V���}� >�'�`0�VJ�>�MjG%��Z����L�ytF1�(�xY^�:�\�עk�Val��VKG`�T�g�ea�	ٷ�h�Ik0���0�c�JGb�b���@��[>�]؄� �Z�� �^�)�Ϙ�C1=:&c
�b���45)���!�Yϔ�qZ:GK���dh�h���LF����TEW�W�f��'C�)���X�}���:	2���I��۞����9��0C91�SX������ә��	�2gq2�Pi{3ԇ#��J$#3�W���>�1{��������r�ß�V�4sԘ9���Q���9˗�l�l�l�sخ7��g��>��+�k:ۂ+��ͥ��r��i�I�6m����`Ik����C����&�j_c���ޡxV%t���e����.q�0T qL݂oyB1*�c�I������
���0%O�SY����P��r;wZn�f��X؜�t�.J�=�+��n5ŕ�MU����X�]�ۘkuFqV��P]gO8�{l�-Љc١e�[,�V|���'E�#|�z�}�i�GZꓢ�b[�M��G�e�qE7�;7G�w�E�e3+�50x�u���bR�w�˚c�ojZY��擟��Wm�洃�3��F|����KO>ƙ��W%�^���އj���|�b�^\hv���$�GRd%�����Tt�R�V�VnH'��)K(Řr�g�	DWj6\��Ls˧㮮 ���؇^2�a��9Vv'͊���7y٫�|n�<��x45ÌI�9����c-���Fn��{��BD�9C�YP}�A��N~Cw�`��qYkS*��E3�4Õ�	<z)��3�e{� \l��3�xL8���dYl�ͅ�^P^�đF���XYu-�r#Åd��V��V�m���lkoն�h��	�]pT�:�;2 ey���ɢ8�q�?��'������)��ù�h�ѹ���!T
�~$C�&e���O+K�V�ϵ7�m��ʹn�5}hm��'ؤ�T/:vg���v��k����.l3nz3�$��ciVJ���'m��2X����~�QL�:���yx�m�Y��A����D5�l�)7�1�؋M�{��}�	�/��o��-�͵���֜��!���L��M�I��^��q��*ԖuĐ��F���^�<+��R>����i�m�~v����8��0�>��H���Ġ��%ؚ�pt5��:��:@3��ΐsXd*r�:�ĺ��;QA���}8�OG0ObP�M'g���VsOFYe�6{���}N��}�O������a��6Դ��r�`m�`S����$�cMG��-�9� y����^�&��b��te�f=4����`�QzOrڅ�:�|Z9ж�\��A;TC��hZ�ɴ3�3�d+���D�!���'�y>^��x��p��Tw�֬�_C�?T���Y����,zmk�������F:��v���x؆6l�x��������f.�-��)X�I�ʡ��v���߲���uruG{sg�	�o69,��9���֍��PcGc���#����E�`�g�t�˙�I�S�l�44��G$sf�:X�d��:��p�P�PәV�jEGEv��s�jf���ni��ZK�h�d����7g�����-�(փ<N�RN��*-��i$�S�.�N����dbk���R�ʦD�l{$]�x�C5^���v�L����O=cJ�iGMssC�)>�{�ɘ�"�N>w���� u��bM��U؎�掚u��h)z����vy8��1܋i��j��S���L�6���̩�heј�;�fϘ�6��$6�FYצ�V̘rX��Ԕ��� �(��>��V5�$#�����TWC��5���iS-.>�3�!%�*f`b5�Nvw����7�;^��I9��7�9�?g��_��F��5b�xe��=��m�}��ŝM,�n��C��d�'�j�%I���t;?�*�5����Z�����w_�m���t���%�޵�>�5~_�
��4�>Қ�J���xd[���:</�	Wd������<�9-���U�[Y�D�������G�K'�R0��lE��jC<}o����I�GI��(�i�h��(�ч���P,A}�b}Z�9M{2L��U
�5�W7��_��"}T
?��/6�Oxd$������u5ٿx�����Ȟ��oy<é&���f-A�%��D������6�/Ġ 뷳(��y�d�4��O�O�A�����wab�O�v䘹-�gK8�i^O��ja��7덓#-�ӫ��`t�t`�>�ܔ�⺝_�	��6�+	'����V�*�3��^�K�}8���޾�/oL�����CC�(O�/� ����"Kc�m�~g�}4�c2�9S��������@�/R�e>>-��P�L��[t��^� �`i�ъ�" �T̆ї&�φ��f�3ޕ)���f���2���h`�a�����i&���� �Hn#GFJ��B���H99O���X�F*��Z!r��>"����&R*�r�+PɆ�u��#���s��"ǻ@�"p��"�\ �B���ȉ.�;��] (D��c!r��%B�d�+��r�k��
���J�ۄ�).�w�S] "��@>&DNw�|F�����9��!r����9��=!r���6���h���m�P�C�P�Ba?h���8�g�,#�9�����"!��!��x�`!y����\h����/Z*�V	��бB�"�0z��X -ʅNB�����\�l��-tZ�=D��an��0!t�h�Z��(�ָ����n�G	�uC-�a��u�%t1�Q��ֳe�su�W�\>��籭Bd�E�'	���@�.D�p�<[�l`�&r>�p!�ǖ�BR��5So������c�}�L8�Vc����ϛ��vYc"���2�ȻAֻ�L�L
��ҁex�R�*��'�d���B��1jO�ok\X���cG�����8�����c����]���~x�ǧ����b}|)��c���޿Ur���E�Ä�.�QBd��Bd�r���r����`!r��"!2�Y#Dnra	!!r��>[�Ș�j!���!2�".�1!�ׅnSB�q.�<~d�D.�I�<EG�����=��X�ȧυg���b��
�[]�y����B�v�^-D��+!��[��.ƹG�<�E��'���Q!�{.�|Z�<��9!���Y�����y��B�i.�
������B��]�9 D�`�HI"�p�,"��qJ%B�.�c�ȳ\ '
�g�g��#�YB�9.���s] ��?v�
���m�y��>ۄ�\ �"/�c��)j��&�w�&}p�xC&�Q�Ď�%�"3ʖ��)�Z�4�R�\bo(7�4�Q��a�cg�o���~B=X|�t���|L��Ĝ�6�C��m�e.ԺE���q�<Q����4!�.�g	�W�@�/D^�y�y��UB��\ w��\ o"�y�y�wp�y��CB�.�}\����;!��*\a�Bߘbm�E��c��E�c�t.B���s��ׄ"���B��.��"o������~NMnt1	��~��喹y3"��Jr�y�y_u���t
���S�P<�8�G���;��h{`��m�(�x"C��C�ld.l-���r���xv;��^�K�^�K�n@��,��ٝ�`ga�j
�� �P�Q��P0#�Ybpp-�]8��^���E,�=Bݍ�E��8�hBg��sP��Jw����,�<~d:
-��)�0��f��N8�J	(��~���H��r]&�e2]��R����|�Uy���r��ҶF�Om�ҦL�6=��ô*O���3����{`��<�gVyYU>�{'���Fn�<�;/�0���|{�`D�K��&�` _1�M�E�|�Q*�kFi�2�(�%�b��~������K�K!��F �WE���?d7h��~XXU�����aQ?,��<��ٷ�[�#��[�0'Q%��갃��AiA?T�k��R-�����c�z4_o=N	���eR�IZN�=
���!�.Q��4�����
$� ����
�����"Rh�ݠ����w4af�o7L�*�mVJ͊�fD(���<{aM�ޮ�J��o��FPU�]��U�����+I���t�RѲ�� ��@���e��������ah�;؇|��8~/G�>���|�N���P͗�5�|,��7A3_Ï�gc��h�őY���V��`�����
��.�9�@>	�'�y'T˧�J���V���π^�L�.�;�s��\�%�7����xH���/��K�%�'�|)�K�>�
_�W2��e��ݬD�%�(_�*���|�v�|[!��Z���*�N��b)y�)��Γ�aW�����س���9���|�P~�}&�e_ɏr.��{�'x��$!?���{�AH�D���C���3|��;�����y��G�R~�������Xބ�ҏ�rZ~�o�_�ɯ��7�E�_t���=l�5��Bx�U���TO���,����0x�c�A/�g%H}K�����R\d�`;����^,��v�{�=^���o��+��	�$h|%z���X������,w�%�]b�t�Xz�p�Xz��%������+.���з�h;]�؛�_E�9�@#�ʞ�	�{��^p��E�a��3��P8d���^~�Q�e0�]cgD.e����FJJ���(J�?Lt��`�{��J�����Eye g�t�`0�!��[1�l �g_z�8�{5d�3R����=��sm(D�'+R��^7"%[�4kvM
ѣ���7�G!��]?��ٌd�t�?�tɫ�2�,���fy]�$O.����A1�҃j>M�c���T>��+�Ozl?i�sp���w�k�B��L%�	c�a��,�?�V��?����`��o8G6>_j5Fj���f�����L5v�7�Tc{K_;TzK�^�+�T�'���z�艈�ȗ��w���i�)f��S�uz�&�(E®<
�Ev�����>�
;�;��;�"���|�Ї���=��iA� ͋5��5S��	�d���+�F
���m��=��Q=�+��h�٤?�Y�N�6Wi���Ҽ���]P_�w�U�?��6l����(�y��YFie$	=O�c��2���)Y��~��H�WF�_c�1P���Y�88D��2�V&@H9�P&C�R��JتL�s��p�2v#�e������u�By�*�����l�A�����}����M�_��Z�r�Lw��u�CD���T� ��	>ҝz��"����5�[S��4�0͐^�ǔN�^��w��i�0�|htN�4_({����?�Hx��$:�T�7�g���EaY�S�~H��=�UaZ�I4ZI%q���� P��"����6@%�ʪ�io��.�l�̳wC)�Ҙf_�
��w��gUEր��,<�g�;8���/��pcX`�ށ��>̹/#O�)�?��E�C������R�
L�OĄ�H��MwR���ӟ�4ߤ������)x�v�i�����4��v�'�����(�4�5�g�C�pFf"U�S�q�Y�p4���L>gZ���ޟ1m�i����C�0)�Q��Pd��Ŕ�{�$|iU�n�$W��+�ƙ��Wo���}P������%
W�y��L�M3�#��c!��k�V�ڭ��i?�i�ٴ�v�.�i�b�]b�~b�.�i����G�������n�\?%�t�
������5C^��2��k{�<����qk��/�+�ވ���x?�o�=��Ě$��i~2?�����x������=�5I�"���X��s9z�z���s6@���ܬ(+�NiE���J�����M9
��;�c��X�FYO(�i��U��%%�(�ue����}%�)	ƕ^V�$�x%�&([�Te+[�lg��l�r�Tv��r";E9�]�|�]����Wv�g�S٫x[9�}�|�(gp��C^���g*?����B�|�X��/W.�ʥ|�r?F��oR~��<�\��X2֟���a��X��S��7(������j��r^������)���/%M�N��J��\/�)7HG(7J1�&�d�f�L���ʭү�ۤ��;�ە~���w�q�*��g�7�`�> �ا�3�8[������)�sڎ��i��%?����/0r�5\a�շ2�|��ȃ�y��}�qj'�ʾ�7!g�Il@߬`$�"��:#ba�k͈%=gE,�i΍�%=bF�j�J.��N���(����r��n�㏰1z<�r��@t����פ*X�5L�#�Ra�K�l��
vzf�1��5�0rz��%��b7ƫ��I{�?c��%u��Wp0�w&�x��(��ք�nu��+�=��7�^�p���|�5�gp\��GA��c]X����G
�2��ܠ틣9��9.��l0�?����43���Z������o�zF�֏�ܥ���ÑV��}���,Hq�����k����<�Q��[������j#��J٬��5μ#��-��k��R�~�U�m�P�Z�L��	�f�  �����ـl��z������=��a��9�4���ha�)��UUA����q�j*�T#�~�9��3��K��k>]g�x�ӯ�r�N�$�o�x#$*܄�
7cA��-X�P����o��6}G��|��&T�Z��;7F�p	\�dl�~�0�?�����0Jy�)�����p����'�Cy
�)O�z�H*�K���2�9�\y�V^��ыЯ��(���W�U�5xGy>Rހ/�7S�b~�ol���P�eӕ��<�l��[���mR>d[��ؙ���?a�+��k��؍ʿٽ����?�E����_���%�X����
W�^�2=�����P��R��&�T�w�(=���G�����/����|6��
��^�X*���}{���u:7�
�X2�%��R����+����!R�Q<O����K�:�J�d/�?��8
JS�ĵ< !�	۰�	m�&���������b�U��3D�}�U����讂}B�Bhٛ�;���O�;������r٫��0/�������i��a ������~ �U�w���T����ʛ�%�8��F���r��kW�[��!����v�����g}�����pnB��:k��=6{HI�H����>Y���~x���܃Y�~CY�*���l��DU�{Ǉ�1�fw�1�3́�X(�/�!��A�	٫�L��|8@�I��O͇Qj�j1LW��X��D-�.u$��Q�E���h�B���`�:�V��yu��N�w����Z	��SW��Bu:�3�a�,R�V�`֧�c���٥�v���ݡV�����~�P��0��Z����1�m�.>WJ���O�,+���pLb}��VZ�^� >�%�����}>k��#��,�\�X2�b�d�`�X�X�0M��R�ލ�'|C_�*�����Q�I}�jc��h�-OOg��Fu���ΐi�%��F{>���x ^�*e�^�zJ�_h�4��}�Ѝ�mz���Ny7�\�ҽ����}�8gy���W�{�c�G�c�ǰ���R=<�
(QW�5�p�j��YYl�Jy�`���K4�`G�`G�`Ɵ�b�$w!�X�	Bq��yB�q�	�ـ�lDq6��x�.g�P�'mq���y�hBqR(N���݈s�P��mq���y�hBqNFqNAqN�.ę@�_�Q��X���
�����'��yͳ�A�Z����[�ߑo�=]�@�?��9ʎ��|��B�__��2~�8��Ţ��\����B+����*6�E/S�/�-Jլ&��l��+X�����(ʠS�
��@Vυ��y0I=f��\�B8D�U/��՟@�z)�^[�+`�z%\���ԟ�/T�,G��u�K��^[��ڪ��V����I,�+N&�%��I]�#�3L6^�-D_�����e ��q�m�T��K�����KD�f`��e��zT���ވ���o�O��f��%E�-�zS�r��[�Wu	^!�%�+9��614{Ի�^_�q����}���������R�ٽ����Ѭ�_����6��.�������XnOc�=���'9��	>e(�;U��������	���(�'(��ߍg�&|M�[�7uq�B4�8��1q����r|:�av��R~�{��5��o�<y����x�#/��g!���pךV04�B��:��a�c�Ы�U���Ճj�O���}�5��Sp��5�o1yv��q~=�d���k|?��p��i��_Hl\�����B,F��@��4n�s�w�g�w�4~����> g��v�sT���ߗ������a�y�6�y+���w\��J��?���%g=~�d=~��O�>���f�����,����e⇼4y1ˇ�(eLT��le>,U@�r�,��08NY
[=#��H8�3N�������R����)�|_�/PK
    �\I+�R�  i*  -  org/sqlite/jdbc3/JDBC3PreparedStatement.class  i*      �      �Y	|�y��=4�et $@H�c�\��aqI�jw�V�����m�+u��m9Nj�ne�8�Ԭcns�q�&i�:���m��MR;��7����쯶5��{������w��+�x�*����t�~䧃��r<~"�맷�1��x��O?�_��1aČ	v��[a���~��21���'8�Ť_<f)����+��q��g+\����>���\���|�9�A<ţI<*��O�9 >+��OA�M�~j��^�v^�p��Vr�`
*��Ok�UP��]�?��V�W�i�x��S�x���^��Z?m�;�:�Qx�n��\]ٍ
o��]���ͼE���9
o�Sw�x�xw�)��b����{���
�P�.��ͱD,s'���dj�#}_<��:���J&Z$K&:�N�τ;���p�@&Kw�b�Q���/���dG��ԁ�P���d$?N�ķA�dFbi�+Щ�PdMǮ��К})m,�Ң�pF��N,�@������Ɣ -R��\D|���ĵpj_8�2Z
w��C��i�lF��G�*�C���𘡹j���j�q���-:`;��t6�Є����hؐ���G���Ld�ɕb�sԢ�ޡS0kk�����n-�	g�L�XE�X7ۺ.��&2Lu�x8�ރ1�ͽ-N���L�k������/u�%�]��Id��fvK�P)�Ebi�>���
��c�=�x\�\_,=NhQ]�}����zGEZ�tǆ{ 1�,h��GÙ�����3�xps�Yd@�G`3���p�{<���H�=���M�e�&G;{[�v�Q���<����L��	g�b�%��+��Z�a�B�Ƶ�p��ҵr�Vx'�\Z�A"�0���P�3v��]�H,���`"���I~!2�D��.os���q.���j��b|z�5���r�z�Yy��푼=:�x2������@�M�D��@�K&�%e�dۥS��`����`v�K��j]=���ǜ�q
�yN�R/���A�|G.�-��:0�L�VH򀮕��]+��5`
� �"����Yε��t�\i��E���'O�E�С�I�3!DqD�2�T�RR�.eE��("�lN\8� I=��H��t��E��g6�w�� �pJ�wGD��:M��b�vpA���l4�����ә���(�%]r�:M0�:��	o2�9ݬ��^�M e !���¼"�+�
� �Z��4�xb��NOaO�6V��+i��P�Ê��BDt����. E�W�t���}���� �ʞ'�Pp��#3����Nt��(:���TD�)���ai+U:L�����*��}*�
�Qy/�Sy?%T����|P�����X7H��|��������.$Mj�@"�	��L6��K��o�|�p�u:�ΐ��8��R�eU>.���YL�{U>���3�ƺv��=�єC]���]�8���@��Vy�#��O1�ٞJ%S���(�W��@�,r��H2��4�hKh��L쌆r�rT$�9U�$S�<����J�I���}X���j�ͺ��7Q�iz�`R/bb�Y5M�EL�O��&��i�ZJL���LP�*=K��O�D!2�ʣ�H���1�rEA�~�)��8��'+��i:]��Q�U��I���b��!��C�U�8��ΕE8ZUB<��E�,f��e�Y
'tgG'S��@$_ߌ�j��T ���ڦ��{N�q�X}�(e2�.��F��25��x@�(D��)8t~��u���Z8#ɔ��Áo�)���!���?2�EN��౮萨.v��n�oǒ1X�5��+�1����Ӣo�%Ҝwȸe��͢"�Bwk�k�)�h\�IѸz�8�w���z{���d�Gw��<]i����XF�Y�d<;�0�/������B�.��Ľ�//8�xk쏧!�1�C16�����e���W��x���= :c(U.��!�F�jE:0�J�7��G�!Bܺ�{���ի�d���&�=E�,o={O�ʽ�*X$$Q��{|w,��5\��iKG1�,ͅ[��QꐞK�O(������Q���:\7;�m�\�A�M^�P21x�A:D�u��\4��^r�_"%��u���.:��o�&*��t���F�cR�B��^b9:Aapa��� }X'��s�
>Gn�yr�=��T6�W��DK񼝪i��r���\+�F'�_�4���#�4T�a��AI��,G�.��Q�)�I�/`�[j� ��A^;͢�G+��V�
Zc�f���0���Z��������u�U<JW�r��j�����i�f_45\B><7A�fh���������Z���M�,���
�<E�=���1�無g����Vs��.�?�S�����C��w ����f��M���b��K���Z`֝�,��X(q�)Z"�ޑ�hn��W�%�y�\g�5Q�.�6�49N���K��mp��ЯZ���.���F)!�9^��S0[J�� ��o�:Ϳh@�$�Z6�kHd��<����r��.�"6ĬEH�C�(m�ۊ/�����h�n,y���0�3�)��3˦���]��n�y�8�)�Mg�8�s4nR�^�	y�-��o
Ygqy�2��p�2\��_*��˘���w� ��[�x�[&o!�A��[���-d�
Ҭ.���AW�~��-��2����n�5�MM�����$)�9j�Q�t���"b�%K�15�14���>p��k!�,u+�k�Я�Kn�<����e]�c��&xE�_��U�ܷ�oO۵�}{V��h�ᶋ�<rf1f6y��ȅK�{�AZ-�D�TV�.D����ET�/�㫨/��E��;��MZEߒF�D@	}�O�	-Ȝb��\z�> k�Zs���}��� ���1�\�7 ���=X�Mx�~A�~�>l�~@`Τ��Q���m��`k�-�p�t�2�&r�?AʿR=}W�%�*.0Oi�T�%GBYw>�W��S��	a>8IS�n��$?�^���g��LP�	�3@�X&փ�%d,.0}Y��
-�͟�fP�;�#�1����Ǣ�bS�Ŧ2�Me�lp�4�����`Cc�G�Q�-F ���#U&v��]�ÿ��,1������j�1�xQ���hhb9�V�fh�(��lm���D1@��� � �*�����>D�8�Jq����)Z�SG<ׂSi�T�8��yʆ�G��&�W_)pZ�>m8��i*g҆�4=��>�8E8�gi	8YΟП:������r�	gE	8l8Ϛ��ͭG}#Bp�a��j�s��Ȓg�� �ytc6��6Z"���t 1����0�\�O�P�:6JrҊ��MrM�˴f�����iM��>Ow�h�$����T��0&��h��gL~���s�)?y�����m�O>�ɕ_D�$=��v��{��X�.o�ѝ�M���V�A|-���uB��5G�r�5I�v[��;4!��B9�4���j"�V��6�Q7�r���vj�❴�{��M��G�:�{�!ޏ��O����0����+|���G�|�����C>A?��r����F�M{��8h�����<���6���b~cccU��������b���;�������_�M��IX1�**[��y�f�3C��Y	�Vg+	J�>��� ��RZx ����_��Kt��p �+��[�5�n�e=h�v:x������<���w���ޛ���ue����z����]�'o|/� ����L�R���B}X��fO����}x�h��)_2���f#�0⇨�?@��Aj�)����(���F��{��Ҭ~$�rZA/ӟC�jZJA��֣��,,Õy}�hM�M��r~Aꠥ�XB��S�B��+?�z}U��(�_d�
6�U�����8�'oy"_����ȫ�ץ��� x�9Y����.�����.ɖ���T�-_���5t�%�2��K���3��\J��*���`�k6[��II�| �+���f��[�mj�q�T�?�]�~���*J×,wK��G����t��k�_^���{*�"�o�S�C�`��8/t:pͶ�5��zMý�a����mg��u�ѯ� ��m����D��ߵ��}��o� ��l������o� ��E�l�5�u�I���Q��-�wXE���A�臥|�d�#�_�|�d�qz��.W��[����PK
    �\I*���  aL  %  org/sqlite/jdbc3/JDBC3ResultSet.class  aL      �      �;x���3�3�LB�d!!�wHB���E��I@@�.�%Y������b-U[+U�Vl�^��{�T�j��Z����ڧ}`o��[[���j�33;���&{��;�������}�����|�q �������x?���=�?�G�<x?Ű�I��=���V��ߪ�m|��*��Ï���|�/��˝|�|ޅw{���Fv/��S�߹�*��h�C��T�*~���/+� ?<��q���|HŇ��<G�2��	�����*��ƗS���
>�x;CW�L�y�_�$wӃO��|���"|N�o��m��;�����wy�x�ǰ���0���w��Ѽ��O�S���/?��i��ė_���/�u�/�R�el��T�5?��(�[l����w|�����H]p�ܹs.�������<l�Q�ט�?��?+���op�x�����,�7%����Wn�MŷY��(�w�U�=Ϫ����xN�
T�P��
Y.U�U��BUE�*<��W���U�b�*�TQ�
�*ƪ��>ZY����#����牉����T1��U1����eq$��b��T�,�T���KQ��W�$��+sׯ�����ɽ����Qd��W�f/ܫ�؄�<v��������9�X�j���Z�7H��Z5|���ZU�U�<<I.!�3wu�X����8O��4�o��־�s�����f���}�����pdn<�:8wC �ţ��G7�wt"���[:Zַ#�W����J�����x��ĥ�p247���6ҥ#H�zC���ٛ��XW�0�������=�xg`O� ��X0������ɞpa��=�s�554.�J�G��$�*'��I�ɣЀ���v5�"��Q_��~$�ۑ�����g� `��t����6l��Є"��u�D�$�8�В��m�>�rZ��`0ԗǢĒ$r���ۨ'A��'�(ݡd硾��I$h��:��t�/'��H{�+[t��c����ئp<���.��p�~/)�5� B
��^��p���p�l��	c�J�D�U�2Z�M�m�]F�/$��#$�5���B�po��ˈ<C>��d�ܡ.�X�C�3�au,NC-QѸ��.�́HH�)�"Te�[��<LT,	����eQ<���D�CzJ-�1Rp_��!ĳ�S1l,���P�TYC
��I�.��@�2�/�m�	�ARd��v�7�]�AN�Vk��`2��c���8������Z���ٖ�S
C�Y�b6��H(��/�����! ���sW�96Y#������dB�0-;�%g��y,�X��HfMYT�d�vu$�\���YF�6\���1��PKk,�m �e���X��'7�vd�a�m<򘔮�c���K��p�0�a��\4oEY�@Y�Lͤ�no��0b�X�ũѕ������=5�"0Է~�>����g��/�_��iM�t�0�%G�,ʁ��?�������ʌv�Oö�QzJ����.j5{]��s|h$�k%�c��$�<+��iz!SC�H�� G�z�o�	X8��3w%�)��9uh\k`O��j�@4�l$j5I7�+� �)\�6��W(b{B�L�W��E��]�`�@�
�@�;��8��%v�M�(��)
R����(lϤ�}`O�7`У;�(ƣ'�'r��CB2��Ms Hc �E�d��1�� �iɒp�)����P�Жx8i�1�_�G#4F':H���O��pw4ԥ�c� �p{��i
EBI�O-�D(�?qצ>N�P��?D98w�R���P#\���0ľ������]:��:c=k'��C&-���Ek�^�ڢ��[T��D�[tA����Ra���R>6җ�vi�)���7��DBo'�����h_���
����ʌS5��F�J����dM�M/�ky�/��4����2�\+�w�8�P}�	 ��*
L���i��� ��M��h̟������/���D�`�ш�0Ѥ�f�L��&��e-_Z�:^��(�BM��2E�i�]���&�"��vx,��F8Mv��e����49��O�c{�{(ft%�Kcd���͝�kw�^�qK��&W��&���b�]���5��X�(��{�"�+���Tl�I*�+���)��$H��ۗ�PB�J�Ͷ����=�(54�P�.���e9\��0���5�)�L������� �!LL��\��sX�մ*��&�h�(4�ѥ�����4�P�Q\j��|2ȴ�I��vE�а}��)v)b�&.E�ѰZy���U%i���Q_ ��u�]:Ɛث�nѣ��اa7Rk?!ѫ�(.��~L1��&�ĥ��r��t\IJ�~=�2���H�.&���а �j8�5��I��Ll�p*N�pδsiVEÑ2����EZ�^�y8�/u��v� �`\��i9���q�}[���=�j����b�������&>���u8[�4lgU֯om�o�����:_dr$d���}kK{'������V�)ӕ�t7�����ܢM�-kڛ����7z��;)��|�l��I�+tm^Ӽ��o[sS˦6����B����Zix�����/��Mm�[(���y�ku��z��׸�~c}c'�u���o��l���uɍ��)4)��7c��E<��Rۭn����N��vG�4_�N$|�����WQ���G�M\���QMd�׈kiJ���V�ߡ�X�����5�	���z�b�IR<ϝ�o�wT|J7��4q��t��R �܂P>Գ���X�R�P�h>�G����M�?%{�C�T��Q$�!&k���U�ܾkG��*��[�m�\��r;*k�.ؑ�$����;U;Ș4�Wz�<�!ї����_�L;�L4�#��s}_��7tf�§>-$�?J]=t ��,�#R�5�Х��H��;JTrYE�?Еq�L ����#)>��i�f�Y&'��e��gJ1�w�
h�7����aOo��F��It��]�S�M˳��v�>�8����O�B}��]�\����GI�	|�	���3m^�8%z��u��rbwR/�]��t�*�70���=����^>b!eEI
v6��M�i�H��J�ݶ��C�q�;Sq>i���Hh��ݔͣ��t�~n�ΐ*1���^c����v���
�����<��eI�������Q5��TB�17�-Ѷp$�)�D���X������"a6�"����o����l[U���܃��A
a���ok��я��$��x+3h!�0�~�cr6z��*ܨ��\�SF�B���g*���Cr3:�F0qx�����a��<�GX`������6]�$�U�H�����R�U�䳷6��im�Xkm�l���dl���fV��G\�Q'�Dތ[^���Ru���Ƥ̗��F00��!X�W�I۷���7#7�Oo�8��U��֚�Ҹ+�Xo��k!gx�"O���[����\Pk"gp��]�~1ȼ�����J��]U}�!j	���B�������g�������F��ާ>��3�̯��U������PkA�VVT=�����ܨ��1Ъ�+�KA8"���~y
ԭ� o�	�x�A#$���.�Px�|C��	y�U�YDk%�l�Dq]��B�.�y:�U4�3��p�f}��%�������K��A�@>c��Y@��.��e��4N����_t6��b��pIU�Q(�'�0�j+��K�� ���"������G����G`� �_Q�%���t\f�������4�k)MLG\R>eҀ%��w��A��$��$������U0�`4�j��h��A��A����WC�M�GLY5��ߐ�P�P>��Ə=u��O�o�w�1���A=��k�Y�u�}��7�c���e���E��;�mh\м
0�\O0�^*��P�1�+��}Pe���dj$�
�$jp?�Mӫ*�����M}��~r/�'j[�eb��GKlDD��4_�8]dr���K�1k�b����V30�'��ݦi�cl��.(`>���'����+�P��q1��b���B��-�z�#��&
�P��A�����kl\�+��U(�Wa�7,�-&fv��cPh8Y�n�-P���ױ��X4ҝ'�廳��ņ�0��@��B+R׀ߌcvK���g�be�_x�ĵ�r��p}/�o�x+�oy����Q����n��(�-�Uѽx��T5�(���O�$�(�o���o���U���j�?3�֜�����\I\c��$k�Q�0��@t |���H|_��'��I2�oZYc��;�w="Ϸ�a>ev7�w)YCq4�[��Y���4��S��q� Tw��y��y�=f��c� ΙX��^�B�&��HL�S�?�a.�0��d1���^�4�ӹ�Χ|&�z30Sp���ɯ=s�2yن��B\`R��X�F�<'�Ws&W�Lo`]nJZ�%}�So�P*J%�2��:߉�o9��jb]��#\ZNY�{d�S���X�K2P�`^6�kXQΙj����5L?���s�j��=ω՛3�Xh����pj���~��W�k��N�N6a�m5f,~���t�����x��5VRk�C��-s���>i�I�?�����%c��U��<����zl'�o/���a9�w�a'N�]8zpDq��l�k��*��"�����w�Xg��%�S� ��<ܧ��;�!ұ�H?D�,������Y�J��m���w�	��q��5�b�IhigI�Q�z��#/���9,�2y$1S��Дs��B�V�C�����˨`�Z"�����R�"X�K`��V\I�^1��˱>�Mp���Bx[u�$�m���ƃ0]]2�(��"8k�d)�%S��q8��Z��%� ��f8TRj9��;��AX�t�άN9�}ʬ�N�I�7�d@�]G�7�Yh�M��29�/0��X n����U�`�>��Y����A(Ð��9)sl�-�ۤS21[����H��'�X&�Y�� 7>�`0A&��6
j-
jGb���C/z���93览3j��Ȓx$�,�,�Q]��z}�TO��8*�M_v�9g����lTw8�˙�83ci�i� �ι��������z΄VR�U�K��ぜ�[�U٨����h�TWS��'�
�r�6���Za�h����#�
���
_�Z�q���Z�)���Z�J^�Q��<�
����
�8�_[+l�V�l�
[��
Y�l�
�s�6�
���
?�Z��T+�D���^&q�B��o�V�-�
��Z�5�^�Z�y�P���|�b�����Y��N����<���p�m�9�v�9ץ;�ќs{j��s{�.�'���S�.Q=bDE1�	�*J���9�L�1��Lͳ��$�8��Co��w?}���ətۈ�=k1�UԖ�n��A�9�.��p)��)�/���d1<b:�3a�����b.\)���D\'�b)|_,��t��WZN��9�K!g,'=cs�|p{�g��y� ���p��h��K�Ѿ%���t�]��K�<�K��Ŵ!2�#{��,����h���:����v��K`�-wB>��|�S��?]�c����;!j�Տ6�������q��z`w��`��e�։M�!.&���Nr�ݤ�=��`.�e�8Z|�9T!(ςOV߅<ͅ	,Ϧ����嬸x>� � ��d���8/���q%^`RUc��y�6S?D�U����Qp4XG�զ�mo1���(io�<�9)�k�#ql�D�?'�/�\����כ��X�o��!�_�/�[�k�<q^�k�Wl�̞V%3b"=���E�x�p�D�e�Zk�� L��9��@�"P�@`���2H��&����|*˫���墫K������.L	@�ԈZx#��_e��
�.P+h�~ě���<�T���eܾ4�A�R����{y��C��x?�^�n��&y�L�;�r��T�p��\���	tx�N�h
-��wx?�4�5)�{��mb�z�M-|]
��M��FS)V^�B<!������d
���GSc��
�\t��S)�:T��h-���K��B��ɸċ0]����ӰT�Dy���.�P�5��+�_��ʨ��U�U��x��[ğ�N�:�+ހo�-8)�
_������=q~&އӔ _�~'��䂷$7�-y%�S%'J8I*�YR1VK%x���UR)����"in��1(MİT�i
���ai^-��OH��F�o���h��R�J-��ވ��˫	�al���hL~�+����Q,&c��Xx�D�ԊE���/��̽�r�T��*?7��?&>7��?�N��-[�P`��a�m>�,��
�ZJ�Y�a�*9�{�^s�{�q�����_-U �ni1x�%����xi9L�V���*�.5�.�	�j�Z,�x����&�|��z����W|�>�H6}�$�ъxwӝ%PgI`��p̒�1(�e�c>+���N��Q�1�cޥ���b�����6�'YD�YD�YD�؈���}�%��X��Ej��6馸���<\-�����]b�_�:_�
��w��J��P*]uR �.��:���-V�MVJ`��/�Ro�B�tf7YJx��l>K-%�KW!%�.�q��PX&˦>캘J�A�G���.zI1(��`��)�%��YH� /n�-��fXl-��Zjih��-"�,,&~Ҙ����P�ۑ���9�Э�Hu"]�s��f�~�Y��U¿�{t�u�c��L��tY�Q�Be�Be�o�ǯJ_s��
��\�8}M�G�"�Jk�f[��Z�8S;��:�����a6�����$'��rƶ+ھ�3��9��p��.Ɂ���-�mO�mO�=�3�`��������?x�.��4�Fh�/��
����؛�WF�!�Ϥ̍���S�UU���p�3��1�ø�U�.e���
L��`E������[����]TP��+��{i�����{��+X�����.���]T�+�/��~)v�k���)v�u	�0��4�AWL7_���.���|�.�z��c}��_��s�ϙ\E]�\�b����~��W���b�����D�G3���0������"���'��J�D�8Z�m4|n���WKK	��B�	ܞ@@�h�TN,�S�	�WS�s�]>���)>u�)*���7*�{�[#IԬ�+�$7�r�|�)�I��-Jk�"�]�I�A����P-#,�\(��C�HV`���A9n��>�N�^xL����8xA.���xE��7�I��<ey*��q�<gʳ�Z����l\&u�Y
� a�\�C�ы��*b[��
��e�p��cT�U����7���G-� Q��Zn2����@&��b��$���B���n�`?��ч��2�@Nƃ+��ҩ
�Kx9��a?���NS�?Oᇨ5N���P^|.�+�5��{�Jj��І��5eX�WQk���΀�>ӡP��(x���#!��HIú��Z�L]�(r�s$�������a��:���xk �s����iƓ�y:XQ���'��uƴ՜�'���o�)m��ϻ��Q�G��|�.�1�B(���+�xQ�����;XdU�>{(.�x�iƥ�?P�}�$<�����~����~?�H8�\|Tq�ۈ�k9��u�PK
    �\I��e+I  -  %  org/sqlite/jdbc3/JDBC3Savepoint.class  -      I      �R�o�P�n�u��1'�t
8WOf�D�.\JH�K���b)���4qq1�W�(���Ñ�pϽ=�;�w������� �P"���#��:n���>�q9y�l30��o�}�!�v��.�t�#k�cZ�c��'�e�O	�S�u�Jv��մ�ʨ�4�����j����cz�Ӥ�}k2��t�����r��l��KEM۴\J唫��b�c�3�B-�ryj:X��2�i[C����
(�˯)��z��+}��q@d�=rZ�K�k:��ۡG!!���&AB�@ک���gڳz�uU����i��\���-WġIE�#1���
r��D^HnΓ��l�%�ɀ��-6�P,���8�{#�z��^�f�������u|��������W8��� 6  �yF�2��F��V��ҩJ��H�X!}��.��B)1�q^ Q]���)���!�$�O���S�a|��+�c�D���$'ߛ�� ��):��ŧ�]����>���xr�J���:��a����4n�%�/l���4|�%ִK�!z��	�[�H/hd�7i�vJ"v�o�w�PK
    �\I�}=�/  �  4  org/sqlite/jdbc3/JDBC3Statement$BackupObserver.class  �      /      �S�nA���º�m��R�T�V��@c��HL���:,S\\vqv!��6&� >��얈�lv��;ߜ�����O �x�"��)d��Ě���u�U��M((���Ȑxf9���!Z,0��nG0,�#^�m!_�M����>��
�3濷<��7?Ͷ'�HH��8B�m�y��;�+���Ѷ|��:m���ܫ�+-���/�0PeH�ە£�x������s"�tX��;t|���)^X�K���q*.(��p�ٿXO7;�� )oPd2��
��NWo�{����P��`G�=�*�h��
2�Ϸ9�6��1])��Za����s\j�O5��s�4�e#�X��/-�o�R�>riR�p|�@����y̰Rl�����t_�3O��ϩՓ�q6Z=2�άZ�͢��Ò�vhs���_�ϐ�Ύy$��U�'��� Yi:IF2���s�Hk"ta�V�4�Ȑ$�<.~GyQ��/�d���F�'��c��8A�+�	�6�5����c�@[�J�-�+�E�V_��iIl"Mk
�QJ�� PK
    �\I���  _"  %  org/sqlite/jdbc3/JDBC3Statement.class  _"      �      �W	|�u�{hV�с��$X@�"	��l�m$��%��r�0�`�jW���(����c�js8�!����6Iq�lC���I��N['M��M��I�������fg!�*���������{���^z�
����� ^��]�b��+aN/Ȇ������rt�*G_	㫸$w/��U�k���~C��������a��O��w�����OC�3ٿ&���?�/�����^�{ߗ�~ G%G?�-G��o���ɕ��͏�����
���go����_�T����?���7��{�!�����W]����ߒ��ȋ���_We��d�Vo�BBTa����/��l�<&*�Pi"DR�R6ᐨR���jE��l�b��c[�Mݸ_7��TJ7z��i�@źD*�Y/����]�d"�w�;��7ͳ�L"�Z��>�@o:��$R����nl׆�\�HǴ�}���sg1�9� �y^�#���ʮ�}zWe��>��2ky4FF��E �%�&)��M5)�jc��ƣ1}L%�ЁDJK&��uE?�ǲ�fEF������:�5�1��k��&=��B�lrK?�QD-�F<�f��IK�P����M��j�x���Z����ެn��v ���k�ٵM7��̐.uSi	=��������j�뎱�6���ԜI[dMۺ�J����#���:JpPϸ�����9�_o:��X�"Ő�o�2�C���=}�a��x6����k<L����	�ȫ�Y
D��!A	��,K8^Ap�=�
�e��zL=ӛ5̴�E����*J�S3R�EGj�
JrΎԮ�(�����Zt���+bZ*���jy�r��Q=���j��@�_jG1u>�8��yiP;�-������T;j�Ҧ���Y/��,^��ܤSq��,�
���N�%�k�0K�D\��g��Uh�����i��`��m�0-7�m�NĨ�CQ=��a��x��]�d\N�یܝ��c�z1m4cژ~����IcH>���*��*����jS�9���X�1�Xx�X:���_���)UB�$=�,�j7�4���o?�l&m�qL��G�o�פ9������P:k��M	��
�2y[�6�b��W�8�b��b&�*b�*D�*nM*���*�SD�*ZD�*��YU�E�SqI	�2�5���#�D�i݌�ҙ��g�F*�AU�п}㾾�[6��' ��y]2���+櫸�b�Uц� T�P,R�b�=�g�]�-i�Z|����GK�T�Ѯ�ѩ��xA�D���-�,�&�RU��
<���8��U*>!Vӗ��"֨�fqK��m&)q��}��I��aE>;�z��X|yC6��놔b/�����9�\U��d������zq�*ngC�ݡ�]�va�*6H���|��m�d�͚�ȰY�Y�����*6��1E����������"&�N��aX��晔~P�$��U���I�ħ��iI�Nq�@[���O�hÚ��M�U|���	|F��8%�P2H��%-�����]iD��G�Fª��NQ����{��MA���0[<͊��ʛx�!*؎q�Q
Mg�LG9A!C?�����a�h굋�ٓ�a%6��PO�bd���.Μ?�m�;�Y�a��t�1z�Љ���^,��]��� ��e�{�������r��\��ek&�ђ��
���g#�M�F��h�uK���U;��o�y�"a�e,mٕ9w3?Av4�/f�<�l���S�8y��ʦ����;�D�N�i�]pخ�BVOZV��Z�{�h����Qn�q���R3m<�c�i��V��e�,�����e�J�ajW�
m����N^z��[j����u��B��v�N;3ZzT>�L�OZ
P�J��Fv�6m��'�]�mȚ���,ZPF�U�U<;T�x��H�Ǐ�-�K�%�s�>��g!^�ȇl���,р�8j�Oa'~ŢR!�iY_pO�J��9���|��"�]g��'����b������b5�Ā(h�L�A3"�_�6�K֪M�a���=��q�V�}.��& H���h��fС�'%��C����;$܎sP;/�����^D%�N�wL ,�<Qşz�j>Blo"ٕ��*Tc5q3��M�az, ����Y�F%)�q���!��hRp� j#�{�5S�2��#���E�o$�;=\k\�5W9b��Ӆ|F>�Pe�R�TI���1K��Gݮ���u�Y̼��Y�]�̡�AG`+E�3�7�tw�	&�j].�.�c��l)�ml,_}�#�u��{�ն,������Nb����#{�qM`V��f�o<���vK�GR:	�[:S�)x��y��fCVo��l�A
�@mSG]Τ���_]����-,uo�Q�x�jx��;z�%�*jw%�d��RW{T��]iX���2�71O�A�b�x[�	���\�l�@k,��^�ր�8[zO��Pmٰ�,Z-m�7'�����3�\��9��Λ@�Y�����L���?�r~�ΰ�� ��c������� ��m�����'�OPQ�Ox�'῱��@��w�u�[!AV>q펌�-����@�*���N��O��z,'�Y,�g<0VƤ� �A�� �$1��ay�,��좁�r��	,���(<tK���A�L����~��9���	,��v�����	D;��q�9���3���s|;��k�z��|�}�QFه���v�n����T����M�;���W�w���!R�Y���ڨ���-�ϢN��b�!N�����Zy�l^�ǟg`x���e7 ԰}7=�8�W�w5�
S�ӯ�7�0�y��z��m)�8��a�ї��̻��_��A�i��[W\D�'�u�Z#��ҭ�ڲ�݁���u�w��M�+rXٚê��4rX�>���No��t/2|<�>�٭2�T�ASŅ�WO"ܭt�ڤ\�8����T��R��J���6<�g�?C_|ƚ?G����V�6��Uj�+��W���̫_��o��7q+��;�m�~�����)����>�3O�u<�����,~�3��e�;�0��&O�L�<ҭs�yZq���:��U���P��=
���G��� �Iƣ>6W�^+��O�.KV[�ފ���yR�pW�}��
F�8���T>q����'�+S|�u��v?��eH�C�M��-HΠ��/�(F>�"Y�	�jmqi�&�-�Pjv��
��֝*�%SP��UIJq'47?�d�'kt�����P���^�5Q��P���1[�x��욳�A�H>����XY)�sn+��a
)>�J�ߑ�ѕ�vG���	�V,�J0�D� �y$ht%hd��T�']	\�c_<��s��p�
�ľ@b���` j��i���DyI��&�Q�.�1u�X�J��P���])nv��v2���(h�G��2}�h��IR�k~}>9��A�X�A�-f��P{��:`7����������;0	�gJ�~ڭ����O�˘�n��;/�.�u��j��}՟��lW�E܇Yb'����K�� N�ұ,g/�W��s�\��a��2j:�j隚�%x�*3��=o{b��8��8�QS�US�S���um�̱i`��g��@��W���4Ƨx�'�!�I1�wO���}���k�b).���K��c����D[��#�}��������$���������5���s�^�d	�@]~��t��O� k�G�>5��V��OI�4ߠ��K��!�䔤��� +$}f:���?���tH?5%�\�B���tH?=%�sE
񱮗4^����9��r��`q���PK
    �\IB���  �  &  org/sqlite/jdbc4/JDBC4Connection.class  �      �      �W�WG�M���T�""h+�����V��@K��Z7��&�nD�Z��_zN��9��9��<�T�;�K��Ŵ���s��o����� ��c��C�h��CG>��%A�:�ch�Bq�>Kܬ��~E����Q�Q��y²-o��l2�j<4�E�.�<ǲ��Q*�UL_uJe�xw�G�Li�3��Z6���幓3�E�tdK�Q\4K���X.Ál�)��E���ե�y"}ez*s"S�mnzV�g�V����3��e�*�9cM ����pb��, ]C���Y�ӆg0$G|A�%-Hy���$ݶ���Y�ؿ�t��q�z|��C_rffF�^	�8،ܙr]a�Yvx�pT���$��^�e�j��ba��b��KDH�ܢ�V�uǠ�TQ3Eå�)���*Śp��e�$�vձ���d�qy#�=[�'r��I�h]�
��Ub:6�;S�q��._v�V���^'�)��J���'�ɮ:��P�[Mt!�3G�ʓ�j�i��0U�0�3�}�9�C�0Ay\�ޘ�2t�<>��t�]4��KK��t�Z�
�A��Y]a5%;�
���\�e�Qg��á��Ȳem�9M�b�FGE��+WϤ�P�t8D�HX���E}���A��8���e��!���H	�c�����B/ʈ�͝!���B����%��k��9*�FO���#<&gÇ�ֱ�Я0R��	-P���o;u�
_3�+S�ơp��I!4>I�<M`�Rl\
���RJ�;|��Xgj4��Y�$˘�ҹ�X
�[��H�6�/���܊SZ�'Π
�Y�
X������en�Y(J}�����7f��d��C��P2����~�K%�����,�?���[2�#Ky��[����7�ͯ��q��QD�ú�J�)~��� �)�g�.�R9#�^:���ѷ%ux��K�_h�nZc���t�]����r��%v�h��A!������ ����]��R/I���[t�^C��z���h�QA}�9qE�Rk?����G��Kk>R`�A����(ơ@q!p�W*��;�-���=���N(M#�8��߽U�{�>"����H�ô��{G�.њ��'���֤����%[%�#�bZp��Ї�A���)�KI�N��՘���)St�m趷е��E�U��,/O+nS"܄H�<�A>F�ҨD�L'aI�=�7!�z�۪��g'���T�Ӓ�!�?�z�̾�?�虠�YL�"��Q�\R³�G��9�o��I���FW`d0���[�g��:L���}F��>;ڱ�vF09�
��������?I��dIj�P���GC�I�-�_�q�%�{T�w�랴iHVs���>�m�Nc�2f[�d"���8���t
+-�f1xpN�:�� �(
YU!�|�f�B-���5	�i {R����J=����Հ�(>ة�.Rќm��7R�8�ņy_o���`��S4�6բ�A�"���J��I��_PK
    �\I"1mE  �  ,  org/sqlite/jdbc4/JDBC4DatabaseMetaData.class  �      E      �T[S1>i�*VE���T*u�ȈU�KE�Ug|p&݆f�[7Y���>9�?���%[j�V[}ٜ���}�$�?�}'�y�=@I�O�B�St�Q����^a4�)�A5�>�R�l�EK��<�h�{��׌��~E0,HO����J���s��;�}�i�g�~/�6حJ�Y�>yp?���k^�J<�;�
|���U$��v��.e
[�#Ϻܫf�.W*7��y^�B
�M�@�p,��h���������˥RnwQ7ZT�n1:T�U��0@��ri)�`%�3ƗQZ�7h�.�5?`4ҡ��p� f���84��`�*�K�q� 7��5���4ƃ�f�b�-�����qhK��EH���{Zф
]]f�)���Us/b5��(˲�����
�u?Ъ��@T�B��z����[��4�a�̘��x���_�I�ƥ���]_	��M�`��])<����7��R 2����4J��
=͠��l@��h6oNiC����ܰfx��'o�J����m2���曨
O\��S���n�]�R��{���R���k��*�YC��ԏ3���'.�ąx�x��x�D3�ף���yJ���3���0V(�7��
"	��3W��+A��ޣ��C�F�,�Y+MG���3l��;��`��MZ�C4҂�hb$h��?;m��8��}XO��x�`����<�O�x���g��)ا�,�s����O�����Êx~c1��50�a��1e1&�h��I�V�{��[+�ET��fgЊ;�Eۥ0f�`\�+]g��#�Ɠ�͌cܱ3Q�/32��d�U��J��wb�k�h���X���ڸ�=Lu��DnX��/PK
    �\I��%�?  }  ,  org/sqlite/jdbc4/JDBC4PooledConnection.class  }      ?      �QMK�@}ۏ��jkՊ�EA�H=U<X� A�J�d�[�]L�ſ�I���G��iQ�J��׾�ff�����16<��b�ź�:�s*�4g��A���ֱ`�R��� �=����Si�i�`䐡��i�ߏè�__���wZ'"nk�Dd�V-�M�Íe.�d94B��a����?Y%6�eg,%_�����T�X�����Q�+i7ښ9���RF���ve�Z��p��o�>UI�{ڟ��rt�S���Ԍ�K�O��/��=S�C���,�-O �H�Q�4%�dx�&z�>y�m��J֯:_by��J��}PK
    �\I���6<  �  -  org/sqlite/jdbc4/JDBC4PreparedStatement.class  �      <      ��[OA�ϴ��M.-QQ.mA�E��%�(%���t;�%�ݲ�&&&~_|2����2��maݖN�Ξ9�w���?��eX� <S�I�xA ������r,c�E�rl�Ss�3�JY��4G��d戞PՠfQ�9�n��}��U`�3�ɲ�R��{4o`$��4j�S[�ߵ`�9�+��FG����nmn�V�٬LmV�9�a%f:I,�P�ɖ�q�7mI������<�� ���]�4] 0K�X���XT��%�0;m�����l�#-��"0R��m�8�F����!�5�c�%��2�Rw-0;�ū�Q�-��E��l�+ɦ+�[��%=�� �ܚ�-�nhC��=J�f��]9=�EE7M$Ѕ0ܠ��¸ 7(du���������� d��h�^o���&�?�#���c���=�M��AͰ*l�LY����)���3Q��j:w����������TO4?���[/�A!0��o�\�+M2��}k=Y?��̡�ԡ�-^��0���-��p��݉_i�	�[I�/����¿���`j� w�4�^ 1�}��~��A�0�'
C����J:,��<Xr��E���'0
7}�1�a�H�jo�� Lj��lK.������{L�=��D���tO�u/Iuϴ�=s���boa�tk�ZA�e�oH�_�>��Ƽ��ma�*o��V�%��{�r~ʜ?h�
���W�؏W�.�Q�')ֵ���E�5������r����ʽ=�bc�N��~���X�a�EF�W��!\���/��_<+��c|�0MOD��?PK
    �\I�,�A  f@  %  org/sqlite/jdbc4/JDBC4ResultSet.class  f@      A      ��{|U��l�ۄ��-JëlSdy
��������Iڤi&��d���2;�6"��
��X+BDZ�""By�E���/??�{gv3sgf�I�ۙ;�~��sg�<��Ǟ����Q����P��j�/Q�����k�o5�����Q�T�z�n��J��ugͱx���ni�d������o�����u�*۳)M��ݺ��-dF4s@IcKSw6��7�����Jk\�+p��%5�\��hk_֧�i�_�Z�k��X
,�h@�c���8&ֽEݪ�Ӫ1oO��|�WK��-�T�j����|��\Q�|�󊁁֕8"z������������c�jLq⊁3��W�Dڠ%��@��D_r�ٙ5���06�-L�!~4���c�՗ݖH)0'�p��1��F:+�M2F�Hi�P
��[�n����VG�4˹ov)�R�-���XB��i���F?�� A�B�ΦSꈎeB���t�VϷ��y-�08q���9'����6�\T�q��.ǆJ�8��E	#�㼍w�2�Ǎ�C���]ǈ7�E�$��nu��_�=���պzح!����ۮi�ܾ;���홴�.J�уY\6.P�����y%�މD�8�t\5դ��ج�wl�l�OSS�Y>��n�sA��B3ٻ�y��gT�5c����U.4���7`[|R׋���'�\���#�>�Un��tC5'J~؍>�����3u�|2��'�	�i�Y6<|�x�-q�=k�
�gJq/��eΟJ�N
9|�����S�j��8
���a[��邘wݗN�V{CZc�ꄸ!�F���M�ص{�L�C݋�;=��]�޾�m��:���Q�|=���O>c����9|D��	��C���U>N/i��� �#��VKO�� �$VH��*pJ�4)ϫf��6������F[y}Y�������ГXesϠ����PC���T:٩N7��J"^��6�ݪd���U%0�nJLv��Հ�6gj[�l�C���UK��J[�F�����#y��,|Pa��u�(��0kD�"�S7�]ը�ocR5�Z-��;+'SZZ�S��p֕���׊��p/��U��а� �˳�vr>��xHxW�Ba�燭�p�A%��a�'�}+h
�Ԉm�lZS�W,1�M�zяvdl��6>�-xD��Zd#0�ձ�&���&T�� �q@���O)�̚B��V����ޡ2�=l�$�y��]�����1�܋���v�"ۙΪ�ɇt���!	��#�9��;ˊO����]�-��������x[�0�o'�&��5��٤	���I^a\��g�2��7y^�p��h��tr��Օ^K��Ϛvb�y&�����
a��������&k�&o���Ɂ�켥fr�J�����ܠ��K"jj���硉�gf��,�x��� �P��/8�[`�g�����L.Ϳ�h�摉f�[Z3#6�L<�LF�_c��"���4��恍�y~go������{�voT`��K���ɼ�ɮM�IQj\�o��,w
�O=ߛ�8j�"�Y p%(,�{ޭ���[ݲt/(�Uf�o��U�1hī�v/8� ����#>�ଳ���(�o�Tc��IF�Ĉ�!p(>_����kY�W��u%�[��Y����pX$ک�_��x
v����G�Qx����'ⲳ4���p���h���Bh�BL�-����{�ٰS9��~X�)�4v���^�'d����1{<��q|�3����bVl��q��0�FC���5����7�]�w�W�Y���<�ɜ���t?"`O�aϕ�ҏ]�ɰ�jO�3|�Vv�T��>)�����
�K����kh���t��U�FJ3���pK�Q�f�����2���,��g�N,�}9�gABJ���.8GJ����������z`�CK ۚ�q3�����]���Rp;Y�X��>��;BL滿���l$v<�j`Pn`׌�s�{F9��2KsP>DR�����|��,�'�i6��`X��R��,�E�H=(����Q��=xkF,�{��<��d�����W8�z�S2�G�3�߇��G��A�;(��w�!ile��d����?Rl�4�Cҙ�̙�L��LY ��&��ayI�����3�h�Z6�c�2��.���OC�r��S��V���Fo	�������kUv��C����#	=��o)nQ�Z\b��	��(ލ�8�_��q���C�ƦʽP%T��j�K|Ա��;�'���]�W���}��\exUIv\�+�uHS��`�W��� �	�
�Q�=d��� ۝�׹R�WȮ�x��>E`+%��`����0An"+��� �#+T�������\�۾>KA'����w���0h�5�.� ��q���淐39mͧ�
��+)@���
��̑~>� �gC�"5p6�YWO�U����k��um�;��5!a}a
��%�/�uk%�Gʲ.qe4Z�h��M��@�B���z��q���/O�u��u��q������8���#pq]��T`n�a��`n�[)[�u�Sc)|U��o��(����= �;���C�����z��}݁m����Q��j$F0r'|���	�Kҝ�
�VB�E� -����f')�����j��a�&%Hw�7���ߢ��"�_D�ߦ�wT��CA�MP-���R��T��C�OA�"�ѻ�{�����R��T��!x��xvVho����S�< ]��1�~@	�C��?ⷩ=�Ä����C
���G}��(��"�q����G	��𡟤�'����ǔ�<AP���
zA��~~JA?EP-~Ny����&��?�g)i|��z��s
�Y�j�<Oy�}����� ��ߐ_�)){1�y�~�����2e�~�p��x����/�/(�_!$ϯ����u`��W�5���	�����W�u
�@hjc��_�^ߐ��_S�I�|o
�o(�΋�7K�W�6A���xo��į,��j�[x��~���w>���{�"����>A�|�w)��E�i��C��x�����PK
    �\IP�*T  �  %  org/sqlite/jdbc4/JDBC4Statement.class  �      T      �T]oA��P��VJK�Z+*ʗn��E��1��@jҷe�ew�]��O>蓉� ����D��Ν3�s.3�������1=HR��q*ũ�
�X]��k0�UlYι�~0����IK�2M�{�2k�SFѦ��6Z�䯇�.w:Z� �ٲt�8�!�c0�.�|P������Ϛ�mO����^TF���� Y��'G�����QS�<W��溵R 9��у�5�N�%�3��g�bOr���N��@G��g��2��*���875o��Q��4���9�*��(-ܷ��Α�0�Z2���DY��	K�	�6��=F��R.��X�1��♼˄=E8I��(]��Mk`\�K�+;֞?K�����#!����P�L���x	aƁ�806��AQ��<iMo���cd<�V��7�]'
�X���wT
DIM���uT�x�ȯ�t	�.����K�$Ka����:҇(�P�
]�	&A��yɢ�Bź��J�}"_|r��s}��.���J�T��&>J�g���h�|fZ�n��X�Ϡ�O;����iT����͉ݾ@�@w��X��,	T
H�%�Ĩ��q����PK
    �\If1�cH�  �
 ,  org/sqlite/native/Windows/x86/sqlitejdbc.dll   �
     H�     �}|չ8>��$��0,��
Ѯ4j�F�Jl	5�@"�����TfCPL�ή�t\)�Z��Z�[ｽ���.v���B �w3Bhȋ���y��f��~����Μ����<o�9g�wO��&���グQ����������i��f֮K6��.�z�9�W<����8��=�ȣJ��Y�y$�GrJ�����?p�ر�NF�lA(��y��L���}k�h�,ܛ%/f��c�+��<K,�g�h���C/?y/��5y=�c�%�Ǜ-��Д-���e��C�ق�<���e��W�Fy�N��/e��X��e�K���>�>x~i��ǎx�Aֈr��5+x���8&����s�_�+�y#f-�>o߼��p�,�[6�|��_|�C��pIc�:�\蚒�U���^ɦ��?O9e�/��a��9O�,{���#��}�r��;���_�_����Urz�1��K�a�3z�Wf���Z�ꞥ�=6�S̭���C�6{u$ė ��U9���jm���g�+��@������g)�D}/mEJ|����Z�4SZ�Sy�zh,�86KP?��C�ݯ� 	j�I����aG�@G�K�6[���A��s��Wq5j�c��BI��;e�8q��)�EN)���d��\]F���C�Bo���k���7�'���«o/�R����CB�eUN3��0�3���tD����R�_E4#�_��XD���3FR �X�z\r�Z%k ����ݧjO0�3�uI�К��	��Mɧ�'W���t�߈67�SlR<ǞZ_�Y
x0�U���_r���X,b�}=&|u�בx~�ZN��"�9�i
�y96�~��� <;����^�̙�v�5N'�t�ObKe �J���]�{Ƽ�i�Vh�`�Ϗ��a���4�*�r�� jk:>�5��T���"F��Ȓ���g�q�w�|ri����>�z`Nf�vyjYy�A#�U���Fճ��F���l�Ԩ�Ο��+�Cl�)���_}��|cFe��Nv�3�:;{nG�wA^@�\������g�B�Ҕ~���Wl��+��ҳ�5��'XjʅZ�3W+u�D/�R�6PT�UNK�3`Pˢ�k��}
��`�`r��b�`�&u��Y������ �>>��T?7�f��U�v��-�x�#M�������,�jP�&�]�]�a�N��]�����:I���<���A!T�C?,N�������x���j}����a|�_R�/n��Z��F����k�d��f莅��A�b�� ����M;�)�+�C��m"�����緒E��s_-XN��m��!��TǢn�M���M�5��%��:���DS�����W��+���������|�:-��Ƙ H:W�#{Qh@5p���(�2yP!���(�zR�g!z��?�O�������2��" ��'�8O��M����&�#�:�Z\nP�}��$���&��Ǜo�X�¶ki�@8���k�E�d�(�V9�B+�+R]4�Sp'>�Ifj%u��p�U)�^���QcỌ�w�.�X�Ʈ�eݹ�(���+{��sӯ0���,��0�œ�Ǔ�Ť�<���w���_@DV���Z�)"� �~U&��.�����B��Y�Y�)
V�|+r.��.(��e9�9Xe��&F�M���m�vL�!��i�#�BR�9a~���"��Ձ������Xԑ�"�~W�>=�2��&��?�*0
���Y�b���0t���D�׽ɑl���I�	��{�,L��kJ#�����D�X'��d#9qB�F_������?S�6�<�M��������{��8�X�e�"g��(:�J/���	��ӱa_ ����������bf&eBF�+I���e&g;��[ʵ �e"�c2=�?�Xb��w�И�)�M̺�y��fR)`�sL���R�AC~���C�pU����Yq�V�&+�����
�q�[�~c�?C�R�H��ΐ�d�j�o ɹWԻ�P�|�\OXn�Q��b(���X��)}�m�ٵ �ح�[�R)G�����Y�#��X��G��2�-�� �c�M��y�C�P�A�X����
����ġ�X񰔵�����MYN��Q��m�	(F)�&a!W.�^d\���C��A3���-��ۜ��Fh���	∾߈}��A���ש�X'��%�9����Rf+��B�8!6)/�@^�j7;���n�K�	L�R�>�O�rKrX0=���ZpX��$1\��:qp@��݃0<��`��doB u%ߌN'G'-I������A�>��N�f�f%F���BNBJ ~�?�Y�?���z�3�Gf���?�3���O�&J[g^r��X7R)�+Q;����g �i�7D��D�M��P�-�W6��eN�]*��=��q�%���h<@��v>6��{.�L`�%I��y����1�~cB0�������k��!JlN��%�;\��Qu�T7�5u�#�>7�.R�r���9G�{cT�|�w1�ی�5��3�:���B�W��,�χP�w��G��+��`@�@.r�F�~	:D��K~���������r'�1���4X+����z)C}���h.@ �#P�A3���/8�@pek�ϧd5[���bqjYchK�4�W�,OJ�<�8	�*���\� �\��(��I։��=��Uƴ��S�}zӛ.�~���mJ���%W���
 ��O��^-����D����I6�j�>��t}����MB�J�{�H�JÆ���Ӱ��xk?�[���O�1���7p<U ��i����N埋`��aDK��0��YU0���v��v������cU;3�O�gP���� -�3�
GRK�N���9Pv�:4�v	�]Q�-��S��*��}����g���I�GЂ~�+��)��C���5E�3T�y:�kD-����Fj��B�{�� }�N�� �+�i��FA�w%���oM"��Dw�E�i����r��y�1��xE{���	N!szM 	ڷ"��q-���?zՠ*����o�۬�!$�m�6K����J�F����O�V#?:*�HH޽>������&�O�f|c�%�����}�7�����C3�6?yP�\V-_v6\v�_� NXj��`���pp����7�������_�f�ܠM�~�TvuԨ��"�f��T��$xNOo�=HZ�	t7y�WH��O����ی�7�S�5�VG��z1MH c/ I����H�2�@*`Y���"Wyp��2}--M�V�ˢ������iȨ��$xn��ʷ(?NaI7FڰrЂ��'z˘,�P,�5�aXCu��
�u6!Ş�2�З?AyY�ob+ΕG硷WR��|������_>g��ڟyt9�:^�~��( l&�T��/Yo�ߑ��A�sp����\�,7�F�#UDH#@I�PbJ��}����aq�\���B�b�π�nkRf��(
��̪]hB?�"0E\�YlȣR�}1��O��)&��RQ�"�ԋអ���%���s{�#1�x����ʋ4��q�n+�c˷�$�ϑ �|i��R��������W$�!E[�!e�M�P O@���!{CV�1���|,#�F����N�E�$�	3�
���ֻ��w��ġ��9������0���{S��0>��H�1���x�������ص)1�����U�����h߃���71��F��o�)>���a�1�q.�j$�%$�ur}&,@��*rZE׾+|���'�Q��'�w�uIN@���ԉ;N.�Jn�3F�[�r#V_zք�
�=�t�$��|"��c��]��y���J���Q;NHǵ���/���Yҙ�#х��V���Vl��+�ՔZ�w.�蛅ʃ� TZ����h�/�Be�?+T�~�V~y"�y������U�Ѳ(�U���I,����o�9勢h-��+�oS���^x&�Mp�/��`yKm�rV���d鄾0���q��o�d9N�}�yZh�o�`����siY8A-��7�+����w��e)^Dt+�*���*6G�e����4�^a����fqUr�iہ��3Ӽ��NTR��F�v,�;��� �tâ�rs]!_�&���ri�[VG�Rr��˧b�yv?Pn9���|J�`n� ٠q+�������"1 ����&�m�m�K)�{����G:9_X{��\�������BR�݄��u)�nb3����|����H��!��� �T[�/�˒��d?���O`�k�C�0Fc7~mƯ��=W�>��U������qB\Gi���tq�p´�hI�����0��F®�̓�_���K��;%͓��
����c�L�� �F�b3�G��E���3z[x�sp��tȱ��-א�)@��c�fC��s-u��$S����**�}?�Q����
`����X��^��C}zz\m�r�]b�\�J)�C�7��d��jp����L��TS�X�ME���5��Ǭ���iI�Fh��8d�o�����=s͈w�J7]��1h�Ԙ�2�e�w��aeߍ\�C����=�@�2$��YE��#��՚� |ϛ!��rg���r�}�Q �~}��;PޢĊ5��ei#���>�aqu�/od��`�Xl�vd�R,�,0��h��*�w�2�� ��w)�i�0]HKUN+�Xڤ*���yt,���M�7x�]���Y��V0ʇ� ���_@"F~�I���n�����s�G������mO8%qO�]F���	O����I�;2B��i2t.b�p�:��F��9��9�G�>*��9>� n��ˑ7E�g��Mb��џ~��z�����kFWL�$ʳQ���BCJQw~y�1��oRGW��ڟ�@=.*��03���4A�[b?���������c+aq�~���UH�\��I��Ŗ���������{�g�;�\�o����튅���Y�M���"Z��ʹ��-m��5,9��A_yUZ[�����<v@��q�Y�x20F@f٤�a���ܟT�0:�?F�P ��}Te�A��)M��}�qKj(S����q�"#�ߩ�H}I�k�J��6�?�M��o\r:6�?ri�V&iV6�˖Ygc+�ҫ����.�;��l�z�ъ�l�����?�ؿ���ͯ"�xw�9�K�W����<�x����_t�����#��������6߰X��n��Ȓp����>���%�D��Rً{��9@�Ȯ�S���ߛ?��O��Ã�X���)��=�vI���5	j(Y���P�h�(R��ե�@ߏ��[�5�&�nhMVÍ�Uס~1��Ԟ�Kc����\]���u�����y��-�����n�򐫃z��Q��Юǎ��cQbQ��an��Ѐ(��X��"�@�C��f�=� A�	�ڿW�R�о�!8�+�5
"��y�*/�*2��!Q;K�*n	�2�WA�Yz�{j��s	:V��Cߥ��q'���j�H�Oԡ�U��3qt�'��Y�eB<~��)�֩v���,��bri'�L����w,؂*l�b�o9�n�����;|m�mh��c�5$�O�,����V�l������-v����V��z}c;��d5�U�Q�;��G P?��]���R�T�A��
�Z{Q�rw�ϭ<��>�ٸhr\��1.�x�0��Kǉ���R�һ[���۩i*�Ty{+�䔰q1B������� P,��=����ы��)?����!9�]�����Oa������Ѓ���}��o?)g�� ³�|�P]���8%t����#[���;�Bq���C����]��x�e��r�%��௩ŗ�g�E� n��J.�������],Mrp|����gz;bګv��A��T�n��Q�?��F.j���GG�wP<h�}�ҐJOnD�yz�;ܐ��j��כ��8�4)'�;�`��R��(���3r�M�T�`d�{`��B3`I��A����>o1�aQ�2 ]�lG���Ũ����cu��Ȋ�m��F�W˾�A��\B>�K��SB���1C=.�)���2³X)w�@�"���UF�yd�����i���/n�)w�=.|�q�����2蔯�����8���*�>�-�]�}U� ٿC���9k�8���El�����\�;��~'4��G�w�����XtMOC��;���4dx 4?�J<��v��>�.��_"?}RB�|S�#���{Xo���hx0cz�C0�^���鍋��ch����Q��F��9؉����	���tA����"g�A0c>� b_B��xr%�7�
��U�O�l�ވ#>}?��Ҧ��1nW<�N��l��`� f��1Z@�m<��U�+GVo�ǉǡY tlW�K�k^�������*����Ş�*y ��ؿg�!��X���	 ���S��9�����F������=�;� �� G$�W �E�9���Cy���D��ՍUN��{�D*"��S�"a���]�D{a�r��*�ETD��ضm��%��hw����M���t9�����H];(ǫo�~�݆��c��L�,�S
L��N���	�]x�h:�,�1�;&������/"�R~z�Ů�?����٘�#������>!-���
4�8]���f� Bv�\�}hV\A�$i�\~���]y��N b<�4�"ٷ�Ĺ�I��è�N4�.Mq��q�#�rP��?o����ˡK��BC�dS���c5zb��)	>#�<��OSE}���*�a(��1��O4.��L�DG��V+Ju�M�!#`�2�j3���p��Xa<A���  '������xp�<��(��9*�G⻪�3Y��������N�P��뒿���/Ug�(�?0������� x�-���G ��|��인~�q���b�ѮI�~���wL�7�`}���(�(�9z�9�����z|���ö��#ء&������.~k�B�ӿ�ua�#*�j���#����Q[�:�⌽rs�c�A�G'�,�zb����bO�&⧱@�α>,�|D��}�$Hn%��cˡ�g8U��fX�렛Mw���!�}s'y�@�˾���r���8}"�wI�gz� �WN&d��T�M��Pz��n9��E���O��ף����]앃{�/�P!r�`�W|
�]��I
�	�XMR;��`��N�C8} ������)����,���w��}�`/���m���̟��e��w����B:\����78�-/z��%u�(�����b�|��?�\y�c���3$�����&�`JH�6��
H[@j��t�C���N���!��3<�Em�P��21`X�	\�$�~�-S�n��bj6�}XqJc>�>s8œ��~��R�6���W�(9��J��lWѻ\�6&d�����$2�2{�,�(g#��&����LW�y���:(����Dz��J̜�{�@�%��$�;�?�j0�+e��0�+t�O��9K�*~���{qx�w�q����Io1�=)�V���2A0���c� c�1C?�D��ڄu�~�R"a���Z��`�XO��5�4V��?�cޘ�VZ����;���LP�!93���S�Y��.�����1O��l�3kOciAF`����{�3���EQn�P{��1jDT�� ��\}������9-�<���J�\(�E����C�j
�C�Y�Yv�,rkt�J���0��Nf�\n
�u`x��iX{�!4��LZ�) �����M�N��;�O�ke��L������);�6 �`�����G�e�=��<�������&0��t�w��M5L��@CY:6q�ڣX}c�hf�GX��X~/��������:�82�:�3��9t��d�8.od륊�ح�pL�n��n�7U)6s��g�r�����Z�O����xϦ�;�m��B���A	=�(���aͷ��g���M9�>Q�\�����+�ǘ��I�B�� O�挬��}`ջF{z�jw�Il�I��=��ENc/�;e�����)km Y�^���p���aǠP��N�?s�M�*�Ն�.�ܜ����͢
��9l�t(U���jw&�դ=#츦g)�Q���o�C������~�?�Kj87�#a�ThU �7 (��	J�����NBҪc�����=�Z*aQ~nъ-��d�}O�vz����`���]!P/z��`�hm'16����]t��:<ݮ��7�>�5��~�N���}l�'Kw�>�}W��b(�Z��ӿ���稺�B>	��Y\�j�O'y�͠��J���~�5P�DKiWH�Ԋ͸4сB�v#�O�G�Ϫv[�SB�	��x:^i0�=��k�=F�7+��#r�~>9���Ta�Q�E�/���f�#�x�\#��I�TbK)���;�韬�tj%�Vn�FUaܔ�ˈ�Z�QS�y�4�ީ���*�M�b�b�`�@��3��v�v�As$r��1S�XX�o�'�Bg��L��F�D���Pp�ej�����3��?�����I��D��L�w@�~���p�L��=����*A(���W;N��ilOx(c�N�s�� =��Cgt:?y��ե~����!=��E�H3�y�Ԓ�]!q��	E|�;fԂ
҅M/�]���j@@��$~����/4�
����-mf!6���U�@]���W@9=hW���SM��N��ZPX��Z1A��:�������Cܯ�m�wybkݯ���������}>���'�G�*(���=�;�ѽw+��d���-�m��"�<�Y��������8D��`��?��G���-�z(���=�`Sc&�?g�mI�t���D�G�5<�χَTꂾfQ+sT*W�g����m9z�粕N|�Sa����ZL��zؤL���;XE�R�f9���L��i��F���f�i6Ӭ���>&雴� �3F�A߭F�}%P��۬���))�Zf^,�o�����0Qa�b������AӨ�w԰�=3�
���"BâǦU8�WoB�5态{w��ؓ[���gqjL0���3��LJ6�v�P�+qh�-"� ��*hq*;��F}�bD+&�����F�$��3PO�Pbg+mjw�ڟ�L8w��������8�[R�;����m���i���m+/�əiaa�!�(L{i3�j�_a�pp�Eok�X�
����0�� �H[hg���/̔�U:Z���Z��*A��b��>��m�6�U��N�_ta�{mzb������]����O6y9ס=�w��V��5i`�)ف
�Vlu�=}�L+3���O��X��3l���ddצ��9���������F{0�������v���j7�w��f�W�X���!k�C.�����gV��;k���>������_1��Z���Fć3�dŹ~Z�A"���Z�B�Vb�K�fv"��szɉfSG�]������4�ԙ1� /E�>�x�F��TH���X�6�2Xotn)�[')����Y"X"���߃RBLR?�"���~�thh�����SqX����YײN�G���X8>����עw��ޱ �=���}�H���B(��k@lT�>1VP&y����5V�O��0�8p_y^��o�} y�/ޖb��7"� ��֨u�B]�V\���3ԗP!{�e��y�9�&��h�X3Aͻ`J�t2φ!A��C	����l�L��4�|����u��<����U���h��uX?bt
�P�: ��I��%� �[�)<�Q��Ǎ3�JW�u5������1����8K�5.�V2ԝ9��z��-��)&��s_��8�b�fd1P7Mof�hC�ץ�V����&%�6�]���]b;;
XKq���|sh�BY��# ���w���B���\]����ݨ}_Ew�r�?6��b�6KR��b�q�^�9)D�l��ϒg����a��~z�g�a��@����p�@�Jj��m�R�ڱ`��眢�h�{ ��_�;��&�o��%1�I����%�r��	�V>?���
�3L�,�X���(l���{�L�B�7ҫ��E��{ ��"�����
Y�4�Z�Vf�?���f���_:������D��ܻ�o��%J�{�q��x`�,牚�<�+論Ae3-��7P�0���i[��E��m�*ӏk�Y5�zhbr�6�z	��끾� o<�M�{�>~������x�}�x�.?='>|_'�a~���i[��E�{`��B�'�Ev�\�7wrN��QA��h��@��������4�T�K���[x�Yѽ&(�t{�z��b���*��QCYp�X�.��`�5�%V�;9%q@�PI5��VI�O�l��5N;�]��4����V���]r�\9YmYDf���v@jV�����I��UT����z6_%�wj���5,���N�g�;W]8}@�+B���0Q��w�<m���1�W=&��R<��#��;}�:P:^J^B_��Z%Rනz&�G۳�!��Qwrzg����|U�OWh�P)��5���I�:5����]��~L��NU�L�t�Vz����:,�ٮ������.`�h�I�u��?�����ԸX[�#� &�ܳ��y��)�qǫ��{w�	�1��+sE���� �!6����$���a�ǵ����~$���� 0��I���̳���?�*Lj(�V��ޭt�W@tIl-Zj��a�M�/��4`������D�S��[�zˊMZ�u�E+ԐU���,�`�ݢ��>d��!o��vɎ�Y��c��+F蓸��NI6{�hߴ:�V,i��1$L����ej�@$jy�����J��2���2�d.�0Ҥ�zT|�(��2�hd��16Q�<PԨ��>�b�~QS��u��=ѽ���bl��c�v��(�_r}/'�/�;���_c�f�-*��O^��H2����h�=G�.A5Ǧ�Ç��yVm��}X@Z�����M~��q҂"�p�5h�~={�)x�G��`b��B)|Ԝ�%�f&
����*��w��"�����`��Ri⃒�tě? ��[��o�8v��q��$۫Lr��/*�����5�3͒��E�[��=�|k/�60���(oX?�'��,�EŽ �7`<�̨nǝϯ_[���x$�N��j�4 7�[gJ��akX�	E���"����`��0~�Y�X�
(G��������z#�-Oe�"���NB�p�5�8E;��W��a�:�S@x!�=����rn�W���ڳ��C �j����8k������\���R-���^�r��f-4�χN��oyC1��ir�+��,=7��i�I�'#i���*���B|`�6�+��A�EZ�D�C��:n����V�g�,su�����և?���W��NE��c�[m��yr��L���Vi��7À��μ���������Rgq�Ȫͱ�:H[�'��S>���<�j@�W���Gj��|�6��e�L<m��L��W��{����$�H�o�è�����N�����w�k�����֧����GJ�����S~��חh�__��o�����JOE0Z�� S������ֻ�B����b���+NN��[5�����YC��[L��d��[�A/����x�kcO�U^����蠓�xJ�;9]Y�t�4��Eu��pH�1� ��y��H��騒�������S���)�t������l��Z�E�hp?���a(�6X�F�K�0FI�ҡ�
L�ˬ�:U�&ƛ��W�.�"��/�5/�X�'|������蕲V����S8>͍�yk��jij�����ٚ5����wh�+?<'��-�<޽��-iV~�\�"WKT������!��b�"�Hl��5�W�j��p>�'c�+����OS�)��s������v7���L-/h�5S�L?`c	�1פ�^����Z��xT��a ���>��
��4��P7�q�+	�G$ܴXwN�u%�}����LV����;b=������Ɖ��ۅ��Dr~QM�d��,�F�a�����u�צ��t�4����s�grm�&ΩY��ދnZr��<˼E7	����P-���_HYJ�:`66���) ~*(z�^���\�]s3>9�>���3D�z���^��au��Px]x�6��o��o�j���bU��)-H��Ȇ"N���UlѻR���V�����mӮ����j�3�]ob��xЈ�mn��|k�<��e���K�(r�b��(����z/�^<�=���ⶭV�O?��|x�h#d0]���E��?����$v � x�ٯ�K�DP��m�����`xV@֭�K6PiU�a���k7�^�>�XW�+���ldc�`>�f���s��^&�9B�v�0nlX ����v���Fg�-*�Rk�@�k��5�r�Ч�!.�m�y6�I����K�U��.|+��V��BA�.zi�I�`�r{�L�@Z]u�;���������7LՑ�IT�L���a��U�+�0+{`��=���yv:�������G-�ЏY3,�@�����@�M<��d��ʽEO�S�[1P�%R��r	�S�o��S��=��s�֬+���c0�r�C`���M��'omH�h�J)쭳	 ���Ur���K���;8��+9���&��ϔ@����Sޡ���x��ʬ��CO�0�L�Ћʜ���c��ݧ��<G՞L�_ ���w_<[0�Ζ�:��Q2ר�s���)�֊n�C��x��"�P�t��}���˽�g�98wbQ檱r0��T�G{�܉-�2��YD�Hu<`�s����j���EX����4 �����\?��p�>�:��!V���]l,�L�'\=�qg*l�o��ۖ;��s�9)�{�����`��XYX��V�'�F�2G�g��%#U_ڐU<�*�������4�[���`�_���[��a$���N-�Jz���]}�zR�[��؋�o��䅚	ϜW�D�O�v344^�ea=j�]�M���j��^ik؈�KK���hd{Ȟ@1��z�^�^K�[J�*еoV&h?�&Ey��O�(,h�����^3��X���ӕ�`�X�� dk`H��~�K�kB��a�$~����U7F���T����&��&q�{�s0�mruD���FF�d�xޗ����t	�r��Q ��j��.�ܤFD�)e*Z�Z�A:����h�����E����#�׈?Z�h�h��7k����V������3��r�m�s����$���R��Пl�"��G�B'X��2�Gh�=_�8�4G�S���nl'�q�ռ�ޢ� �Ѫ �>�h����/�v��%�`vU�c�@w��#���P�k,wN�Hr�a���L��z���4����ԠV���.ٷC�d�A�=(�T�p�=��hTa��2O�dz�8�	��39��q���d`,��H9\_S�V���r��)�!y�ΐ����x��2�r0��0U��B�S�?nC�ʌ��i\��2���I��|��^~�ڿ8��#�P�b�f�@3w�Ⱦ?s�yўw�"X����}��j�ǼO����=0_�z���n���U�G+�V��WW���g*��*�:�V��Q�y1[b��ޡ1@/�yb>�m�n��2�y.��5�� v*�0y��\m��Š�F]�G/²�T�8�[hH��ҳ�+E�I�2�����͢�)B���빃��#��*�^ݑ K��h:�����z+�>�OƉ��M�ni�ɾCg�Ɨ��A֞���UO-��Hհ�O�ɹ�b�?�9���r��U膯��e_�W$��Q�a��
����(�vj7���ik݃�Z��Iԯ��Ƽwh_��Ua\����=������tY��Yc�5�*}o��0�Q1:���Tx�r����-�[k�eᵇBX4��l5�S�_�?=
H�y���|�Gy�����@Ԣ���o`м���'8�z�F�v�.�K\�����z�C=�)e����\!���6܆�w���Y�ZH�Zyi��E���ٲv�0����ѧ_E��+������N#�<���8yf�}��4?YD^������[Kr`��(�߀������De�������i `�eg���蘳~�࿮c�y�F��z�i��Pz������q6Pw��o�{�`�{j����3Q�1q��^�Gr�#)��1Q�{���`8Y@]�(4��}�4^i#����y�;F��ޮ�Mjt.|�~��� �rd��� �0^PC�f��u����l@u6����7���ϵ�\�	4���\6��η�D"Ѫ��I��y����)��A!09��@���A/b=�n2���2o�7�:ǩ�I�w�/kX��s��̽���Vߎ�a�b	�Q�
�V[�Wd����G����c�G��"�M���R��x�1o�����:����L�L`^�Q��r[�*���7��&�T<^�d̔;�7��e�S^3O��u0�1x$��u�qr”�aV��-!pj@
O��y�,>��X{��~2_�>���j�̽:_��#���`EW�y�w��"ٷ���
@��	M��8�����/J�v�u�<0y~�Y�99�e`DI�@�v+�?��Z;{�Q�5�%�s�X�&�ݛ�rg1�K�Pk�>r��)C�.�At�3�7�Y
ɩ���&}<����h���m~��O�6h�rp�d���=�*J��!�k��X�6P|���v����j��0=p��c��l��l���+e�����I�Ec�BJ���=g�+�`���y9���*N��bK7n�?���=ֵ���B�߅G�?#�SiɔY�t<ެ�*�UqZ�Uʭ~����P���M��i?/���=�ef����?]q��ɰ���rh�+؃6tv}ƃ�57����2ME�%��Z��?�MP>Qo�?mSϚ�tm~��M��Pߊ�]F���'����	�����F<�l9��Zڳ4��P۷ᚤ�L��^,wZ�V���2�*o =�i�g㖐�:�AJү}Mq⎤���.����n�oqf�}����֨=�R*oXn������S���,��%��A0>v�!Ž�y�e�Q~D���ˀ�y�F]�t���|h|[~�B�з2�����]>���9�f�Y�p��V�j��]2�ܙ���7���f�:X(�����5��Ne�iYhfeR������<ې4��7�;��{ ء�@�8�6�`"0���+&����Vȼǚ �o�ލ����q�`A��<Gnl�f
7����0S�ٯ�u�_B��{o�8�ƚ&<���O*W�o�<'�t�reу���Ӓvak	���*�� �>A����[Ҧ�	ظQ����ߒY�H<�:%��ӓٸ�{��Xp�3�[
0�����f^V,����ǯ�/Y�p�X{T4��5W�60��寭@��"�6@�o��@�KN3~X��z�2��F�y�_��ge�#x�b�
[��1���z{|r�{�d�����Ḩ����ᐍN|k�z�Ҵ��4�	 hB�O��j[��$���ˣ�}�:�\_�.�~��)��΢�S"ŀə-k��a�����W��,U��VXp0P0m���tПͅ�șܳT��ʕ��٫@V����Y����`�jhN�D��(2Ǔ-o�	K O����ƃ�8�i�7P�� Cv������^��e:���jG��w�.��z���9�H�?4�!J�Mt����0���gs�)��@׃T��ϱ�cq5ZR䒟�JnEeJC�D��:Ԉ������sg*�t^I�ŝ����P�p��;�k�B�#�@]��O\E�ʅ��O�x5�N3<��"P�(�s^_�dW����m"�Y�$�8(�@+�/�9	��l v�Q�7w��/�	h��0�.p�I�����88_$C��L�s��ZO,��&3M�����+;F���ӿh=�o S��'P�����@5+��2����
�t�_��H���+B�'�)������&�?Ձ4��8�p28_��yy����ִ�L�aԾΨ�a��H�}ߨ^���Q��O��?���vS1�Z�zS*��Y!+�bT0���A�����c6��-Mч7:��>��թ�c���:/�7����p�9r!m�S�W�=2�#�|d�0^�-�,x��Di��GF��iN���O(��S�|��(� �����ϑ������=KA��p.ZFV��'�ف�tUf���PI+O1�F�l�k�ݟ�	.�P���ø�o�(i��NA5�\�}�%F�fLc�04q����V�s�9�K��A��0��C������#��%��Gx�w.F:�~ZR�	�`������ÿ�s�2���t�Ө�xwM�ř�U^�)�x�l9_��Hzj��
�+���s�_�zy����WZ��D1�6������Cc�7���������y��}�o������ѕ���6�g�]���>�o��j�g�]�����.���϶?�����	T'���mt�d�f:��<hQN�%~O¢�Y55���o�J�l���<�-w;�e�6J��%�g�����W��U7��O�ⅮE�_}#�:��x�7��	 �?�g�?%�}Þ�n�����YR��7'�	���H
S�6�{6����.W��T��f��^[hu���<!���d�1%GK�_=����_M^0�����xM���c)E��^��֍���>.�`u�x�ι�/Q�����œ�n1B�w�}z�M�B��֐� G�BG��[�E�P���ѷ��s)3Ѿy��yS�[n7]�.�������Cמ��6\Mou(~TJ�,��&Q%�����B��x/C]t+��	<"��A9��=�[f�9�D����GX�S+pʿ;��h_8G��iW��0L�׽�Yg�s<!�.u3�h��^���b�</P)o��[�D�H���^�T�[���Q��o>��HN�dבI<Y�*7V%L����nGV�������T�N��@הwi�;��D�ޢjy}s��r0���,!E6�ٍ��xZ��/��}m�d�[�|RXz���n,�&�æ�қ��!8��X�l�K����W�D�mѥ�+z��y4\�5�y@ 7�[X5U�7���o���ZL_)%B�qu��~5��˼��]vr�)�3i���ݹ�.�YTC�;m�D��������{�����O9u��Nc�Y�K��,���u޺tA9�����wՍӾgG�Ny}�2����mهʎw���䙨=i]�]�&�\:H��ڔ�z�̲o9zr���:��	]�6�9ة�vjENv�k��2A[`}�(l�Ĥ�����Wl�<�海�Pb�5YV#�(�Y�<�W��Zʒ��j�(���Kb����P�qk�S���cz\6� x̦��֙��%<�iן�
�t��8/�y�.��ˆ�bؽ��rK�5�b���ӵ&&��
���s�['�7Y����Ã��_�i�2/�:'�Z�`�S|�T�;dU&x�rd��nc/�K�Rx@(�/�L7㣤�UQ�M����C�j�ÃZW�.�S�d����N�����Lu�7ܓ��e�6N	<&z>�0�#X�q
���N:��f���u�!S��N�*(s~$����|C^e$��x@'^{�x�t��q_1]�`�}��&�m�wH�O�p���$B�I��y�vu�����*�x��l���=�V�x�`$k��g=G]]�c�ˑ�T��Hq��t�> $?�`����ޛ(pf^z�չ�`/�y������)�|�%:�8��ͲF琓���Q���k�F6:O�M��M��5�<���wGp#ޚ�]�s���'.`6V�����W�BJ���T��,���@�����2O*�7���H������s��$
y��`�Iq�^��;U���7�v�}�J�b�c�~�z&�����~�h.�z0)I�h�Ƽt�$��Ȼc��cP�kѬ�ُA���ُj�K�2�g�h��O���x{��S���o��y:�|E�-!v�bޑ=D��εILz������-Ċ ���7ପ�K�����_R�_�����휾��ʖ�����i���5�xt�x�lm�rI���EM_��X���.����0�?W|�=�9/\H�O.ZY?��x ��?T�;���o5Mx�+�_�c{���oLX=N�X�������P\�X�c���D۹�u�B�z���\�/p�*�B1�}�q����.N�r�w� ��Q�i�:#�sp�+�X+n��;C��]׽tc�����Oyv3Tnמ�j�Y��D:�z�/	{ŀ��V��[��{��P�ؾ�{	~�R����LԯQ�F�ר�]��t��pWb����LX�t$�*����+	D��%Z�z7���fI�wMD�ӸR˧�ep3?v�8%K��ܔ�
h˾��8�Y>�ӗ�(����^�ǚ�`?.��bc�̄
'�u�1|��$$Ƈ������u:ޢ�U�9��i(�(��A���̭ESj����EY�
�9�D	�G�c��-tnAMM��������w������)���C '�ђ���힓)/�p�Z�L��x�s���-\\[�\��~��v�(��ʣKп�ׁ]��s/;�먳�[:��BU=Kه����{��u�[�ey7S�kx8����������V3{RT��R���{~߀���N9X��bP������9���/�eR>e�Q�#�7C\ǪY4e�O.�/�.e�wh�'C��q�c
&����~��-9�Am���g:/����(wĕǨ��'x�I�d��w<���ظD�� ���QBl8`kw��@n�%��s���oZ)��J�?�B}7�:��J��O�FWȽ��jN����70�𥳐ӵ.v֊����0U�O�3��Z��X)�oی��Aw�6s�)$�I&h�>�W�Ǖ������u	����󙬕Sip"Lt�:�Qc&65lq��)�2��ug��St?�E�3Z�N�O�i�79�~�z6�c��>��'G��j�A�r)�U��{��0J��&��K�7�Y���~	n���#��D�-N�;P5�ib��7܈t�|�Z,���b�2?8;�B�ҍ߇g;�p�@�G���f���L?�lf��R��l"�	���Q��UAD�`N�`x�~���+�i�X��e�w��zl>�N�d|��Ex��rY Э_x�_���_�M���^�nP����tL�u?WS%�E�iV y|�[��^-�",�-�\�9�N�N�0y�!H�a��I��xۉްӭ�
4�w�r��~�ꏙ��M�~���7��a�[XP=,*�r�6��&���>ug�[X�uL�
���kl�k������=��'pk�}�����el�z8�&K�7���� �<l}�6��2N�1�-&h79����Ֆ�o��H���4~�������#v�L�O���x�g�ß��4��5�7��`�͑��quȿm���픐n$X��VJ�0��n3%dbz����=l;�9�t`J�,$�~����"c��fJ���\ y%��?n�>a â���0���2����?��Y���ݤ�$���C0V�PIo���ܻ�K��σ��a@؈�]����M��pE�A�n�g���7��[&�-�AX0�l�?��X�C�e�7Z�z��t�d5{>���p�5��m�د�e,����������⮽�;��\N7�{$�������zD���x+c�p�x ��$��z$6�#X��|�-�]ݳ�o�g�&�࿽ڸ߿=�~�OX����y�#�������7���m��ǮU��0�Ӥ
�r}�� 댒��]!�8��Ț�'����'��������� ���������m�i�+����_��B<B'�=�p�s��n�S2�N>o6�'ƚ)�����%�K��$?�2լ=����V���X7�}>*�{����uQ=nE=�2�#�b��g�j���I��ޗ)t��'5A�`��~N� ���R;IJT��ZE�>z3���6k���V98���`#F���8��v�����!i:�j��]L�|>���ݤf^�U��~������k�瘹(~��q������Q�9_��F�����b���8]�XA�E�t�_�]�(M�d���jwuD���S��#�jġ�������L�;��L��Y-F8�1��>}���2�V���(��gA?����oY��O�f~���R���~=�+w_aY�G?�[Z�k��O���DB���k�BYJ����>G��~�!��a�y�2�4��ȉg#�p��[��vqF1 �uҵ�j��d�p�����{԰���~��/�{��? ��u�w��~��f�c=}��SxO�')��8[�|����9�NX�%J�ڜ�X�.�W�ԟV���4}8(�u��������RJ'�����X2k�K�STMo�_�P� �(�Z���r~���]΢�D�1w�]Ǡ�0���i���%˯�E�j(y��%q��;)��|u�|�g�g�p|���W�p�ɸIU�~�ӓ�A��Bî5���Vm��/���鏓����J�<��[1�{S��?H�ib���� m�(_�2�W��q���F~�BE*��t��y�$6��T$2�R�&�`~�T��n�@��l�w^��J@]���e6|�8kgg��x�;`kH lS�q��r�(�B���A9f�SrZ:�ƿ��K���r�ˉcf&q�]��cw��7kÃ�	�QK[?[`y����װ} ��Z���Y���{�����%؍��3�]:���}�{�k=����>߃nJ)����l�EZ��A~�K���SӒsU+Do�I8_F�a|9���l�����>�B�`�6e�����X:�0^V5�vp�}��Ls��]��гR��"��$� �:�b�J��ᵃ��{`���zͼ�ͳQ��,l��,�7�ȗy�f�d��c���Tv6�Y�����_�)�̵�*bd�D��}�W\���irYs���I��qɷ77fp}�6���Y��v���Y�����|��Le� E�6�<�(��Pb3�s������gbC����(}o��}�.��8���9������'���<����/���(��}�>/L\�>t�9�Is<BʤAN E��˕�kљ�����m�˴�<X��[+r6bO�u{�|�Ȇ�R<	k�|+����B/�ba�ﾒ�b��/Ě�	`ˏ+���7�-n�q�ȳà��\�{Ç��a%�TH��j�!�W-oig;�����=_hG^su�A3����I�{b����uTp��T`�B���5K1�痛S�����J�[�hYg���~��-��o���ч���g�n�#�Y���ȹ���O9|�v��V��F-��~��\��X�����>-߾/P�F��­`d<�5[�ձ�L?[��]�����l�����^tC���&n�HW����l��ݝ����=	O���=�A~�vx�/ڈ=pup�EX�+I�T�Cp�h��3��^�[�!�����O3�G�����5M����?qs�.��������"��]�C������ֹ��W��<��moUu��IN�	�0J��&�jFc�1��0I%�@B�@Ѷ6�Z
g ��OF��;6�Z��^���ڷ���i�|�L��!\0@��g� �� ��Zk��LB���}����9g�}����k��`��籪\^!��<s���VU��h��W�XU1����R^����xE&�*�VU�+�XU5��aU�x���0?I5sB1^Z�K�0_F�b��5A����׊B���=v�sO�ܓɼ���`^�{��'�ys&Ǐ_��3Z���J�1�ך�6��5�f]o�?�L�3�:S�6��?32��usM�ӕ�� h}��Z^�Wy��f(��,�ai�2Ǭ@I�r�;~`�B�[]�u�jB��銎�~�X�IM��%(��~D�ň�\i��L�ո��}�b�"������X1�1�d��з~�`�#������J[^��6��^G�!5L]��k*�&᪊r�=��?����� >�{+�� j�(y(m��Q��
_��O�����6����h�J[_�_��Ƴ�q�gmS7@-����wM�p��ncV	�A`j5�Xi�{��6�M���c� P�Z£��$v@i����h>�;��Go�3�����6����f���!6��۟���|�c��W�i�D��<K.���-�G]6�n�5�N�|������0qυM�KL�ԍ�z�H�4�#���)�I����ۆ>�!�e�5g��zCiz�޽QW���L��*��6��f���-t�
�<��Ǯ��n�5ww#���w�P�;�71�)b'y�JO�9e׹��IR��ax���{��Vؠ��8�� ��:��"�ʙ����|:ȣ����֞�=�(OrPJ:��~y5�w���]A�,'�*O`�0Y�>���A	����$SL�:G[�>&~�P�$�`T�3���o^&��׻����ߍWSL� b�����zWy�A���X	sR�	�S"ĳ$�*h�X�ݸ<"�����R2�?�9�NÜ˽J�,�dcz�ˣ�O���Y�[q|Pc}�'��/O�>1��� ��1�� ��i�	)�9�m�1��1_R���QS��l���~2� �������w��<���1��a�oӂd\��F ��>�9��t�Pu)V'��\�|����r���2�A��1C��y�R}��ҼH;Ϻ���d"�4v"�������v�~U:r��>X�K��7F1�L�t�E�kŪA؀,I�Q֩����	N����ۮ��-��?b�&..:����O�Uo���1���P�Q~�JPS\A�}��\���:ܟ�. ���rŜ�VgYt*6�${��2�Zo��.� �G�/> V|�h0�Ό��f+u{!�����hcZ��e��qmH��7|�X�ʭ4u�-������ǌ�?t0p�Q�6�����B�q㫸J�������)�c��O�j�P�ö�1��G�r+��
����[�)�܊��
*I�Hp!I2Zj$|��b�;pق��_𯾞����o_��&����;�5�FW��a 7���4��rq�]�9B��(-�26����T���Ŷ�-G��?�<~�N�+���hI�E�Qn=��hԣ�h�R�D�ߘq(��*�hP2:p,Jt|��o;��\�g`k6HcA�ġ�a�osw���V��m�������W!�O#�6#`����2E�_%�����Q<��0�htH5r(K�C������x��P,����k"�	A���G��l
�}����wPp�[2� �P@�r��4��j_���P�T�:G���H��f����'�w*�A�Q�{��Xd�uG�89~��*�
��iEd:�z��s�/|:������_)?��q�Q��7I>����W��B��XK;�5��c���c��cW�?v7\M�G"|�h#��T�^��aT���l/������܆G��jK�z�����'C ���q<h��&J��sl�2�׮V�A�k��<��é��������7coDW]����|��kB*��2CΏ"��$#`��'q�0�n�`ޚ@�����SG�̏�;�?b�E$�|�[��12Տ3|���Qe�h��d�[f���P�5/�J��"+b^grmPa:1�(/R1�y��t��i�d�r`.��E����@g*������K-�+�dɨ$��P�اUdP�T?o3���xJ$����D�r���?fq||�#����a�����/� ��l�;r�"x��>Y��&@s��J60�y7�i	!FG�,g��Oy��߮N�3���rM"�q�]�c�ᵤ呎^LG�V���3�T}-�C�¾E��ȕt����kG�>������1}K_�?_��l5�챲�͋�j5Rf�u�����x"�r�AO�а[�F|"P6��A��+scx���4A�v�>�a��`1X�k���W�<���}w<R��؞���?R�������7������h���F�c�B��'�7q(އ��k�~����GJ͎P6le�z#O�5�v�Xej���/s�C q�2���}�c�E�k�dQ_��?�"-�qnQZ�����CξȜ���Ж��K�O��%�������T���+��6��\��a��9ʮ9�\�À������W�7-���ڝ���������#`X3�"t��z�}C��*��?��m�`ڞ���̣��F�����'�z3����v=�Ȉ�z~��S�)��!�8��"��'�<���e:���n���.|u(D�$�W*x��6g;T1�[~��kBi��5I;-���4����	<&	{�@���5�bb��Vh贳]��RǙ�G��ff�#��3�U��r�i��Oxq (��4�����aj	l���Y�h$%����*Ѻ��2�f�)|7)�Wkz������{�'���tθ?������s5��h��m��gh��!q N��|����<r���	N`��e}�l"nv�=�Q@�5! �&�'��X'�L7N##׷�H���t0٤>.�w�����K����0�P��X�y���b�+�uiDu���V�g5_�ۥ�a��J���忣|!������3=��X���|Z��P|�����ҶS�QX�'�R/z3�I[��;��>L�a�Їp��T�B�!-���ڭ��q�a`:v9OY,pT�h��q��%z-3c~n�	6�˱�`4T�@��-��MZX��{Љ���~ ��a�od�yRg�9\1.[�����wO�l��!��rW���WʁEv���V����z���V��_���j��䭐wy{׉?���l�+����gf�r1+1?jL��3�]�w��'�-L���:� �S�^�:~7�C��������@S��}B���'W�-h�%��9�0;y��M z-|K�cE>d�ى�Op���.P|��5���M����D�β���qp�O��H{\�ٸ����f g��~��x���u�,���}��	!؇�o���&<�A;�*�#zծ���0��+���̹�
L��2۫jz8��-��*B���:#)�*�K�O_��l��Id��Og�Cl��8����-�x.�:ع�N38� gr/��8��JS����N!�^tS���L��Ͻ��
�C��܋��]��zq.*C�%��/�C]�/�g��N*�b7��拋��*���<������b\9k��J���/F��z�]PE��\1ﲐATݤ�E <��7u��n,ܬ�QKBr�y�eX��|^��.(��A�~��v<y5�h�K���6���WYC)����W٘'G���Wٙ'����We0O!�kE9��dw�ne����*�yU�XūrXŃW#�����_�\PL�b,j��^�bo�*h��'dE�`$�&>�%_ae�\��od��o��e��R����c��k��c�M����E ,�z���5��E�q��_)�hԔ=���&�����X�B�	��&���d��/��Y �|�W���w�C�yDn�n���:?�-�)lF<u~��@%#���"�X��hJvo$R�>!~6ψ�q��׉XZv��.h<4��@1� �pLC��O�Îf�h#��,�r$�x��fF3�OY��d�X~5v^�9'��Hj����nv��H��ω����꠽��u=C�&��Z��<�D�JP�I�Xз�X�)���-�_��} l!:x�cr��u^]b�Wg����}�Cȉ6� 뾾�aw�Aw֣q�S���tX��A�¿�l�<9^)�Z!?�����G�H�RI>�') �r���� >WR�����X�3�r�_*=�&�;��3��tGQsN��jT�EF�A�0O>���k&�����X�,�����#��wY%�Q�|V:
�Ry�<�#�&po3�÷D[Z����ٮ��Hy<����w!f���(�'zׇ�����Gv���g򹼼Rs��BnbS�a��>VZ��+���������Gpy�������	�Cz�=z=2�Ӏ%�P��J��J�r/�z�%�����#h>��(�+�9���s�%K	0?t���Q�W�����T��Ց�;0�D�y��f�O�QH�VQܹT��w�Qv�#!�`�pSF�r쭠�5����I�ю=�'W>O�3�2���j��̿@���v��ά�ň��,�.��~�����B1��$��f-��}S�������#KX��Ǭ�cx^�HJv'Ae���k�����B���~*w��$i���%��Mۺ>_Q<�^�4�#:���[~l�Й�є�w;F,�#��d<:���Ǡ��7�Yuf�:��avs�T������G�9'`��ͱX���g���}_.��`4�?�����L/�?x�d:�ҍ�Y_��:�D��:�n��a-OV�q�$A�itk�7���?�D�Mj��2�+�	FuX��Ld��s�Rd���&s��"����͎����ۅ$k�2�%J��:�����h�.�����p�#�M���A��@�ԇ�q�ŝQ�?Qp��G"3�c�ځ+�wc�m�M���Y���dI�ZF�&��+�����Sb�)�[�N���N_XjFڝ���ӛb��"X���;{�Ղ�s8��c����\
(��+g_�Ť�}�W�>K�֙**��M��v��'��ė�
�}S�f���әД�����8���L�$R ,���'p���F����@Q4��r_0��g�F��LGP�d�� ��Wa6hSl<�g� #������M;���?z�������b�\��pU&����E#0�&���*��U��8���M�ɚ��� ���yڪ���H�)>@�v_�itb<�vǌdA�ո%ۤ�h{�+��v�j�`�k�A+�[<���|-_����K1��R�/����22�Нr7��#)���Z�3,�����>f�(�����!R�Li91��*��xҜ�Ɏ�r$ܬ�К��s��h�a�{�Z��S�"P������u��f����;W}��y���M�����|�G�ϧ����qF���/�#ߙ	E��s�Nl]J��D*��u��.�K���er
�/H)�_��n/�?�~R��M�ڔ��6��4]��10����S]����I��O�����ڌ
8u���%�j�G-丘ŧ�����Ɂ�1o�f(HY�r����0}�^1�쁲��M�&���������&��}�$c��\�j�d��d�����ςe�ů��ha�'3j�Kx�='6��x+GT����{PH��8V�����\`�-n����K]�J�+h��v�P�5��Pr5�j&����x�?��/
�F���e}*�+̪if*�*u�e���zH��=2�]���OE�jɱ��w�߅�����<i߁c0S(Fב�?��[(.�̆%JJ���]93�;�.u�t �u&�p��T�=)��-��;g\��X���S:>���r��T�ْ�ЁN;�t�L�rzҁ��l��uOF/�6���gʣ�c�r(M�J�{v'����P�|��7K��n��w�G��Ї�=&��m�9����-��ʱ��}j�Ҷh�`��͊0��TÚ��������7���7Z�͍B�˃q{��^�[Bi�H:�}�&]T�$%`;���}*�:��JáT�r;+7cyf�Dyb"
��6f�i�u���D�	�-:xic ��0�.����-��.�~��HT豪%ξmK�I����/��^��p�k(�����Vew4`i��r����ՙ��hO.B���\5��������R�ɉx6�/[��-}�!v���[�����D��C���HI\��v���G�7���@�ԛ���%qo)��l��֚����0o)/�P�*Fxg9R��tx���VȾϠD䯉�h2�Yʂ�c��!�<C����9o�ܳ^b��;��va����ȳ+��.}$�I��&��"�ǘIh�,�ޠ�/�]s��>��#�W��"����s��%1gf�:LRV���:$:cD��o��.sdW�c����Ic����-t&��p0A��<5���00��]2�'�b���Y|%(�cb��&�=��BW3��rܞiq��"��K��Z�ሦ��96Z�v�����W�7�����x�t#����	)@ݿ?�v�dbՙDO�ǛY�=�y�w	�,�_�(^�۟̊rYy^�M.O�D$�g�r3[���m�g�zdL�%�0�����aT���ނE=[�}G��y+rW�Z�֘�֪{�zK�w���d+9�=vz\~9�"��{���tٕ+��l/��d؎yB��lA4�	�G�F�x%-�D���g�������0�!��&�!mNU������bB�H�K�[�O҃�/sJx���1��6��!D�Ay�K^��M�ԇ�׬�lM4�tL���MK�K�*hj��[-�os�-�M2"҈�^s��K(�8��N�~��~(����T����{�y3|3����y���հ�G2��z\,����x�#�o�������oxių%�6�0`;�<l��Z��,V����j&��p]T�Ң_y�+8	�߆��dow|��}(�QmP:x������+�Jey�us&4�����~lQ0�2�]Mc���P���)u�y�k]��Q�`��c���%Ⱥ�ރ�$�fJ�u��&y=������|�4f�~������.,��T6M�Aꏽ4�Q�^� ��)�O,�n13�@�U���a��@���Ҿ��B�~/�o�Ro�����Y	����@��$`��
V���;���7�@��F����� \��D}�0_"�ĉ6���&}���!����*K�4�ـ�6� ���9��c<�X<�*
Y@�m),�̘xB��_Á�<\ÐqL<ë�m��x�zk�����Ėb-+a�n�� �1�ZK�e$�� �
1x��D�V��(j��U��`V�4A6�0F�n��c�b�C�s������0:n�l�yF��x{�+�eT}ƲX#&{�?f�З�7��7����x���:�*	�.��!T��-D=����,�a�R�Qx���V!�]��k��w�v���%\W,�����+�,�%6��{Pw8#��v�.��mRZ�����c��3�U�l?���p�6��8�c�V#�:�����0~�8��H�����=������G��̬k�)	����@%Ƹ��ц��W��H:��oy�R!{WY��7�66�:���B6�}��a��U��ُ�_nav�|�-�Un6�NvcF�]X?}$�߉��ǲ���t�G���!|nځKO�i �hw`(����eJ�:QQh!
-(���B��C�_���
6��-��I�Pf>3ۊg��xޚu�>߸����(ǭ�;�ƙdM�_���"=�՟�L/D�pK�0[h��$�>KژA����vh���)ðl6�W�_3i,IR�g���E�L%6CKA�#u�� ���kҟA9�.W��łW���w�ڜM	��T?j�Y�OC�_�Wj�7D��;��,�f45�z��&��zMAb�l�QЂ<}�UJ[#*�d��$/���IBX�w�W(��rX�ʰw����1[B�?�%��&[�c������J�c����Y�����_9�֎��@i�xK%��
R�V���oט�QF륐$b7An�h'2����^C�]4mJs��.�H�W�Ȉ�+���
C;��YHiB�>�F�Gi��4�u��Z2j]�g�Y���-Y�a�%��-<���d���4� ���t��0�T�]:��v�W�҄Y�DtD��ïl�J{W��<��T|=�E�dcMK]����8��M-�C�1��Y���i�> >�� ��"��݄Tz���G�����pSD�mL�W{��s�e��'!©�A�^�-�8%��GH��e��[<�n�L��X	�@��~g%�纆�#�p������C������2�#��c��c�/�XhU���^!R\'~��b�,����e����-sp��0KI��\�ʖ�%z�l��{�\$����Rmش��kό�_���P��οFLʓ��wBA��_1_� ���$�jc8܈z��P� �i$��+����%��A�@��>`��'G���Mb��/~��uI��J����	NZ�%TKmq ��xKj������ �^�
ߊs�Z0W�9�q>�`C��A6���۶��3k�(�_{	�WQ�K�ڈ.���Dٻkw����������?<����%�������< 2z,]���0ȅ���e8��'0�1�+b��;F𰕂gB�L��.Zl_�ue<���B�}㈘/��,�&�&v��A2�;TE BSK�Pg���c�g1��b�O:4�׷!%[�ʰ<"���y�~�"3b���P�y���ދd� ���*V�����F}��W_�|�M}���1��^��¸|����ҝ�g��:4YC1��Ф^�32��涄��8���lR�'N��������aT�ٗ5PA���
*=�
+��T���6�E��\,#�on�R<��q�7�X�j������]�i��7��$ ���{m��y��("�0�f"�]���gB�;@8}�G^�A��]L��XOîГ��"a,�N؋1�Jo��ɴ\1���C�y�AM�j�Y�8L"�q*��F��+V�:���h;=<$���!Z�}�1�!�w~��R�k��t'��cԤ��(����P\�
�%S��q�2��M�[>��� m��yh��Џ��[r���z��Q�����ك+ԌwX�(!��
��'0���/��d�,rj�s,p�f��	Q6�	�0�����>��>ʤãrvU�����X3If��?$jT�Q��R���
-��f�X2Q������7f��؟��u�5;�����&==�������A{Ok�r��	��-�h��8՝�b`�o�����v��]��}�C�Ȯ�.P���{<�#m1�x/�@l�7���W�w�|�[I�lB"�� v#��w�]�+��(;�qi^�}���cW�ղ~�B4*|��<�p�7�����G0�B9f�4���L<*�ǧ����$/�ϸ/C����$3;b��b�]+E�!���4h4/�Ë��������?~��+��q�������7�N�������$��U��Xe�f<qdS������$Ԭ�?���Zx!�a���2�I��ye�Լrr����N��sym&�ZOY[˫�}n�T����\^����%��)�S/N�<GiG�}���Z�uM���n�Fi��VZ{�Vv��3k��M�ޓ@0���5#N3T�uڴh��F�_�zh�i�fy�Ӫ򮣾͍�9|��`|y1�����k�����R�"k�����"�,a��uK�q�<��0ck�C�k��>�MM��>�1���M� �pv��
]�v ����|��Sb�\^T�����~�#���,��*ߡU��x�JCc��q��ȏ�=�>��*1>�A��Դ��f��gQ�i�Tw�J�N�H��-3��S݀�_m�;w������Y � (ɾX���l=4�/��M@K*��L��9��[�ޗ��a���hx��8��-�@�:G>aO����F�XH!^i��o��U`�C���y��/r��!�r�E�xu���9��4ps��]+~̩�F���>��`[�ט�G�ۉN4Y�h����@M C�RM��6dj�Y�n�Y^ᆭ���2���z{����0����|��$T��l���&���Ob�؀u�p#(x� ��|<O�����lKF�\�hvϊA�n4���Z{���ֳ-�3��>�����<��zi���C�2r�<���3���J
y��)>[ˣ1K����1�$�U1��[D�3�����lXw�Ov�7��O��C����(�����ߒ>��0��H{]�(6>Cy����|@b��?J@"��޴I�%�aL�?M��?�/$�1�8��<�?a5L|wý�#������9
�,W���N���˔d7���:��x�e:�����3YuX��=���cߓ>�+sw�G��s�?ީ�h���s���F�\uZ�1+��}G"*���y��K{7�j�E��Lv"��ͦ�
,'U����绑yQ^�E{����X��Va��a<����0�̨߸V��Y� ����y:�"��D}��J�v��Xդ]h@�bL*4�e��lgAP>0P;�Z|�2�����p�"4��a�G�`��@@N3o,�e�x��@59|�������4F�3^m��<�1�r�գt�;O��%�OC�����T�&��Pc�Q5o����9���O&^"�5tJ��)���p3��a(����N�W��}�?y=�'��N�Z&�'0��<'Թ���4��
N���x�;��������xO�O[���
��Ç�i�ZF؀��]Z��Y	|�2����!�$�Ԏ�U�ٳ�o5���|���!��"�L����G��bIj	<@`x_Cz�V�7ṁ���AÍ4��v��-s}]f� H1��p�Y���~�XA����O�d[>ƃ�n�G*�~���c�C�"P�������T��m��`��ށ�y��گ-�nB���=LO�a;�$�bM�g�4ϰ`+n;�I1��`U�$J�*�8{1����19�����	Vw�8�w��W�5G�!���,D���G,B�e+�oIcQ�\*�>#ph�	#V?:!1�����	��	b��GTA���6��v�9���Ag����at��r�1c
�ѭ�l���=Dd-<M�9m������q�/��x��8����'G1Ch��<����bTk|؝gõZ��]����tm�U�f��S��.��� x�uBi�g5˳)�5Q(O����8�6+;K�*L�qjs̣��}rtyo�!1�۴�$�K��Xw��p�/F/�nt]����t���^ �V^%��X����y���[�B+_fC�m��:��:��=��otO���lBG��6�7���wCK]�j%�g�7����7釙=�K?,����P��~�س�v��I����ˬ��>�/]_
�z<C4[� ��B�������]�A��&�Sk�L�����F%�$���Dx�)Z�U�N�o���&�(�nQ,������צ�
��k<�F��LɄ�*
D*�hBD�Ar}�o����6(�?~�"��,��	��C�	�c�Y½�0���j<x8��<���3��2��TN�D�&fOU����=���h��";�˙�R�e>�9b#zut.����8׀ݚ�׎j�8�
��8ćGs%��d[þ��[��Ӏ]��� Ke���T2��[��V~��ӄ19��x�rǸ���_i+7o;����4���G��C��<���`�ɑ-��ډD.�^`�߆����m#S�w���v�ɗzcy>���K�g��*����AS|�(�r���Wa;�#Ey��*�uw�Ȋ5��&6�-��p,�$������Y�c�{�W;��y���/���F�c3��.�m�e���	忑�Ua�&S�tm�X�{|if�?&Џxyy������V0�K3��J
+�?!?���rz��I�s����=���Q<�"�u\v�tX���*����n ���u*ŝ�x�$�	s�i{�`��{�muuS�E�NXuf�q�+�d���:���g���҈Lf�2���ձ|Ŧ������W47q���1��_���M�*�,��u�s��}-����ȯ/t%���
�,4a�	j����T_�<�/@����0��P�Xۋ�v�J���J��+��sK��[b�x�+�;��0ڹĎ��%�\����%foWv{�a3Î��N�ކ�H�O�ry���&�w�����x��,H��� �9�"!c�ɵ���c��`�	��|}��?XE�N$� ,u��Ƴ5�/0�s�"i�TI����5��s!�m�{���5=�C�Ie\6"�CE�EB���ZÊ젱m�dU3�+�F��t����X@�O� 1{0{�yI��OT�GY�4.ŒBe�r�b;���,����K��)�G����7;^���{�}������'L�,��X�]T�ѕ�?��䗣��םHϰ��X�W����g�v�s�yT�^D�b���,�������w��!qcXZ�FflJ�}u<��,�K�F2*�+M��@l�%6֏AD��A�d���/�o��^���+�i����س�gW�OxAU�*�1����|	ji/%Y՟EX���$��T�r�Q�+oΈ�&�|�/��.Ϊ#e(��@�����ߧ4c����'����VeW��#޴=����{<�G\��(MO��-~F?L��Ï_:H6C����0;��VH��1:���F�Eܿ�TO�0��D�>d+2A{&Y����V��|�l�������`��Q�Z��R�1� M��%����-�r�F���]#3�A�����] Z�t���.m�`:�3-*�Hx���*��A�E���J�F!T��)��?S3��
�~�s`t�bU���|X4��8�N)���>�f�F��R��G<�Ś�[{i�f���ϔVkS�:Ki�SZ���VB[���3h�� Jke�K������RP�>�N�S���׮�s$r���Y�Ť4�B�=���"xxxxxxx�-v�	�d�ϟӁ��ޅ� Y��PA��YX�-J����k��q��R#�(��"6dL/�㍘Ҩ4a�_4b��DH�IJӋ�K�=h��u	�`Aԩ��l=H����2\��m	|A�3�S`=��C��7퇗�tr���
S�ע�z�"���ک�檩Jk�T�TRzo�w*�Xa���תm��^ #��W ��g��D~�ڰ�<�y.�t*�w���n�:�"�8��bt���"U%є�$������d�1�i$��I�މH��P�1v0���3���:��)�E"��z�L�sQ�dR�E�q�{�9W[�K䮌�����M	�rxE.ܺ!^*�-ȅ����T�T�24�(OMf���xEa�M
L���W��V{r�u��-�u���[�V�<��"���O~R���\�W�%x�1<�R�˓;N�Pu�2o�0QA��(I'��`~��0��
�/�F�F��
��v��z-�b�.�^�&-����u{�:JV��g���U��XS�ڒ��>�ln��&�O�|g�D#fO8E&�[���jv;���7�}���� h��ω�@)bf��?����щt���T�D`4"�F$?�_��ٔ\GG�cj;���f��[�mF�F��s������<l�������n߼�=f^�i�Q��R����<�8� =��L�]����Q�ox>��n�ДI�������1�A�A|�J �Iڞ��|�����#^eq"XM�����T���J�$l��[�Q�h���h��ϵz�4�o�)|����;(g���Nh����=I�F�9g�i��WT�Ц�2(�����,�-�zY��p�^j�ɤ��Ѣ�r��"��
�����4�M(�:~���	�$�d��z��J�b����)0��N�>M���9�KxT��;�ٽD�(��!�Ea�,jZ���[��Ȉ�aL�l�[�W���_p�����񐿽X^�P��/E�����;��K���HfI�6�SW#a��[��T�ԛ��́f���T��Fa�L .|ta��k�i�Is4��� �&�
7i'/�������.��Sf��mU�{{v�x�)f�b`.x�`USj4�C�ĸP���|+r�����gH�e��H�E!��rO>�P ��K�ѧFn�x���9c�w\4Ul��2\�6�Y#�����m����go��}�A�il67�K�!Ԃf� ���&{�,��v��"���c �\�?0o���J�y���w-��N6t�LK�e���ē�u}R�{W���h�]-��^C�<$��Si;�E1� ��8�� ~����;�i�^�v���'��W/���U�nPv�(�{�;]G���:Z_�а"��(��~e���F'�u�k8���:����#�\i��;��Z:�0K�]-���7|tWT ����rg��5ڨH5[�Nٽ�<��/5&SMǰ���t\L��� �Xj��*�� 	;��@�T�G�w�5�Ť�;��BJz�}nh )��h�f��g����/;�у'��2���������Eν����9���<C�:����sX��l�������"?�����U�w�ہF�rB�������L�vs�`�R�¦�E�	�ԬP�[�4L�	ýrh���̼���1�:�oH���2 �c�|%z���q��/�ҁ�����[�=�J�~���M{�ٷ�,}�.آGI>�
,7��x����R�Y��<Q��gv�2�խ<��,�aI�n	ڼ�y���uTi�����6I�ހL�F�>���z�]{Tb�Q����Z/!ϸ�oC�,�� ։���!����]��f`��)CM�2�Qk�o�����;��x��lWZ��@��2)�t�XJσ��8�A9���s��о�����̎DZ)�z�@�J�,g;&i�S�%�(r[;`v����
a����N /�X0����P[/�������B�^�h_(����́��`�,��}hvU�r�`����lIp��y?ZG�,�!oa��#����>���3x��9�?�~9ҙ�Cq�1�А �Ę �	=4���U�y!�z�W��,h��m`j�@�o/24:Υ����?�����c�<E�%�:gh�w�=�˨��p��K���=�$��
zr��U��ۛ��NfG�8��#�����*��a�w�ˏ��@NC��X�@�^AQ�"�A[���p>�=��2g�R���Toe���B8j�D*j�#zH`�	S�3���,g;�b����m
�E��Ev���
��c�0�lb���dm�����U�v�� ��}I�����S����`̞/�Ѡ۞�K!�#����� zv��-�h[�ǌ��W��|Fcm�I=�$�,�O3�'�6.������˳�vݍ	>%r��}�l�Uk��37��1��?��;�7[���bԲ!���=��]=k�r"�X�I��MtN�Bɖ/� +�"+�"���|��՚�!	Z:���P�&�9�>�y��&��MQC�C�GR^]f�����H�o���+nq��Hϴ/:D���Yd��
E��o�G-�3S�8��� 5�\��p��;�HJz<�i�}���, "�&�����%oOh�`�^��l�/a��7��̫m��SM�5���[�E75�'kk��<���<m�`��S�:*�}v���@7�pOn��\��T��r+w[]ݾA�[H�ɒ`����@V�����c��
:�(�����n ��Za�<���U����ZmgE6m�C
�- ���M�3V��"�S�#�Z����I���!�6�
w�_�~��Q�;�׊�ei���:(��H�����`�	�˓���q��[o���~
�4�fMK<~#�G�׺��� >�Ǭ_�]�-�����j`�wy	�ߵ�$-�H��1�E��)!�������}q�;�C��%ϯ���<�ccU��9%��U�rЯ�D��!�LT<��sf7�~d�z�u'̏17|	�6�$X�`�������
y�
��5����|��7�d��}��F>�$ce���{���R̡g�v�Q6.h|�F911�?���3�W\37(�̤},�#[ܘ9��+��Jk�4����[�8�/��f��c~�-�1�5��b�E}�)��E��K2>��׭�.���aDV�G^k��Yh��$!(���o�bq�O��(��8L,�|���ka��$#�D؏݅��V��+��E�;M �qIXv)Իw'�4<��ʞ~Ɣ��N�I2ݍ�(�{#���,^[h���BJ����������?�B!E����9GYo�>��;��*)嚝���r0�D6�hy�D����?G��.ᅎ>��.�?o�U�~B�軸�<�~,Ui�Bޠ�X��~/�z}Rx
���(�k���H��kX���-V�BY7"[���3�;L(-�"��@j�ed���~�_E��YnCwy���5t��2?�j-n#&���p��5��p��@Q�Qn�X��?2pŌ%˒ȴbg&�sPއi/�(�i$�g<A�ʥl�&����L �ۍ��U���4��)C?�!?4<,5��Q#�k��޼4x{&zZw��;�p�Rf��2(%N&�}��!v8=H:MȜ�WP�x!Erd��0FGd�9<�m�'���-*S~T��R�*I�`�LG�
�wTT��)O�� Jw\CB`	xMkVH�ѥ�ס�g	����y��9f�kߦ����a�kւf��Qa�~y��[Ew֐]���S�͒�:-d��(�?�N��<5�EO.�i�g޼>�����`:<����������Xʶ�E��u�xf�:κ'E�7^�� �Cv�[�i�����7��a;p�:�N+�ߏ��}d_��<����5dC���+��-�T��܀����l�ݎP���v?���2��,:/R�i'����X �R���2{��ߢ�'>��.>�{k[T���u�Q��?�?K��a�ߍo� G��`z�%4_��?㐱��p�h����4�:g���[c�K�D���ͱr������'h��XZ�=�1;�D(P@b�a�z*�X���Q��L�s���7]_+3�f��~��f��fp��F��.����ѥ��a����|P@�j��J��S��^�dv�x������C���N�9���6S��>�y���-)bg�%�DlI~�7�I���|�{](S�<$�/u!93b����VC
���2�\���?A��C�	�~����=l�2˄U@��X�g��%k�p�ʠ�����Ӎ[d��	�2����6�h�M�N�hÒ:�ot�TxnA��\�f�>h�=��@���Rի�����l	z��D>J�_��h���U�e�^�.q�NK��`�_`F&�(�ݰ��%B�H�
J�u'������*��}���Zx�4��ڋ&�q�?��� D�`��8O!�J���+n�	{T����־^_�<��� �y�5�/J,��1ׄܰ��Kk�J��\)�uJ��F��^t��e�&P����7ԧ�Jj��O!;�p��Q�b:��.'��[;/J���*�wRl�d��kQ8M�9���R�*<�����5ڞu];qM��|&`�|_�](���L��^���Lr��$%YD�#G��_����V��-_����OC?A1�[3�z��)�pY�fq=r�o�v���j(P����I� |4��|;���\z��%��X�	���AX|&���{>*�e��Hc���ctu�����d�:�^$&JȎntA���O뼒@�y�.3�6$��lS��U�W���x��q�]�d��h�pXzE�(g�`l���d�P�B�q���<�-|��-SL��S��"?��>4?^��o����v>�Vx�;ER��7Z@/��_Qn��r�CFUL�Y ݏ��"�f\`�1���&u��H�����]�9���_����_��'�d�^n�hM���m�s4K�*/���r~"P>��������j,�v�� ,[7��X񗝃1����c�?���+Q�$�<k��k���/�Ot���gq{#��,rیҷ�N���w�I�?O�_�X�����L���>t���q��,�g�5� Oa&fO��A�~���/�qqD�	���9����گ _Vڊfi'/a@^�,�/�ʳh"�ƲQ�v�u�X4r������ٗ�߇�r�e�%�CgԷ��=蝕�����}M�	�ב1*�v�:�k�k�^6����l��y�&)�x�;�F��D��U�i4�Rޡ=���z��U�i9�;7K(;����.=����hG%Z�">�������� R�,�U���._�Pw���Xoi1%+����Cn�Q���m2�s����ͅ6w�7w"��R|�bE.��3~#X�Ǽ��7��X� �����݉r�y ��Wږe&�r� z�_�H�-��ݙ���p�^�C�y���-Th��N���O��#�D>���kH6ԨU�Ȓ��w�ټ�k��b������Y�
bʌ*�-|�H6/��JitTa�U5���.��>_��P����"�����:4a�*��^iQ��ja}��ٗ=<tNq�:����&כ�c��-5�~��]Ro�8V�5��
uEz'���Ap�(�s)�r/
�ڥ�M7����@����K��j�x/8����h�����p��xL�H��M��vLzLڐ-B��9�J������� D*9�XRZWK�/:Ӯ?��ӡ�c�����U�l~^��J�b�!&��Ns�Iszf9�$�y<��U_� ��2�ee�uMqumΚ��lL���&�p:�S��h��JI��-��CYp�/�S�*,�O ��C��q��R�dc�#O���8�D�*��,CEY�TZ��a��cf�dC$��5�q��v)�S:��F����M=�����M�'�!�3���̛ͪs�C�^M�Bӽ���m����-��[��:dh�44�2������'�6�U�e����h�M�`��
~c%~cl�8����J�=�~m�o"v�dڜX����x2���E���!>H��K��<ԇ��_�{DƯF[4+)r�%ׯF�~�%S|l����s��{�#�O�N���i��Q$�*`�*����?ZA;��w����i�x$exՙ�'��9��9fc�مG�����X������s����Y"?���:���<�;��hۏ���h	��.��.�.k{�D~6gT{o�z�W[h~*��=e�e
s�~b.�j��V�O��V�l;Oa]:��X2�^3��kn2�"��1��et4E?�gЍW8�T���r�`��7w�S�]�����:�1ʟ'��2}�D��Q����#c�1vD4����(F�P��|>r�g���3��b��h܄�Yh�ۏ�;v��QECrq���H��V��'�2c�4����8��؆^���o(�vQ���;����SJ���5�阚C����v's�@����+mI��J��@31�v}�o���
���/F�#O��(/OU�k'��@ǐt/�b
B{{�x�{TϘC����S�_����0,�9Pa1��������GW~h� k��n
�u�� &�rc]�9+5b�Ds8�7/��|z��v����h �yf�?z��mY��q�F^|,S��dJ ^�g"�	pĢ}��:����Y��yH��I|i���Z�^H��2:&�5�`}���u�������ht�?M��:1���.�e;$���:�;�w�G�_�O\t��n�-���y�9�N���f3f���6�Mv�sj���v�++��Q �����x��a�m�]����"Zx>F.(��fi܈�1��Ҁ��6��
k
��~%k��2%���������eG���N��@��������)�U\^xI�AˏdpY��O�����Z�]�\~x��H1���N�����B1�_L��� �9���� ���?��]ֆtLo.�a��[~�|�\f����8��1p��G ���������m���Ro҆1:�#�m�$(I��B�$3@�p����b����
=��"'$}��<�[��1���h@�i#��-�B䩖X�� ��FSʙ��p�����;���K1*/;��w�I��KܓC��oA3��m�x��J�#G��W��#���M��!�H���/P�(y*F1{� �
�� J��6����S\Ur�e�-|��'i�INh��,���ɏ�Z@ ���k����XD�K2I�p
���d��m�?�?
�U�D�d�ټ��c2�}�3�2�C~�F'��ԃ`�+�ُ҄�>�w��u7��1c���i#��)�K�$�p�9���R�K(���|��Of�7��	�0���[��Ks��!탴Ƒ(�EJ�'@j)§%��O��w��Sq���]�`9d�\u��9*�����0C��[���4,�dg{䵚�W��U_.#\���WJ�%�Y'��}�8�&��c��6��P�iߵ
�ָH���1���=�,�*��� _��s�K<�˗��U�x�Ɨ��ĳ_�en��W?�L��z#����ZPU0%�~�P1��G�M�T�H���#=��^��<�Y5���������gf��!����wd�x<�I�m�W[�j�Y���_�>�N'M�TcГ���@��]I&���p_��B7D~�(efü¦^�K�@���n�10��G��q��i��i�&>�o����D�jA��:�P]\T�^��71����u�ڥ��H�;��p���P��ֵ'�R���������WgY��}����'Tl�w��E�����^{�*p�ɵ�S$����g{���l~;_!Ӿ�9h�LG�.��c��r�٘z$ο&�&z�N4���S�w�ϱY1���f��<�+I�V�<�|�����VQ�/�9��9��K�Fm3�xem>�X?�p{ka������@19/P�D&;�V�s"��@�$����O���[��f����5n�k?Rl��'���=M��Ƨ��O�����p@��<���HÑg�ӭ�BY�x��p�<��-�h}���Q�2Eˬ��))��l�is]�@$@3��x$#�Kؿ�)��.�oG�]�4���by:�D�Ԣ�o4�G�Ct�g�P�p��n3��]Z���?���'a���d)v��Z��5�?�ؿ�Cr���]�2���_���������5���'��,t���O�M5J&�V|!��)�7TB}~��[��|2�'̔hXVb�
y3�u��0�W�V(Dܣ(�?f�G�G�N������8�H�5��F�kt���!p�i#S|g��Q��@�oM|�C�U-�k�"�z��g��m� R�"+/]�6�l�3��!k:R��j�[]��E�&,����`a�Z��܄�U�B+��|wQ��<�@Z0��S��p����M�܄�~g�kE�:Wk�\ݾs��,��q�gj�Ҽ��E�y�M��՚.5̀��ŏۻxQ)�J'���?���\�ŴͷJ���8�b�
�X�k����SvAi}�U6�URs���.H�����df�]����G����ֹ��R4�IGa���,)�@	Z_y���{((���|1�Ԭ���X
5u�Җ���z�;��5����	�8��xJ�S��4�}�W;�9;?o�HRZ{Ȓ��d���ک$���}Tψ��G�6O��$���֞���e˝�*�`��1讵d�b�X��c'8f9����7���q+�K;{�f�QimFw���<���R��|�s6��m� �2��m���R.�~������9~�V4�`�1�Ѻ�����e�<'�J������:�m&�z�.�t��T�v��3k>����Ρ���X������֕�5���?�n����є�Ǹ�೘�濞1 d����p;X����VÖ'q�Hp���	#��l�=��=���� �x@��M�>���3��c,=3��c�J;�����t�����w��:��w�I���Y`�+la��&1+Q�&�B�!`$\"�V�"Њ0�EB�]e<���R[�*_۾V�j�D�@��BRnꫳ,(�!@��<ϙ�l��}$;s��9g���~��!l�2 �R��Z�"��C0�<��E�o�8^��jKl�0�?���4K��y�Ϧ�Ef{����l��e+��k��X�m�8�8}�ȕ��4+�7����Lk|���\���Qv�l��&{ٕJC�v����!#E戦���߼c�t"��}.߲�덓
�1�\i&���_y4����D/��6^�G��v�Gl��'酆�D��9�V.3��D����y==�LV�#?��0{��r�Pu���菿��0�P!s�u}��ƅ>��a���G�ӝ��&��pZ�ԝ��N+������d",�C?v4�d��@T���h?�i)�ײݍz���_Vk�d�&�s7$�� ���2�C�Y�CF{�03�P���1�{�=�0�����K� ���=Nm�������z�������0��M��O�c����#ک��"�燴a+��і��M�����g��ݱh�����c�l�X�~�)�R��հ�G0�Co�11y�M��0΀@Æ	#��X��˹��iP�nf��0���߮��y�}�����`���@�-���l$��헗?�|�;�s�\�+�[{����+�w�e!���	Sp�C�3q0̀t�"�螔bf�l��%��>�)`q�-I��;��.��Tl1���۫��c���B���9�'����Up{���Ciu�C�z�R����8g��\$�2�wAP�VH��.�f'�pe�1�mJ�O���/��}�����<�W_	�y�ڥ  �% *�,$`��rtϯ�*����;�Ø�����g�N=��J]�z�f�٬�C��Խ�^B�c0����J��كaυ������x��`>�ҭ�p^$��۪'p<�21,�5|���F��b��X^�%��3�c�-.3��ӧzs�<�D�IC퀧G��ʻ:�Dw��^$ߌ�E���9L���۽�Y!��A@�Sڢߣ=!������lz&�����a�!���z<�}l�ÚCk��Q[<�r�&������PעF]�$7<=�*;
�����]�}��X�M� m�fJ����p�/hS�)2��6}G�f�l�@%�~\�9�|�Uz{�T��-(}18r�Q�B��I�����=4m�I��d'����@�%Y��DQ_�oQ�a�m(=1X.�r�e���9&mZ>����j%�)&�f7{�F�K�l��e�Q��%��L{�v���!K2��F���gK���Ѷ7a����X80���d��\�#����x�('��� ��ɛ�tM�WlOm}�g�<� VW[xx���t����M>k%6u/��R�H���W����g�^�??.?��s� _��+J�;�����-���6�;�R�l>R�F}�kdV�g_��!�ʱ��R�z{g"P敍�f��m,�� j�������$mF�@��M�9�=mU�b�T[d!bF
Ez�u��EM�L��m���o���1�^)�k��M:�
4��X�1��k�ֽwK���>$zݍH�Ԭ&���hZV[V��Q������/FH�X�?<ZTY'�os1��	R��G!������)p��t
�G�#)G�R�������U��-$������9��xz#S�E����!�O�T�R=���s�ů��Sj�����b������꛺�(�Ƶ�"��
���z<�.��WP�x"E%u/��K�sc�.ٹ�q[h�P����Kz�Rt��C|��$AG	nX/��:Zܚԛ�-&T�՝j/�O-Ae�ť��F��c�y���R���L�+~\5�V���#̡{����W�J��?��S>����V��h�B�A��%�ׁ:53Zf �-շ�\/�o^N�H�ȿ�H�;E�����^��l���i�C���?Y�;.d�s��2��$���>�#՗�!���'yN{����ٱ�|�d:NiN��v?>�HՓ�'éAj�P�kl|#aAv���m�C�W���
��R�S�dN(�O]Y���;'Ճ�~�����>3�*H�����@F�M��?y����률�^{��,N
�&�jhQR�7̲�����	�0����#�g��o���wvm���+�V��p'��v��Z�g�bW�����6P��MwB��E��J�͈��[�,��/4��-��Ƴ���$�B�G}L��_.P�c��q:�%�0"^�J����k����=���©����J��W�Bd�\T� [�' �(�҈\���é��[����{��*)�K�o���yC����
�����������c��㯾y>�{�g��c�%�#�b��!����0a׈I��=�zo����amU� �����M(��E|�m�	j|�F,�]~����)ح��IK����<��>�W�1��,,����}r���F)0�^��sz��'�J/����ҋ�ڳ�rz���R�m���|�_�H� 9>Đ:�\��6q��0���є����A���}�_��|8�OD���N��6H��"��z|�p���oc�����W�,~_�K�Dw�r�"����k����f��b�Pg`#��y�z���o+�7`�I������Y�����k�]�S�}H��©��;�ǧ�fJ����h�қ%_�~$�ϴ���C�0�����@3����S?���͜x���n���4j�,S�s��f��~ٵ���:�"W{���T��]��G9'֤��݅B&��0lm�6wW��[���n?A���Z=�Q�1�L������9N.d��v�l~�����K�U_ĂB��/G���[��R�Ǖ��������G�����2m�[��&k!4���
z,���q����`S����8��;�H�i�����X�]�Qm������f�	I����;[n<����+�cS�~���1g�E�_������ �'�~G�|����;���$Q@\�?� ���6���5�h��?�v��C�5���*U�L̚�Vث'3�퓏/N?��=��a�Depmq��XC��HG�2�N�K/4�V�"?�:�������:�v5�[�|#.�A0Z0��d��S�d��jA�+6�0�v ���	���E�e�K�Ų�Z���b�k�g䪡��M;�x3&��+jS�8�p"�ί2����ݬ�R}����ZZ�ʇ�=�.V_n�UٮO�`CX9�_'XO��ā*��pi��y)��\/x`���]����5��)�],?�����񣁟���o�|�?��	�pIL��Uޖ����7Fw���ux��(���r�F��߽�Y�����w~kq�jtK�y�u@,��6��>�L��k&��^�#[X^�1����Mj�+���Vw�����h�z$}φ��r��+p)Gk�q	>�%M��K�q\~XA�5�L�C9"�$����$�/��E�y���K"ak���5�v)8��cȞB���]��+��B�YlE��P��a@#E^�d�j���9�y9��ϡT)���� (}Ãذ����O�s���-�K<{�*�;��o��K
`)������)����o!��)��B�a(C5t�M�U!Q��Yݣ"s��+E��w |.��-"[��nk�1�Vm��Ԗ�|T�x<��7\z���� ���6����C��}p���ԏ�ظ�]�����ݒ~X
���h������9K翂�$��Zw!�S�3Խ�őJo����'�{}7����������0xE8x�54p�[����Y�gbى��'�Rc�d�w;1�~�w�w@cPt�xێ�O���c�ի���n�ۍ�+�q�^�/�]W�v������u�h1�%N(���M^�xP0Q A[u3�JId�
��Ť/�/��� |B򿇾{�|�w��=�=���	��~�� 4��.z��@Y_g&�Vr�D���:ޡn���?�"��dX���8.>�`}��D.��D�xJ\�R�1�n�r� ؙ޵�Z�yo���p�́dh_V��K�v�K{�`�	�
�:	_ �zU�8�/EB3
?_
�F4�t7xfB�{C3����1|��%��.��st��*�yм=�3=���	�j��P'jH��vW�����҂ܾ�"�c$"�7�LCg���Y�LW�� ]]��G��*�����������55�7��/�!��@�<R��*m��MS�/Vz����ǘ���R����0��4���	5Ym���|w�Z��.m��Q� x+�����jkv7��;��c4]���C��S�k�M����x���n�d��7i���d��:�AT~t8bKxr��L�����mj<̓��%��|C�#�E����/��z~��8��R��2 ��<��}�e��rY�����fw�f���R}r�*�V�Z���-�B����)��6�Iځd��{�E�Ow ���l�O�x�-e���+�R�+����]�n����P��V���$��P��C��{��L��&Os���W����^u�@�GP�"�M��@_&�Go{��=\j��%j���c{j�^��۳�?���K��p���&��h����7 %t5<5����?�F����{]�'8ӛ�q�l��v�}�b5.�s�R�p_��Д;��1R�����^2|=�OSw��5z�����֞���F���?F���{����]���|5�B�sV��Cu��©�_�!�`��)C�.�I=ꔊ���>cO�^$m�/�o���o�f\ⲐiG�S��Z�¶vxl,&���A��[k���������<P{־2�����B��x��+�<�g`�����P�J�FccO
>c�������&����A GX�ݟ	���v�Uҏ&��K6k�d��=dIn��s����S��fՕ�翋�5eꞜ�Ư����?���E�n�m�6�ᚌ�m������ӏ/^	͍yWG��{�i�g�Z�6Hh�4J���D�e�
4����lJ�:?���y`�V��t )��������[�odk-��b0W�BSOg�Ȑm��i��1�qhF�/�5_b#:��t��s��iT_��,�Ou:�Syk&ax�짢�$�;�т%�F#���N�8k�0E�W�S��j��*�S�/E��L)x�<���SҀR�oV��n 
��(�ƨ}�H��n�K��s��08�r�ճ�jj��7�\6�J"��~��Z�_4�Q�M��{�� �fۥ�ǒ����'&55alչ!�Mi��ex#0�6�zid��`>{h������IJ��>[W����|�����LB<�H����V�I7ſ�3��:�|V��8[����~���X�Ww������e���C��N���(�
�]��(v����D���myh�i��L\^���@��Ym<d��PRWD73Zu}g+zs�rX5z���ʛ`�|�/���RaK4���Pǡ����)&���bG~KNf��5���z����2�`;5w{txg��,�3 �p��v����@������ǝ�@{�فv���y�v�r����#��,M�*�A�,�4���E}�*t{NW��e"��{�OlJg�s�H��C��x�|����9���؍� ��S����Ш8��e�'q�8��}04�����j�����=��[K��w�����fn.��0�gd'7�t���$�P�-zm�Ds�3�U;'��>Q��U�<h�"d	R���^_[�%���Ck�����y�\R���?&G'�h�6Ji��\�Ҟ���SEG��_��>�SNi�S8�<Oi(/��A�`��˗�Q|�j�`AW���$]���I���]��x�f�ݭ!����$�/NV{a�����Vp�p"�.4j��[=)Th#^^*'W�^.�ނ�ݲ�P�nriB�izmp"*����M6��1�9h%��œ�%�\�� �ZYZ����.�&�iT��Y6�=��C_eǎ����oJ�v�ʹD��MT�N�!?��y.��,i*1�V9H*���T���w�������W��+��ύQ3�rQ-v����7�������C�����	�ϸ�u��`ը�C��˾b9�5�V��p��P�o(�٦�Q��y���&Ϸ+?��� �b,a� rQ�`�,�r�	���c%�`e��M��|��$�Ž.\pq#d�Aaz,�#��h�l>��cYM��:�{�	����ܛm<!��e�t���{Ũ��_r�kx!R:�G��xC��
H�k���`�g���ѝ����Gܼ٧6[�)�s!��%&��!��O>��7x�H��b�j?#�Ҧ��w
r��A��d#fPh	�9d��ⷓ?��N���/ȑO�_�N��j.y!ڥ�1\Y�~+m�C��xLTϩh���I��Nl<���y
�͐�3�kV������rQ%�p�S([/��tBtA<��I '�	"�C��P^�G�XhbnZ�W"��o�&��'y�<) �cH�yzv*��r���L�٠�^/a&��s]�C�I ������J�V���{o�va�<�i�Q�S3�zbm�hb��u8<���-n�}��g}t�W��b�~xm��[�*;~<5�I�PxT�p���ܒ��@/�����@gk��rk���'9� _Y���G��|��A��K����5~�n�{?^�+X����*Lֶ߆��M�T}�����ը��q������M��[��.��{#��1�^��q��{V#�L�e�n�������/+�T�%k#�8��\ɪ�`L^���,GsT{U����|��N��e�:�L��:���'�@iS�8�عS�]�+�Am��0�"+��Ju�uD�]��E�9�2+34�:4M*&>�����m�h��UEdF?��}�0��?D�Ǐ꒷b��sH�C���T�KBl�b�<�"`��:i��a�=�ɟ_��y�
Wz���M�[W��Ļ�1$6J[K3��W<�r��u�x4��ȡh����*�+af�}�X�m�R�Y�~�qT�D�y��Y.,�c�����]�>�ebRQ����U�[�?��׼ڣ����0����@��2��PhZfs7Pׯuh���aW�Ɩ9<-j�sՐ��,ёx��h&��
�-�`��Y�%��zU�-����sd'����PEיP�A��
�]�Z�B�!bC�S�v�B�ޟ75Bx���;��P���?OJ�+�{Ÿ���bC�I��c�PWE�F����@�=��(���I�fds�G ��.�O,*}��4�G���$�&�� ��?)���l�"C��UmO3���Pa��I��#�y�Kr�����F�॰vw0o6�C��D�s�+O.`Ӑ��c�1\rm�Mj����C�@��&u�x٘�����3	�葌:�#�7\��7�~��1�D�R�3���ceW����4����Y�d��������T�gI�����e���D�����kuW� =�|�:i���I.de��|�i&Re��/���7�;�L�8��?��
U�|'M�N=�}��}<�R�ړՑ�]�$����t|WWM4����d��xFfn���O��Bǌ�a��=P�T5���=[�6���ƽ��I����"��J�G�1�3#j ��3���ᇑ0��C?���E���Y�3I�o�8�����&H� � ,g9���21T��vsg_�ݎ�`����.5M�#�5_)�6�X�sDw7�?��!C]D�o���r���'Ś�N#ekV���r�\S����أ\�gj�o�����
Kv���� UI3�~���,ơo&[Y���<y�K�;��'C+������'vQ��lr�7K�7Ɲ�P��<.���a&�6K\�Z9�|�e��J�� ��� �s�ɮ�������M�����F���O�=�L�(����o���#��l��:��ng�=N��)L�CB�}�m�xP����ڈ'�	��2�\�98a���ӗl�l���gm駺���I}��Ho�~)����l6d�Bw�}�>mC�k4)y��cd��w�-�k�����t����&��$�7�V:^����_�w�ϯ�[�o�Mx��d!	���mi4�h��n�U���H�n�\�3�D��Jw�����4H�;�Ʉ��R�_}<W�M�h���(%Z1Ѫ����%�0Ѧ�s!~����'��{�фF= ~��h�XQ�g2p����q����i��p}~�[�������9�_�2)R�y'[ԃ���jd�{��7��.#�+�M���ĆB�0!N}���F�C��Ԃɲ��U0Mv\-�G�w������[p��B�Z"��|��h�Q��Z���l+޻���r|���/��׶:WD�ɴØg��ht�O��lQΕ��@R�QQ���#�?��Bb_g�x�O��0��kEb|a��l1��͙��Tz^i�ܡ��,����WYvG�g��Zj�����"��r�R�Ht�gY�k!�&>�w��+�)t4��F�D;�BG
���y��n��݈cG;\Z�Z	��Q�����ˮl_�\W�6�v)p+
�V�
�ί�=t��e����Y����N��@s�rAN��"�'��O檎��JύR #8*=c��J�c����q.T�MА/4��ۥ r�G�Uza��J���D���˞��ߣ����E�R�]�Kȃ�'�o=��kW\����y��DE�(�@iI���m�&;��Υ0�eTqa*�d��7������Op�5��0�WuA!)���#
��BUr��==�W�|�S��:�"�3e䍊��:[��Z�zB��{�\n�l���Z���;wu����<|+;���7�Ob8�"�t�B��ch(&=��bHD6T��6���Z�a*�xw�����w��k��+op�U_�[~��g'�2Y�\�>Y�,�[����x��l����9�
�/�r�U5��������co>�c��$`7�y�7�f�.t�oCy_�p�~�D�rV�CN �Χ;)�<�,�HGeJ��/̖�QH6R8�%l����0���W���'
$_�
��Bs~��p_3x#�ى��|�(�^�@�h��z	� �}@�0�O�����ԟp�"�Q
��&D+r��[�q�s��l��^���
��>��-����a�-Y��=�鲻���XV��/s���2�Sڥ ��f�P���N�B^���?`�<~��.��A6}�_/�e
g��R�0�
߭�@Ja�����ĺ�EP��>H�ge>1�#x��%N��ؑ�:�	D9W�8#Y|�
1y�9��h�Y�a�PT�{���.��_G�C�y;p�]�%IO,�k�0�Jl{��e`n�A�ܚҎU���[��%2�{)�4q�YJ�/vݲ�bRHo!ݝ}�+=c��D��z�U�*d1�x�b��V�&�~����Z7�w(���y�rJ��a���1��m��RxC����Nz�O&�۾��GT��'����"��D�aj^�Z�縺'���$�Z�pK�Wm�`\�ځ‛X[�9Þ[(��*	���)����[�����{
>ε��!�S��-�!�H���F7�jK�~-��]����1�����%�KR^��s3	3_��4���YZAB�����¶Z�v��¾�A���u�����Q}`MjV�v!�糆|��G�I���k��l�.1��;s0�b�g��AJà�6u�Y�l�6��R��ݭ�^�Ţ�)>���L����pv�Y��0�b�f�`^܋��/7���a��-h&������ rչX~��G�SA�䖍f Kx�I�����uaѵ��4�c���A�&�\ �:7���CVyU
d���hk45����9L�����fn��1�U+K҃��A6
jq�T}��j0�-����#�4R���L�b>q�ّ��~PuH��Vm���ۡ�x����8x2M2K�����?[�����ޤ��x����K���INw�f<P�����:�V)p�D���P��kP��a ny�g�A�i�S8��r�<,Ƭ�@���f�Y�S5Ԫ���/����T6�<�_��(�A���ة����#h��E6a���W�Rw���t���񐳙���,`M�NT�y�_�糃4hwO�MB8�4�`����>Nd��$Ad�pm6!��7���n��M6%;��Ι��`�4}�}9�g��L��-��LTwi�|�SO���&��`֞���})��A��),Li���PFz�{�lU��es�d��ͤvW��wo�G��"欖w�z�@
|�sY��K��\�D���4�g{��Y-��>��*�݋i!�@Us�!6C�:#<{Ó�q+*nv����a6H�"���r���f��Go�0�<ޫ?��4��ǁQ�r�镤/M���p�\�5�߷�[��L8u	���<|�r�83���������;�xL��Zx��
�Z(r�3��>ݞ��V��l��!����ݥ6F-u�o���7���	�\~1zq�!4fK����k��`��U�	�s�C�ظ~g	+���-���]��?8��`]l^��;�a�'/#��'���	۪���z\S>!/�#��ð+IR�bwd�p�r�!겥OKf)PP�QK�d��1�Ofl���(�u��1�4Ѵɤ���H⑈(<:�f����X)���Lg/KtF��8�
�Pvu0��g!�4��{��Y���̱P��o��e�(��J�B��B󑞝WV@H&��n�#[2��B��34��U�-I�nJ��M�\��~%��|&��-i&���N��@1A�s�";�hH�LH�F;I1��W�d8	+A/H/�q:�ymǓ��Z�M���;�G��������t��S$�9Ũ�d��܈Vv$~FK&Wu:~�R)Y�l���t�s�l���S�ݕ�4�Y��}��ɖ�#��1���h�]��2���^D��g"�I��A��Io�*/�F�������L�G�Q݊�{*֏Hu{M7Q�ת���-%�9�!����������)a���,�29[�/�,�l�9����
�v ��;"yF~�����ó�R񘪧p��0��ŏ(�$�	O%�P�(͂��t;��b�އi�$�'\E�(��1�!!���#���x���<�(Y��R�!<9j�I�n�`��F�$����+��q���l�MĞ���,��[�p������-n�����ul�5�.(���L�=����q:�h"z^���/@�u8��:���J�����i��Ǆ؊�Rk�>4���,Q{W�,��~� ^���e����ٻYv�:�Y���X�Vj����n���� Φ��N9'�C��Wo�Jʅ�5~N՗�r�Է��y�)��0��5xB�1��HIO*�Xd2��M�\�&T*�I.)�B_�� �>)/<�l�oGG�_���������x�;'���dVVl����=����`"��1��u��I�����ݨ�(��	�b!2hK��B.?=��OW^�����OOi\�2�S�1�l����r���b�)83=�L5�G�w�g2���%�G�	��!��0�z�DMl8� ks��c�dc���u�r���,Y`4D����UЦ�~����p~����lk����:n�x��Rdv�ԦVҞ��F-0;&��!�ս��ԉ�����`.� ���wbF���W���^����n����<��^��8t��.�K>H��G{/�woyA4�p�w��x�4ܹT;����}�C�'��u��|%V,���?�%�>>_���~z��rX�2���b�#��@�}:�y-����fp_����g>�[o��&ö�|�I,����?���'���oc�w�2�\���^���_w�3��9qp&H�
m��� �*�P�U���>-<+��h��q{h�ꞏ�Qb�mP��{�!���i��O���֍�?'�>[���啵�e��;�]��R�/�0uT�_n<*��O=���D��~��{�Y�b3
�ȥ�_��K_���fo�bd�Rct>������I�=ڏ6�i���m����
�\�O?����~�_`Ms�;�k.nߪ=�jj���[���Sޏ��[��bS�Q�_�4� ¿�؈8��p������o�6Mtb`C�%��nE#�q�qh�x\.GL��nIz(�z?>�o��H��fB��v�P��@Tv���sJ���@1�=�GzƩ�5���L�~^�3Jt��y�����0����P�l ��{�r���������Q��� ��b��HC}��v�?d�������l�F��	���h�%��C�7��F>� ~�-��	��r�4~.�&�l����"ꞔ*JA��+ÅV���X�v`PP`�7��Ц�\N����#�8X`c���!����w?�q�:$ixDN�D�痽�f
��f9ƻG��}8{����Xl˛o��A����,��S��֬��襀f������űj��������/Vy�|����plv�'	P�q�Ɋ��l�XdT|����Ǖ?-zʓ�����:�cg��qU�q���Ґ�Xq�N�����`�}"��B6á��-�MZ���ء;ʍ������x&���<~>�m	���9��:���dfs+���U��K�a7�?*7��D���ѕ��s4�U5�f��Sw�f6�<~�����h�����,{�c6ǪmÐ�sl@���� Q�r�A�n�88� 
�~���a%�Wm�f��G\��,O}6���2�>�&p<_vؗ��٘/'�����̗���w�Z�t:�P�b�����@��U�
A�ڕ<�Y��}<����Q����"|��	��_���zT������Nã�7=�#� A��W9�W���S������m<����G�g��_#5�'�W0�����Z�E�
ǯ��K����mb�^���ڇt6-��d���c����O��o<�3ц�F��.��7�f=^�U���
D�\n��$8M�E ��`Du��H�3]m3N�k?���Mݥ��������nc>6ͯ�E�����8��"�u�g(3͋��m�~?��~8޷��������_�(��s�W���X�	[���<�~��)V�Ɇ�M�5���13�
��a�U�����쿰�e0dK]�)ܭE��jU"B�٤U#�4���+T�*go�\��������BJ��`��ڙ��X��{�v14��@j3]�d�TB��<�����m��h.�>�5������o4ܲL<r��,���R[��F�cԲ�c�e�(R�τ��ƪE���H�K�d�����%��㟵���J���0ӂ%F�jd0���pA�����|�3Ғ`Oe��TԮ�
��]��Ě$�k�1�OS����[IƏʆ�;PT#nE(���)���R`%�����բI
|��4�)R�0r/�K�1*c��b)�e"4�\��x��~-��HA�J�kR? A������d݁�5�>	<ny���4�'%^O"Yg�lڠ��
��k�3�fI��dB�j�#a�D�t�W�J�goW]�#�_�*��'�4��T�%0-��-�:�K�7���.�#p [�uwC/��cJ���=*�V��ad���x&6�O#���b�vI��?�f��`�Db���4ȹj4�%�c��1Z"�$Z
 �Wz�a��b����p���	=��u�v�f��Gc->� M:�����\������?��������^�}xa46�te�JEt���qp;=�Y*{�O�������A�ٍX]���
ғkl�V�/�߅��T�#|G��rg�д
pA4���x-8A���V�fcz��7�W��> �yknN(q`yj8�XPu�(��GJ���I)���Ev�l���"�~�]�� K�7��D�a�åm�n�t��a64ć�<;��햇(��ߔ9�/��G@Z�����7�\��h2NQ�6@���j�z�%�z�o��?;�����<5�9fJ��J��u#+�s+5�S�(<�:�x��͓���ܙ&�"E׆������?�����ka�E0H���&:�'Z�߿�Ą��{S����K`��iK����d~��/������Y�3q+�b��!]��h��7�ҩ��w�\�C���s�]W-�+͢v��|�?����o����������l�p|����2�kne�)N�k���C�Vwn�
{����P6�d�I�4u�gou��FA�����8v�#w�l?��!���sA*^�7�	K���M�<`��0
��
.��s�ә+M��:<�[�+?���3�[�J�gs+��N��C���Q^��^�������T��{qh`>Io1�E�ڐ�E\2@�]�,�ߡ}:OoD�-{�_��C����`��`��^;$����~^r�)'�`�]�T����chQQ��=�)��P�Gܬ|}�s�c<�&��'�jA�+|��4Sg�k4��<���s��q��e��Ѱ�f���'@d�O�
!5L�dJ�����������c{���q��k�n�P���ڳen�={�\{�$m�p�����ܮ=���y3%�&0�;�����O#@[�2��Qa�Q/�8����ͬ�tz���.���_Pj��<�ʩ�T|��SK��ݹ�}	�����i/3��3U_G6��������u���Ε�aq�G��JQzL���{���7�ة���U��!O��7�v�7E.�h�3�ܚ�i�bc��.�������L�p�S���D1�~�.��b�O,DH[D� 6�<��*�<��̞D%�T��2
��4gz���B�������@�v�1�ë.�U��W�Y�tjM�[��:+k
N�#��a�h}���/F�0��o��E�I�,ҶE�W�e�������D���D&���h��Di�謵k�, �����$��Lڶ��D��cB��ԙn�-OՔoDmdS�����2f�[`H�����:���fPZ�j(4���ɋYB yta+˅�]-��+����.��ٜZ��N$2~N(NVg���%����T�+W��骱1�{�_Qx�
���vq�3�$��wLM�4<����Ӈ��j��V�I ��=09?8y];�[-���'/��9����%Q#C�dr�^�)II�9n0��֨7D�3!y���O*���2dI�Y��S.��D�ĈU��ע3M�`����`���.�a9�	�]�MA��俐�ԛ��(�o�E �\�������<��S=,x��j�P;�9z���r��¨�+"[��0�f��>�ׇ���r���J���n�ut�6:9�XF.��s���X��8��Ho5	hU3�ƒ��^t��(~�V�`R�[a����<�4��`��[��V���gF��C�,�I�N��
�>�>�j�h�?q���{HԮ��Ò��P�}�i����\��.�WV�B���PEb]��}�w�Ғ�F�Q���gEC1o�pJ��H>q�M��#=i��;󇳇J\����Q9�2��$����m��Z���\X�iWB�C�zwk�gɪV�����#�H�B�|u���@O~-�|�k�2�5&�ԩ4d�>�Āx�3	�N�)E���"9�c�tO��^OaxFX`b�rs���6�ӊ�͑��.��Vڑ�|��`_w��r�6ɇ���Εy���I0x���-j����p���n�V�Nr���0ߝ�+�<߮ؾy����4�M��������F�v4)+�\�ZnF�r�kU˭����!x�~�y��J����E�\�'b�H����V���9{�l5��.����y�.rH�M�Rh!��0Çpû��ciSY�Z0�u�����Q�C�`<���_��C]+�
V���a�j����k���3��:�~6�S% ��x�%�'s�6��3�_�u��0rit#R���?�#�Gs�����㋷ D��c �=��|yMU��uK�����[��p���Q-=
x�a_�/�����&���^]���M:��0���G3�Q�46i�q�׭�G�A6�a��7��!\{g��9���-xR¹�ѧ�� @U\{�n�~д�/ E�Y86�}�\+���O�ؼ\����q~�S��1Mhv�O��.�R�	9~r��R�T���L��fܼv
ˆ�$.���W�ϩh�'�S�v^��󻑃j8i�.���B�_P^=$��r�Iɏ�y#(Dl?UpPݩ�靁S��#��i�Y��i�F���%i��'CO�k��,ϒ�o/rI�h�x���5a�D��~�H�=�������^�j9R���X3�?�m(7�G��i۽#Pn�6��|��%��a ���pm��J��8�|V�������k��6�Y����� 3�΍�B�*��F�q̃q�Z��S��}P�����4�N�A������L���D�������a��ݾkE)8�t�d}�>lF&zA!,0�O�Rݓ�M�H�4��4��J�&�P���
.G �S��t�H�c͛l���6��ޗ�C�k���;���������Y�xw4��Q�z�9�gb]��q��!\��s�B��s��L՗ɦ�H��&鐙�˸�	�E��������^)��������"�P���$��ډ\{�[M�]V
��G!՗SI�+��Q�|�ϊ+�"kt{|���K���:&���G���Y��;[%��EQ��N��*�V��v���;����8���7��NDk��vw�~�0�s�Q]R[=�r���U�XEMA���F_�Mw����P��L���o�Ҏ��Y`�a���p3AU�=G[�&Y��Q;��l�Mi��Y�L��b�{��7�8��CYkV����~~|1�	�G�	��d���T�	�ƻ�7�@j����u%�d����XF�sT #P�̸<dI�#����!+%#7����zѩ�Z���bm�#i������6�����o�-�Fw��4)��R���~�T9g�k��Hg��*_:oB��9�g9�Op�?f���'���&=�AB�H˟��Z	L�	�8�-rK��l�����5G��Fn��	M��+䥀��~�:�_#R��+�9�X��w��&[�h˒C���$��	�S��7�׻�b��B��^�s]�[�h�Կ�;�̆�c؜��M�!y�0~�TO��ꦻ����.���f����_�?I���6���I�c2]���h��&[P5
hwcr{�Ԝ���z,�K�g��o���i��XJ�&�����Z�"4�<���Hh�4�����I�y�����cgS�lЕ�_�N��=jV�=��i�^��J.CB�whY�ɭ�oq��~n>�8��s1y��6� %T�����7D8\�]����J:��������Ϧ�C��|��m������m/����]��j0]���yt}�X
6���X
�m�>�+��lD��!�ef�~b�G��1���N�BM^��/�hW݆u�V�ω�`�?���+�`[.���oET����Fُ�eO�<�+r?��G��NZiƱ@�c�/Ϥ4���/o�~r�AGL��c~+�#l��`�]��\�~�m��=H��S�_^���퇥�E�-�<A9)O��q� 4� � �o��}�����#w!$��*Z�<d��PZ7W��G�i�-�.�7����j'+�e5b���<�|�l�ໝ�\�8B/���|�j�}`�7��3q��H�\�\�T;��>~l1��;.����<�|fC{z�M���%B��~H���v����ذ70���1yf����p_��պ	!���f�^��/��Rq�M�Y-��/=��0Hϐ���yb�6�l�@w��kY��2�F�N�es��/�S3��ӛ�i�B��D��I,�̆D9d$��f��� iOA��K~H��{	_[��hi:�O��,=~5�mjWp�S# ʣq�<�+��xǦ���.�dK�ȟ�S3��6��\��9lj��%�B΅+��<>(��G�:��\�,����۠Щ��*�3Ւ�],Y��R���b�҅���p��A��:�#���,��TO+͙D��=�5� U&��>#���&?�6�F��ܲ�G�!��B��-��=�}��<؋6{t�j��!Si�A���@z_=��Ȣ��<>a��>�1`~3[g��'.��PoV�	�C��e�u��[}�4�kh^j�����~['&ˮ����7C��Y���ģ�=�'J�J�4)�y
�Q�P�=�#������N�i��e�P���!��B������"�-�%���>e"[�}��dG^r�E[{�{\ah:6�Xi@���9�o����F�DX�U_�Xޒ�yBX�u{�Y����p�e56�M~�u�O��U�;�ʷ��r�{����=��^6���N�k�I��66�I&f����d"ā� �M��f8�S���Y�=�ߏ��x��ȿiA�S�Խ}�'���l��w6B�7�8�M��/3G���$�1"�ΰ���ލ�#�:ٔ������P�c�,!��+��{�g�~�j�ק=8T��˕����ց0-�f�e���~�<�'=��is�1Y-WQy�xaN�o_	�T����.Vj^�X̃���ہ�v�-��֡dNݧ6af$8Ps�����9"@EC��q7��'��/��4��\���N��G��[�0|
�s�pT�L�rwI��%�@5��;���<�h������J���:��R;1�6����hW�e�R�jg�D����A�M𵬊,�����~�c�t�F�	�:��ץ%���D:�� �A���"m4<<��}PǛ@{�B��=ԥN�'��&�^��!�l�2�Oa	^��Vw�У���=.���)�|D�j���J��\B�f�]]�g�=�(��)��{Oqۿ���rEW�z�W��dh� ��#�]XZeߒ=y�.6�k���((��'l�R(`�u&�(����~p����+K]0�
�V����0_�1����s�Z�Ǵf�Y�Y����qk6�0`��D7�׃)���T�����|�%���(�k� Qړ}���k�:;�[�1�,V�G�hc���A��3lj�Ba��=�,�:͢��k���@W��.rY��}�(g8��8g��W�i������%W_J��q_��;g�R~.z� �&�@�<(�F*���d��ap°y��zmp#�7�D���·�+#bۃ���"[���"/�QX��-���Y�C
����_edP�?ɗ��|6`�'�#0�-��K0�s���vt���9����i^��Ms��Y�26�#��� ��}�wI������?�Q!cp5����Ҫ��u7)�N�N�7E�(��U��7+�W�7*�k�L��['�p}���>�׏
9I�hځ{�[)���#ǖ�����0!ge]n��"��hF���ȷ����6;����P�f�rN2������m�.��w]N���ˊ?���s攦�)���{���SC������85f��n��ziEY�eV���%1�x^����
����獶�����Cq��0ן��4
H�E0���w�$F~By'�#���PƸ`X �UI�"��ݤ�o��:��_T	=߰~;6H�o0�m�aER�}��`;���J��2>��˓��*�*GS�?4tEP�^�"��8��oĺ��O���\�Z�hT��<�I%iqKI�LD��
�j�Q)ƭ�KE��m,�A�~�e�+�/�f��f9�i�n�������E��buow6o���V��9���k�al�:㟼fVA�p���z��*
~"&����j��[�xn�1�����a����H��ǆ�
�Ti1놢�~�4
��������1&L�Cȟ����/1뢇��}���[�+��Jo��|�A��B3�	�!�U���忂oA[p⩅h����i��S,��"yM�t���u1[f��,D�}4���Vf5����E�A.c�����u�#��)Y�\:����VJ�C9���Py��bWY=��R�nb�Ū\x�%�l΃�2ȖY�k�h'\���L���*����h�"Wqh�j�]j���A-~V���e��E>/R
��&�!�JE��<q/��`��or7
�'�4�"!^Q�7�B�xxB��x�[�4�K�t>_�.B���E��@�<��6}��Q Hl+���c�fw�v�*���X��I�4\�Z�x4�ݮʹq��(3�JOX��T��"S";�52[;�$�ab԰6�J�Z�:�	2��q���t�H\q	�NPi˯��A
�A���ql9������LP���2���:	���0c�E�ut낋�'yj��'�V�X�<O��@�\^ڭf��'�q�<� �ɻi��^>'�+��jǼ�R'7��G�.���7&��ȟ�K��P��*m4������@��ep��S���i��4z�����0��OHnAZ��>ň��[��Z?z�;0�&4��?��b�b���Q3��K�	++C�je:X^YsK~�Lo�`��9�����S	��P�5�J�q�V�m��꺤�a�{V��<�}�
8���(���y���]�
}��5�
jO�k�
J}�R�R�4E��A��~M���p�".��)Y�_3�m����.�RQ�Ȥ���M��)�B��(#�.HˑQ ׯyyKېX����V@�Ũp�ʨl�TdT�Zjf\`ZjaT�Z
y���ƨ`*��҅�_�#y�a��_��E�k;y�9L��N#|	4����b�K�O,5>q����U~�:��X��� /���*��hN�ќ�L�.��S���F�]Pjt�L�ʍ.�0�`!��� ]8���w�;y���l���U
�	�p,�۲�h�2�-�і�F[����m	m����2��(��.2Y��t��2^��hӻ���k���x��N��*��H���g�=�?z���[j��2c�dc�V�We�^-=�Z�Ja7ЅK�V��L�Z͠�����K����4wwE�<ϽN^�||1�O�k�3�c��N� ͮ������y�w<p�P��&�Q|��d��C�w�ޭM^��)�#q����4!O�m8儾��(%w���SFzL
샽HI����҉�����W7��'�����!��\�=V7 �mE/a�&^�+�W�s�Q\�F��mt�ž��#M��mG����M�D��F�\���,�!����?��Ń+�ҳ�k��)�N��ک_m�X����߁2&��s,�F\����3�O�H~Y��6IT�Q���<u�woJ:o�%<o�x�;A�<��V!_r<�kXAJo�ɛ��+�z^3=z�N��T�8�uq!_��Hƫ��=��3��q��*fV}/�UB����+W���ށu1v8��x��g��~���!-�is���o�╏/~�J���wo���)�>�P�#va�[дNI̫u�F��|�9]�u��k����s���-�덴�Cږ��o_�[�ڲҴ'�v���@N�[�כ@�}�d#���qbK�kH,��"�Dt\�8���_#����e>INr�Ч��4��6u��D��}m;���ȩ�3����p��p?��:}N��.�/�c8���FE�5帠��ԼP������k���+�՘<�eGDy5�k���)_���;�F�'�y=D���1�iV
���2�Q�k8�R �CÝ�_���p�q�ޭ����� HG��3���.��Z�aG+������VX{���'�J�����Wee%�#�r�g4���q��؛��3&�:
fy0�f`�R_JAt�D�.�`o�ֿ�T7H�i��%�j�������$`Ӳc��7�mٰY�����u�,o���B�DD��ʉ�z|�9H]��h�L����2����|^S��q�o|7��y�|[p#��%\�|��-Y���+6��9cc1/+	�:��B����S�)Gm�%� �G"S�-<�ИcNgjγ� AB�k��$y&���-+��Vl.�˩��]&�ģ�ӡ��E[�7�Jg��_д��u+~Xt��_d'I�es��if�����0~�D:�1\�K�8Q��������H����Ll�Ə��X�3DDH"T�&�:QK��̌�<^5+$pT���jj�,)T49�p?vd��.qb�j����#�V�ڱI�V(J�S����n���_86#W�1�����މ�ݿ��s���ك ����$��mo+�(�;��r�ک� h�X��I�/��vHG��8v�w\�q=�x;�Y���]�-4A��,����pr�St�%�����ol����$CJ`D���-X����تiJ�
�VD�Ȯl�,V�����:�vvv�Ǻ��u_���wWt����b-*�RA�u��R
4�sΝ�i)����:��s�>�=��s����jb+�O�ŋpȅ��;�������*�,���ƫqB��WyG�!��;��n·AG!��u"��%IX�"�kum_9��p�z���j�a�U�2����k��L��o�G+G�P?���r����E;��~�st�P3��`�K���Y/�A����)��.�OV���.�[i�a)º��	E���Q�T�L`_�X.��X�=�1w���P8K�D �����{F[����r8gg�m�T���W�o��G��OA������#Q����[|���3hn��A�A"	ϙ%E��+<� ��նr�U�j��+<��o�����Kb���j��,{�J�8�V:������DNO��#ϴêܪ|�d���T�o�<ӤEtӰ�|>x��G{;	|q�T�aM��s������V�.�ӆ�U��Ҥ�G/,�"V���[�ٮ9�i^�к?��PC��5HZh�L����=�
�c@�)G�F�or���	���<������x�ӥm0��9y�����R�.��ٱ4U����r���<<iS�J�A7Ǽ�*��LN��,4��ܑv/皛�z�������%��3�)�h���"/5�Q]�+o���(`U8l��ֽ��.�C6(���}}P�G�|V��q�������y�s=kϬ��x*��mOG}G_�򸻫�}�0܇��иM�����2]=iz�.R�c�5,C-�j�-Jf�jh����21�7E��9�Ȣ����͉F��?���y�)��5��C������{/��Қ�?rb�1���يމ���c<�u���J����/,n�Z2��@�ۥ�
2nH��(�(Y�qb!Fk�Os���o�of���_^�6h�3�P>�0Í�{�n�W�����7�}�ҥcu�_��:1߰6UW������m�DSmT����uw��Iu��9B/��.;]�'p{1p����fr�,�'t|����mC��	]W�?/3b�3��7���os���E6�ϯ���c���=��m�DG938A�������(���7�����<ؗ��M�I)�{�E���$��V=h��G�C۳�	�um=�n���8_>��=�Ud���"�,�+�� ���d`�S3�G�$����sČ��_|��p̿Z?��1wc[�Ww#Z����{k���S�Ō�E�cߠ��r�� �ϣ,��_���CQ�=�@=�n���d�_"u��u���5�#���G�3�K��t|�/�u�܂��JS��Q�70h��\u^
ۑ�('��<��h�Z3�m��"`��3��?2�mx~;}�S.��Z�H͕��m�^���B�p�>�A���g�Y�cɮp �ɥU��:}���ߜ��Q|���:�_aVc{鏆���`�X9bis)��ȥ5,�7�K�`���]�V~SZ��N���� ��[tz\��q�Y�z�>��$���!}y�j
��h����r�bg�&��B�cܔX�7�XF����d�*Q<J����hp�&���?�����#�(�}��:�ᄂ^5@>�7jj8���k7_����� �ۢ<}�U#�Y�qBf�7E��\���6�ZjO�7����.e�����W,�く�0p���ۆ��Ѱ�W�1,��	���������ب82麷_V���-8���	\�7���gȹ�)�}�����<����{y��>\5q%�(�G5!`�-�q�=�_j��)M*��sR3�1*xpԈ|6�|Gڎ'y��!��ځk���\��D4��i���>�7�N�\K����G�P"K�Q�ĳ:�s�&��������qI����G��wPD
H�b����S'ۥ��]���;����ͤ���*Kz�1o��Jt>�FoO��P�x�2�4�)�|ZQ,n�����:Q��Ⓦ1G�pT1�&țC��?y������\�\���T��摿����)�-�'��p��C�B=�)U8A�VLj[��i���&��S1$�n檅v�=m��M�����������4�dfp '���4:b��w��g�e�s�%-���DY�c|��X�5�s��3xy��/��s��M�]F��*�s �	�!.��%����G�F��vXي9+��q.{D���L n���jE��A�xRD��0m(�̩|omb����7Uε#���}h�U"�Zc7�,���k�=�m�A�Y���5���9�Y�jVǊ�:,����Z~8y��8�s7��� �b�\�4D�i���ݿ$V5s!��-g5�.���,�?<��w}���4^$�]����؛�"Y����!����m�?:�1��s���w�;��8B�����:O���X�Sg�)���;�T
��? ";��ο�t:�7�ö��C��"�ۃ�ڢ#���Z���S���EV��^��f#sm@6;������O]��N�>f2>�Oy�}�=1�|bزW�Z!{���x�oU�Czc1�J��%E�{����$F,ΐʍ�I�)\�)ZÖ��B��8o|�H��B:���K��^���a�dW�"�������ؚ��H\S��x������^��Oh��h���%�vS��K�N�2�+�<����TB�;�Y6&��.u���:|�1}]��W&���~ie?Əd�L`�Ir�v��("���D�q�)>9`��%��x��`{f�N]98C�ד1�&��1����HMB�_8*Cњ����ӹ�MO�&���@�H����I&�8a�1@݅C@�+65w�8 q�C�<-����(`�C��]%���M㑏��D��D/?5e�`�����Z%d��<����s��j��N}�O�J�>`N��y�ϧ����V825�/���"a/:�Oj��t�ge`	�@�"2�޿e�w������~k�?�����tO�p�?s���8f��,1}����~��,�j��c�H6��X~<z���<�;��i�����"���)̻p�����[%��P�+h5�J�z���pL���9%����0?n�P�6���	L�p}���Q��O���No�o� ?�?oy/ܟ�S�ϱ���3���?�/�����s��{/֟����}��~�d]�?Ş���|���}��~
F�~�J�n����'��n����νp����<i~~꒾;�ͺ�B�y�u��ti΅�c�h��<|�����t]�?o�ο���p�'.֟I����!���ȳ�L�5���e���������[���f��5����O��Ӫ!Y�Ҥx<�9�����糛���1_�?o����؃X�� {7�?y#�ߟ�ߝ���|!z����-������.Fo�����_�߽?����e����h�4ߟ=�w��#?�P�OM����q�b�i�ߟ������q�����ߟ����?���ӟ[t���M�7���i�-�����ÝG���w������?�_�?��\T�ѝG��O��p�E�>�/�.�[t��;�V�B�|����?U.4��&����h4�V����1�IG4{c���c(H7�r�n���&��_ ?��϶)�8?{��\߱?5�j�.��R���ҡ�폍�j�l8�[lם�CP�����X���>��NP�T���Z>Q����h�H],�Uj
?�@HK�(������H���y���A�p��!��FyY=g�F�;���3�|كA�a�Pi�A��S�����
O����fZ�ږL&�4M,]�K�u�X�03wR�f��1C�l�Z	�'N1Dr�l��L֍���+)�@�i�X�w8;��xt����$̞���@�R�oM�&ԧ#8�{�d�K���U5]���2�U]���y���!"O�������te�+����IqU��������>	#�z]΍(K&��<�}n>�����:x\"����B��.ɬ�p�F�P�JXX|/�5���E"3���Z����cD=H {a����w��C��^J�n�8��'�#�9��A<�z	��-I8�	�οW�䷟�?��X�������ɱA�㕚}1?�D�d��Hk+�`KewZ�b-��ҟZ"�>�?RХ#�F.����Q�,��4�w���R�1`��1�]I���H�2��\K4�4���F�����M��q�L�-����j��ـ�T;F	�7	���p���ŷ�`/� [������ʣÂ2ώ��S:�q�K	[��9|6'�5a��-�����5*��>Z6_����a0�M|��FN��4|�2��[՗�(��9���nNm؟�m{W���:��v.�C�5@\�~#�5�V��V��BS�3��E���wފ7��ej���vQu���j�z:��
;�7�O�u���gjF���3��D�hv�Ń�+�ڮחJ�Bm�c�̳�hT/HQV텁ȳ����܊m_1�A5���Z����������bC�z6W=]/���Z�:N�<YT�Xߊ��M}�t��«�i�<F��gH{�I,%,r9��5�v/O�%�\u!Wm������3�z�z;���3u�6S��OG��&�v��p��U���di�����F�V���҅����z�w�gbs�76r�Pk��>O�<��p5���Vm<_DO������Uu�0��u�u:_��Z^ua�|?Ã%�n���a�F�#GƉ�1�GR��ҎꫤHC$��H�x�^������8i{C�(4�G�z��z6�4�it���bJ�t (U��iG�a#ԪbM�$��_�K�&X���j5Dǅ����R~ (��!�����)��g	:�����_e��a���79G�������""����_�;c�7�SD6QI� �| ~� ��<�J��I1<����{H1˟B(%��Pf�C��C�j8L��%Q�<�=^}�ls@OT���AT�qD*�l��2c���RE4J{c�u=n�އ�+ŵ�,�]�K�� >&�c�a#��1�!<C��� o	��#���M"�Kw*eJG4ʂ�w+��gOj`e����ʫ=���|x}�)Ç���x����\��1ʹ&�c�#y����8�v������1ZB���y�Z4Řݚ{�Iy��0��kßw�p�&�g�(Oo����J�r��?�R�l>�O�09e�!�My����m�ߝ y�a�&��bx=�&�z�^y����dt�i�ߔ�bȮ�3��^Z5Ө�ke��W�Oȼ	�^����b�;�#x����ߟ�;�m^%�X������U��ub'֛]��j���U���kW���Ƙ���o���Y��4�E���_����SX��F�E������ItIu5|�s[%�T�W��W*4��5�Z�$ֺs�������ye�E��V�+{��ݾ��yKq�Z��H����I�k�]8o�ܥ膔�F�ᅼ��M����(f!�v0�����X�%T���l��?��M�|�R�#��r�ߧ�>��}����<�o8�KE��m�9�'�+��.��"K��;>��b�{�4��G��c�a�I����n�N��[�D�F���ƴ&����S[�z!�O2�/�_����O�/�9[�8�=Ѹ^,��<#�>b��A�F�i��򌾔�װ��_��j���I=�l�ks�e\��<xP�R�#���>P�٭|�O=H���R.�F��S��؟��
⧋�\��W4�����saZ#p:\���(���f|ګ��G�� �����A�P���?x��/�;|����V�i�3\�,߃��w��*}��/�M)|XP���^T���~�c4ON�n��ryy��֒Р^�k@��P(�c�с\�,�&=:Lx h@��[#kb��i�z�y�Q�j�>[]�Jy݈��;y�F��*飺Ku	Eā0!��0廕���7X����^̵K��ſ:]]PcN��E"Czov_�E~=t~X>�������R�Z}J[fQ9�K��'���O��<]R�r���a]p4]h�1��Q��8�ڇ���MwM�SAh~�*�R�@��w���T|bb<��rb����V���K�C�N���D`�-��5�NT8�7�K
ds9�#�L	���r8��s�'mCW����k�b�`�f�<�g�!Д��^]8�D�14�nUF�k<����uȄ�,_�`����[[��0���-<������EY��P�ё�`N�&��d���a����p���)��;*����R���R�]���Q4��IG�K}$���;�SR��66L<jy��`P�u�����w4^Ij��L�z��o�k�����ʇ��/q�|�\dG:o����걻Z�%�M�$�/�r�&=эWʝ��=���.���/~���2K��k�V�n�l�	��Z���TڬX�[�t*��zh\�ڑ��K�\�_[� J|{1��Q��@̾���nK���g��8��͜k�e�a;4o֮� i��@e0Y7����#�������2EbYBc�]͏N`�c9�˛jq�#��OՌ�F��}Z0�.t���J�U���<9}�C����D�o»b��ZX,��	F�$B�<aW��PDeGCc���$���]�	����5�M�dq�,l�X��g��/b����G�I����r��������ɘ�k�z��n��f�_=��4"���Z+�������}I�2���. ��'Ϋ3���J���?�����I�i�&"-D���:NK&�7�>��9ҷ��5=���m���iw���`��õ���e�R�§��AXM�]�g��F���Rq�{Bfさ3L�A�_��=�NJH�`L�j��8��C�MB��Z�*!�6���_�#t��t1��������SOhQ]8�1��(9J��/��j�[�T�4L|9���wu+GR�ܒ�ܫ	/�:�����dBO��f�?~}ߠ'�ٓ�%Yu���ȷ��0S{�3�~��*k ��Wp���9y������"U��:��r��W�_6Q��Ct~$�1��,�r�,ǆ��,��k����x�枊7����,!�@�f|��Tm�r�4�D*�Ӥ^��O]�'&���}�H�elo#��E��Z�-uy:4WA�]�m4����o������ I)U�鶕��7�սq�=�G�x-�g�=�0�+��<`�ˑ�1�

<���p���q�����'3��|�QDnz���>{[҉�*���7�f~W��l�Vy��`�g��� 걅'��s}��u�>5U�m�g��TR^C���ax/�ξ�p*���"R�{�Q�	��LD����f���)�,S��:\�s�0.~X���yv̼�p� w�Qȕ<l��ܗ%���Q�<���Q�>�Id.<�>���]�P��+��K#�Ώ���3���LʳMi�tJ���C8�7dK��	ճA����[�;�c��#�	>��R|�����	�'۫1ˇR���[	�_`�a�����|�^�
�<d�io��Te���1kW`�d���E���g8�#X���<��ty�����p�x��<�Քꉌl=ӧ����{L��ozv�f܂9�F��W�[�,�p����c�]~�.�㨄��OD�;��A��@�X
�~�t޵�ɛk`3�-�=�48W>�?"��n��_�S��]�,#�j��t*���Ơ��� �z��³�^���� ��-&[z���'MC�VO��ў�v߻r�9�ꄷ��p(gַQvl�$�:ֺ��Jx�g�^���Yu�Y�����XC+��R��<�w5!m�B2�\M�Q��z�g��l��&R���e��yQQ�K�̓'Y���$�@$�_��	�n�do�f��˓gÖ��+�L��M�W�T���7��\�ѥ5Bm�M�~C���;,�V�,"r�ټ�)��/��#��Ǝ̜��Y7�2�Uf�eDF�~W��6�g�E�Q�qL.�N��¦V�B��i:��ӧ���Ӎ�K��R��?�~�<�KK��|B{�O������������n��
��g�1MR7��:�xO:n0h��~F$=�'B���>R�#��5:���-nx�?V�O����7���Po�W:�NW�d�B�3��2f�:�Ő��;J2�W7���w4�� �E�p[4`���-���$�߅z*1Հ��Y8#��}�:�G*7
3�2i��fK�Av�r�f�Bӕo2�u�������H(Zm6����՝�e@��rc�P�+��k�b1k��|M�;���w�Sy�zo4!��DYt�"��W��GY�X�Mx�"�q�Lw������c g�ۀA-�pZk×�pv*��P��D%�@we$�E.F�ÖV�Ӹb�����!읐����Z) �m��\�w%�.�b�7�#-�(I�����n|�h���ష�d��R?�����.��k%M)P��ì@�@�P
Oh8ģD<��/�>�AP��?H_�e�l&����`���e��gg
/S^�����e](�֟�5}fB<^@�H���VZ�}�O���=����+�����T6�Ì���[�QDP&�5�hd-��TK�3��9�WZ,:Vb��62�8�e�.<7:�����´���bQY���m�z2VxA���ђ�F���)}�R���)N�qãI��k�p�#�����E����ds��+r9����B�w_���%������ ��j'��*�K�<Ӗ5#]>�S�X��f���@{P��(�Noh���:D*�jg^#��f��k��i�= 9`Z
au	�c�֟:W#n��f�����$�q�GYZLQ��q�,��(=���W��{l����R��=�B���u�7	wУ¦���F�/PۚkJ����d->�3�Mi	)i:����_���GH��m��Mw�M[���\X'��}��6��$��1�%�B���'/���|)�,O���0(�{A��͐S�|L�����C�끳Y\��:���e�K͚k��GXW�Z�5���jQc�1��FYy����g¯M7�c�Gig�f�х��۪1�tO�� <4vV�Y��4=U���G��hWMm��5���J��X�Д@�;�/z�,/3j�PUI_ɜ.�=�""��i�Ã���,�ѡ���Û�<��=�/��d��yUc?+ْG#���E�~B�`�*�~K��#[�	��Lh�1���n�l��/�xE��"f�~�4$��G>�����a����fv��كv2\02ƴ WK	�DC[}�ɹ K !��ip2G�Y�7�<Վ]��Ů����0n��-�/�M,ĉǚ�"�ǚ{�-��Yᎅ�0���
�?��S2�i���������we"�E^��2���g+�5�ve˗�sd��Ǡԯ���w×zT�@	jg��5����VåH��(�I��ˆ=��!xk?Gb�YCf��z|�ބ��?A�]��Y_�r3�m�|OΥ��2Č���_0�V�#�O��*࿼��Z�ş�F�
%fzL�	������{a���s,�>e�e���N�*C�0F�#�
�Of��w��_�W'��!��i��n��z�#�
�:�c�����ï�,r�u�TZ���1�m�c!~�I���y�b�i�tͣM�dk�o�#����k)��LƆA���Mx��ei�.dVjhȇ#��h ���^̈́���uiGu�*K�D�E�	� @!q��K�#����T�~k��s��|D�QK�c����;H���o�G���E1���������P1��-Y�j�_��tð'&0���}��ى�h�lyIR�&N�|s�u�#F�Uynʗ�e�fboJU����7�9ñ���J�V���~:�9�Pb���P@�d���*{�gd`
:������1�&�N �:�|�V����oa�9;;n��$�T�R�g�m�e|'��\�wrߑ�v���`����yf^�cԝ/}"x{�<S�N� $�#&M
hL��P"r�e�8\���@4�cw2#����
[�C��!��LŰk&�T2�&��:��تŁ��#�W��V{T�1�u(�[&'Is�ʗ(��)�9�hT��لj�����
p�f;`>���*/�����4�G��z�-�G��.<5��`��I\&�(u1��(	�r���,m�q?�ھj��8�6��/�O�9O&��L:����O��{��쁦0�<�.�� {���2�3L�u���LM�tu���HsiM���X�����WN4�3JKYj"���,E��qJL�֌����&Ї��Se���|#���(B�:��vi���}�<���u	��9�kx�'�&���+����1���P<��	1���%��RJMY��T|l*�Y�Yd*Q�����-	m����،�Ҿ�r����a,?w�o$�n�������؈;ya���6l`����WA�&�n؊�fNy�����[��!&nb���	�k��{�Z�ɭ폂}S��$NK~D����)���A�@k���=��4�@����lx���WS��0r�D�����G��4�J_�
�t:<#Zy�<�(�\�M�B6��L��t�W���h{�H6"/��:�WN����xB��m���t�M�-��"셚�oT�5y��O6�p1>������A}5lXB�7�S<�^������%��k��;I:��'����FK���0��˞�5|��&�R�A,@A!؍�ۘ�a�V<�~]����?/���s�E:�T�_�3Om�oO�"B�a�a��tBh���u2���P�x�]��H�B��8�=�B�S��6��uF��2!�1������PyF�A$I��w��q���>�P�]����?�ǭ��/��,j� �1W8J��0�l��cj[��B1P#����6N#�~�Ҡ��!<凮s�.db.�������\d�ԏÉ��N��1����]��u�GĽ	>M����!؎n��mp��*����h�=P�aS.6���\��!Y���mqX2��!���u�κ�ǣ����)�fJ�A���F�R�|/6����&M��u���A/�N��(p,<�!~n��}X]��5����/6��F#����Ul2�E<H
h�����%r�o�1�{�`��kA�ѡ]&=��Gj�$d����@��!��I�ϙA#.���R5��`����O��o�^/�W7O�)�Z¬��Hݰ�ơ����*��<w��X��A?���� l�?b�jB��x<9�ya��c�+`7Ɍ��O�M<l����)>ogRX�Y���3BHEQkFeOp1� ����@&ԑ6�=��FRٗ�=���7*�c9[�+��B�"�[5O.Ā�&^k�dV1��ֲWH�ˀAJ¯a���Z�A��P���%�ѱ	�z�/<��l�qb1��-fq#�����k���CKjD����?յ_���`�:Z���]^������
�?k�~�WG�>�k��&!X-��ݵ;���H#��s���p ��}��l�Јz�,C� ��D�!�Wl�(��;e�{�����NJ�����V�H�_a.t^B�)@��Ѭ�Pkơ��h�O3��R���`(�ER��o�9����6`���ks��%�"��gq�q��N_�O��W�[����޼���1�Ќ���Qdw+p�C{[}���/�ZC��Q�0g=���g�]ݾk�-h����OK�2?�.��ο�T|����n
� ����/A�@����f�#��P_��\��/Hj���ݑl�_$D�&���]a�g���s��n��J���q;R�x�SO�q��5���Z��[��2�/�h���TO��7
�^�5��M7y�һꍧ�kg7l��`�����N�I~�XF���wd7i'�w+p_/T��.)�-~<�^���(���3wz)pK���g U�MK��=�I�,�a:Nw��sZ�3
����#��f��y�0G��,_)W
�&!���<W=���)r�$(�m#��]���>�î�͗��eNeGj�D�a���UM���4������pu���xu����?g,����'���=���F��Hհ4��z�Q �L���OFm*�E��%��Y���ʗg(D*&�HN ��
Bp#��'�*��KNƧ����\��\�@d8M�`��t���h
�}�d|��>1�#����$=������XA*ө�O�~�����"����8r�!Ti�ٿQ�J"ο��ZK2���a�ʠ=��o`s�^,>��q����өvuO���a�8�����c[�e���F";�Tutuv�vlc���E�U����ۄ��+�{� &��kwG���f������(�D�[]{`��"c��G�:�fw��V�o�����v��qw+�#<���j|k��#�k���-Q]�Xc�V�kh�W����r�@u���
Mܧ.��5vo�xĨ�<��(|Q�������cnZq�k7���'�a\:��N�
���
��������/�u/	Y�Jqit�&8�K��l�	v��뢳�m��!��t�5h�Њ���Ƚ�q�N���&��x�A�K�p4U+�J�h��i�c%�g�3/:,A���Qj�ŉY�� �s<F�=�k�S<��y���O������^�u��r�s�,����a�'�h�@w �$�)�S!C6 }�k�!l��z��]�|�^��s�ƀF�>E�{�c!Fi���:3�ׂ|Q���߀�ve&Lu�c9�+a]�c�;�R�C���Y�X
��g��ݥbCz�ױ�3uwkD�����t����(E�
�����R�/��0Z��eҶ�ۛ���P��	�y�]+Ğ�Fr����;��B���i_1������W=�������w�N[}�`�~�}|��00��f��mG��T><"��8��W�M,�j�v�߂��\k@@N'�T�� p�&5�ib}
����_�f\����8R}���$l�,���W�-�H+􉽆U�Ċ)��$J��$�9ϵ�o?���.vs#�|�p�H�o������H/�D1�~u��V����W�`��F�Ɛ���HPӤ{G�Ξ�[����B���g�.�I�ܮWw��Wj�M��D���ڶ���D���	���h�v��Q��ˬ�	ԵJ�G����^P��?9��~ާ��D�P���S)�`i������*<��_��]h^��"��&��t߱�B�7L/�f��@Ӂ(U�֐�NЎ]���k&�l_���5��L������}�vu �*�q*4��J�J���D}X=@}a� �Q�R���Ѫ�#$��Yx���qIs�t��l��i���˨R:�����LA�9'�G�uӑh��Hxv��(:܅�J���8��̣+�T�+�}�մ6u�17Aks@���Wm�DZ�pׁ�.�?Xi���
E�<$u7�^��7brc87���P�"�����ş��a�W\=>�ӫ=(��_�F<P�i��f=N����לF�+(+Y��n�*C�?Sq��~2Ӌ`���N�mzu�)&����|�Z��AX�Ђ�-��1����{\xd��¦�p�˜�G�5�MI�]M��Bx2�-�~C��1��n�	��t���?��Ԃo4�'�M=j�1�á4��S�������paT^� ��vq4v��E^t�7�?��m&�Tסtl#�����Q�}4�@J�n+�ê�
�oO�\q���
mM��5��呪dk�!R��:�B��z�-zU}M�K煽�+8����"��1�rT�T�����09:e�!:Q[�&#\���fOW�9H&�Ax�&r�) od�RA�v�����"v��8�ŎT�iB0�kRk��p�-x�en8`P^c��G�uJ-�W�(���q|���I=yr�c��-�N`���J��Q�v1C+���<+�K<�B6d�
��HI?,h4��59�r:�ZZ/�-hݺ��YJ�7��R�;0h�"}G �T���S�>�.���EBm��I�O`o�jo�n��������kN��yx����
ÜF'z�yE���k���AڈN q�8ߑݘ�"����D��e!xw��+`&ӠQ�G�~�V9�I���1%g-M��Y���<`k��w�t��y���D)6Y+a�$�f�OI^�(IcpCtP��}m�f�?���ًUx��\�N>��6�4El����!�X%~�ڊ^��# A	��4XSxȅi8��Ѯ��m՗�"���Y��S{�)�Hx��ꤘ�-�b��!�z�|+s���6��W����2$RI��s���<h��u��h�����*ѱe�.?��08��ȝДP�/�5��e�?*#s�W(u&��	)��+�Mg�xn����$�\Y�x���y{.˨��´Qq�Q ���בrͳ�]n�=H&�pA�~Z�G�������b�-����m��7;۝�Y?7���qY��&�56�]��#2?V^�!�́��V ��t@���yZ����v��0���J� �?�rx��X�����'�H=��h� 2@��H�������G?Z�^O3�ʞ�b��`�l"�5O��(s�e}�4
��
��L�Z��Y��2��;u�y�x;�C/p-�A����%Ff�+�(���y�*���p�k`��(���R6�����,}�(V�W�&}�7����?Y��	���%�{oi�!&F6s�o���"��2�3�ൈXM�_�({b����l�8������,g�������$nB�ؐ��O*��gR���Q��2���Q��Ը�;����E+G4{���5��p��\>��^�Ž2���705��b����(�H7�I=w*� ��K������V����O�äcW�����l�Uhy��t{GE�Ɲx��N���K���J�r��4��ù�q�l|qܐ�&����`�1ޓ�W`D��ݭ��1҃n�~ā7V�u�$b�)��
�|�y���s����v�Ƶn}�Zt�K�Z�t {��K���uT�#�Y��.� �(5��Ť	6�<6��$��8�qǽx�%��T�_�;'d��bA�RV�����-p%�"��
�1����+[Ra9��[,���?�[r��/���iiA*_N�C��'�Z��"rLSB�
(d�j7<�������<��Z�!�6����ϳn��({m�1�p�Ϙ���7�(�8b�Ю�MK�,����arQX���%(��]K�}��t�4rh͂;ɸb��/ {�����Vri�	_�=)�ɋ�p�':y���=�����AD�k�L}|)0���D�Qz-ޡN��Gy���1"��kO����+��_��6EKL�cq�*��9D�ʃO��?�~�6-���P&s��]�M�'�#7Ǘ��a��4(u�S$ƻ�=T|.I�����KU'�k�_|�?zn"L�+`_��^*8A�)�q��y��e.E_�(��m���\��}w
�O�y�G�\ڦ�Ohގ7��Y|��|{���-�������+�;_|K[<�RN��b��<J:���a�Y7�?��"��Y�(±]�n}���U�H��_�|á%�~~��ro���_�٘�� x���t��\�1�E~�T�[�<0�1�4����#�������
�����F��m�ELDvl���07-�v9ӗ*϶8{B��W����L~s���n��gL����� L�r���^��ڸ��#��w�,�IĿ�-�V�pl�bs��&���8i+U;�m�\��Gb"�P�J7 ɐ�g��{�k��Wd�:���w�u+/���wYP
�f,c|U�0�Ui?F~�? #�M:�44h�0h������($���T�i@FĤf��SL'&o��œ�W�ɡ��w��lX�մ_�]B�������Rc�;~�OB̕��J��G����S���G�|�Z�5Xia���3zU�D��(SxuR��Z���nPĔ���C'/=A��Z<$]��RM��	������E�X`�ڱ��|44��<��=v\�T2�[Y�+j��|�&�߁�鄔��G���FD���g�|s䍨����eQ�4t殇z�W[KnZKO�9:��9�*����!(�M0�_c�\�2@���J�I�|dGO�RUO�ʭ�t(��Ց?����4��m���b?��� �ߠ��N�M��A���m0\vs��w8&��JM���~�G 2Rb�"ƻV���+��ņ�١V��B�����:r�_ �A��{bs�d$���$�g#%+�)��d�%��x��� �cS�tsS����U���yC"��q6�ߴ���s\tk�Bx�*�������i�Ô���Hu�ֳv�0��8�?��=���cL@�
��\V�>�-+ߥ�|#ҹ6>�����F[�F/���4� F�!�wʠ1S".�<C�SOnE�{�"�V��W�#tCX�I-���bJO[i�WzP�[�<e��y���h7J�a�<-�,-;������X�S�t$�����5���ʇ�<^�j�NXWd�i���ĭz�9r�Z#���6J�.�����o�W�C��im]-�gq7�w�ZW��Y��Q7��&�5��
�Z���n�y���/t�7��/s,,��8�W�C�hi
e���C�ݚ��#�ȹ���B�1�j��P�o*��@N 0�_Pϲ��*ǃ�+[���l]�ڌMԒ}�� ��\�On���Y�T�^1u _��&�O	I :�M9y	�Y�ʳVd�m�QU����=$�'KM@M���7:c'J,
��r�O��Zh�1���AS�o�݇���c�(��!}���3�}��Q 1%C��c?�p2л��~�
���͈���~;�c���x_-�ť�0�}uר�=DR�>�EC�g<ߙUS��'a\ϧ�D�D�����x	H}����W�}[��9 5����Ҵ��iF�smb>ϕJ���E���E�+I�t���#�P�	󒳵a�J.�v�)��f&�e��U��O��YF�@��q�dQ s�|SG�� {9�8 Ԉ��ȿo��G�����> }�h��\�G�վK	�e��uU��Ό�'w\),��cl�\���9�.J��qԏiP�k'����l����_5��`P��Ҫ�!�|���_���s1c�t�Q�e�f��Yfi�Y�e�f[�YVi�U�e�f��Yvi�]��f;�Y���TyV�4;�L�x�����G�K:N'MG�8�2����+s�~faoD%�I$�f���p�RC���6i��5&b�������x��Ҧ-N6�,b�.3��O�W�A�$?j��GF�r����'�w�����������Zp�^m��h���3��|TCxS�/[�s�����cyd�̅��ǅZ�0Chj�,��w��O��n��ʦ�1i]��w5�*A���r1��bdh���(N�C�%���ėɰhf��|�&!+8A2�@d�&pB���ʛ_��&�?�����
b����[�=L�,����%SQ��La��?�Y?�;��wT�r�~��[����hU"�
O��[+)Y�K^G�T�YX�1m���P�K@ҁbKaA��B �]!����5*�>�`��DF�QJ�ʙ�Q:z�=[bi��m��<�<L�k���ؒJj��&�f��ea6�7J��b�&�jW�03�I.MP���d2���|�Q����3v�t�6�XPYK	4Y*i��O8U_c��tlfv=�e�
����n[O/���!����8��iA�=[���_vvƎh�|4�#��M��G���w��Q�<�$Q��dWF���l�O=lP�^.r�#�9���x��Bh	<v�� �~�-�	[`���<ax[��t^lnz��PeHg��0�"��0#=r�����!�%r�^fj�nNsc^dS�M8!�j���1u<��.^�P�7)�)��ȵ��ώl�Λ��&�lge
�2if!N~����u2���ɣ`�V�i�n�436vC�LV�ʟ��e�	&ϬG{\���HN8+��)ʿ:�+~7��\��P���T�5O��.ڤ�-�����@�bG9���ME��
6J��Utfa]��Ƒm�R3C�ra��3�B2�Ik%��o�<2Jϔt�_��Lf��,`0b�Ǟ\��?��v���w�Gl��F0!D�{�����c�����H�Y͟i�`v����@q�uV^)�{ܼ޿��唞�.A��F�k���L�a�<J��5A�ӓL�)��u����R����1h�˵S��6�0]����f���iC�ט64��0e]�eGl�d}������Q��h�R'@��:Q�@?:!�S�w�xb��@�'ϒ�--���1���x�~�|YV�B\³ۡpz��5�^i��A ��"��~��"_����kmM��)�Fj��0ߗ���H�/`L׼)��L{F�����d6�Y��e��K����DƱ#�&��v��ճ��9{<�9H�#A�y��K͊gO?��U,�f����(d��(<{��&��Z�v~e�
���34<�
D<�����OV�'��<���_��c"pLy�:x�5+0s4G��:u���}Pi�;�jy�����hD�a����]0& ��~����{� �������)g0e���V"_+a��0jOܯ�'=�cOA�2!�KU�.6*ЭQk����xy��c^�g��{��?�ř���HV2�Hϰ�ǈ*�|,���0��h@kGa�m+���;|6ߓ3��� �`!�&M������A�X�����]�ߘ�lQ�F�mԬ�Bc�T����_�ŗ��^N�=�b���H�ϰ�1��^W�i�YD6��EZ!���m��E����bG>�ءo�X~U��uF鐶�?]+����$�2K���������1��%��[�50y��T���ܪ}�q�\�ޥΩ%,08[fy�5K2
��2�C�C<�Hl�������	�!3�I:oD^�WKx��-z�L�1
�S
 � �;���+Ƭr&��I=���G�i��1�$�k��NC��4�+.�����ǌp1c�e���ęM0ʅ�V��ʢ���C��L!N�r~�:{u�����V�3�m�
�K+�d�~���
��5,��o��.C ����c�,�[<tX}�{���G�oBR2� �K,�Õٔ�>��Ϫ"cHJ7��� �w���\��,D�o��w�0����'�H$�P�c�v�;�����d�v�P���@�[!n�-Fv/���N��ޯ��/_X����Ar|��Y��A
"W�'�+�>��wT.���$+R�-��yF��,�O�JO�X
�1	��kw�t�=v��MGzF8��V�:2���S��:�՚~����z�E��q��Tq6'nɇ���2�m9�+{Rc���t�r�xF�ؽ�����uh��Ƀ�
�hd��'�k��g��B9����>Bp4�V
�/aB'���B��L$����'ƕO�͜��f�e�y�;���C�˭y5;�MK&��᤭~
c�z4������#ŕj�.��0��������1��ӥf�1���-���_�4`=��Q�d��;��Ĩ�7.^C,��,6��T�_����?bRV�<��HGNa���}���&V�F��-�|Ԋq=�������y�栁S?������2���]��H�>r�X���͡\4B-"��|����N.�i���c�ST���y6Y��1em�v
�vtFz������-Ԗl�{,'z�1C6R@4�<v_Zi���ڗ��6�N|�va�V����`��5c��쑞L�U<��L�։(����3�zR�i(��%b�mԻ��Bp*��UЖ1���T����� ����ĳ���3�?�4� ��XV�����r�{��]�T4Q^���!��/&�0�L��*�T����_������Y��t����
e���y�tD�$�����}YT���Ҕ���/a�K`��@�@2\GE�:ᮈ2���4��K�l����W�6�Y�:��0�@u�cW_?�x(��L�G#�� �е���#7��g	���6&��g���rz�S@�9~���_�6-����b��WIh���ͭȃ&"*�����&p�{�i�SP�B9��vT3s,�s�T<m0j�ƀB� �B9g|���l(���d�k��0p}
j�=���=���QΖ�{MR�l�R��� �U6�$��)���?�M��MB��u ��9*�gs�g-H��U;Hn�wݛ.?��F���?�-'f�X8-� ㍈ �6�n���?�D�R����wza}�.��N��7r^S��mgD����𐿫Z��,����:��M��y��<�|yhd�S��֮A0���oF���P�����(֍��� ��)D�����c|�>�GB`:��o��<���5��܄=y�sDnf��P����_7�C� /C��wȏ�a�a�y$3F-��)F�`/P���x��?Q٩� �@'�[�w�=li��?�F^��gߐ����4�Y����3l�{Zش]�}B{���i���~��U�G����?�V����Ã,�
7�?��1�M���k�e�N�1�r�o�
 �B>�!�o�i�������m�T�g���x�]٠|��(�V\�B3�e[|����=�I��o��A�&ԟl��c���_H�g�~ܷXx]�W�7�c�m����Y���:iBO�f��.�M��")���t0bvͲ�dq&o��b�-��V�Lã�1�X]3�=Gy��ȼ�!�cfO�Y��(�aD�8,�U���oa�g���7^���;}�C��B����f��#�����-!���$9����{�lfD�Ct,����U�H�[��}*ĳh^��]@�-K��%:#@����f�5�6&k�e�I�$ Vk��Kd��;[	W=g��}di{�˃O�p�2��N�Z^!��@��f��[���C��v(ş�XE�&Qd4��m��#L52o �&Yε��_] ӏ�E6r��i�%��i$�w�2�g���m�T,��K��H�'à�)s���4{`V��餉�/	G�0a�H�/���%���u��#��lf�� kMF��M�	���ŭz2�p��T�e���d��3šV߇�5��ʌ��+<	��w�1xpn���LP��������M�y6��H>3��v�/c����w������+�]NVz��6��_��"�Ս2��o�F�g�he�~MqFE[������m9����=$>��}�^���2Bk�ұ�����U���GDVt��TI|�Z�~�^N35-Ǫ��5�5kcŨG:YԻ�j �ZW�}cpW��
f�]�m���(�ϼx~�����h��1M���_�Qᘺ{t����`L�T��4�4��G*���dv� B�Tf�5��/�$k^B��pC�C��k���3fuș�ݹ�ᬱSs<况�X�T8��.��\�dضG���/� �T��D ���e��K�_V���<Ʃ%>ڹ~��AO��&5 s�P�^�0M	f��t��w���b��/�v��hP��q|�:�BC��ҧ�����(�J��n�cXrx#=��e�Ӂ�������`��(�M.5�BQ:+na6��X!�^s���V�p��I���Cgy8F�O��xy:��R�E)��u}.����(�#X�qV����d�t�.����O��o�J�|��Óg��<�|�
�G����(�ٛ�cg򕷷�%PPPie���Y��u��͚��}6-�(�����5@�	K$@���7���uw��/S�����M?�^JO2H�a'h���r��Ԕb~�Tg'�{�����H
$�����4��[I��#^]�qK�9��#L��sd��&p��/0��N�BR.[+�!l�mc*ű�	Fq*���m���p-m�P�QtA��Ѭ�!���VY�^�.��Hk�t�,ο�����6��\��z��KC��:�r��s�b}���b4��v?�+��G�I*4kq$�q��cV��Vr:F1��"~����영盌L2�[8��������Zl�^���~�6_�](g`->\�6I}�q��0�l���C�|���6��������Z�j�CMf��ҙ�$g"��;�JvP���Ճg�(�M)g��X�`g=�������ا�&-'L��3�si�3*6#6��ne�`������|�-�t鿑�,PI�r"*?h&��鐬S���C"	:^P��V
ټ���k��y���y����yf"��9�l��aŁz�D��a��|i@	/B����e�}rQ*�2�����Ǟ�&�ï�ٯt�(~��~M��܈�~Y�H�7��z�e}���'~��&g}�'!�k��wu�5�Lְ�E�����V�o�*'���]Tӳ��g���Ϳ]�˾�]�
�w���$����ɇ.d ��˘��⬇b�\3�"�n��ThT�X3�G�)�����*"�C�u�h�멜�쉘Jk4�͕�]E���(�ZCL�����ψF#�	�]�Z��'��r�O�2�x��i��5��d�����K��n�S�m_�LB�ǌI1�i�Ey��l&�Vf�#FYd�"f%ڬ��I6!B� Qbk[�-jjv5���J��"m��X{�J�}zxl����V�P5BQԪ��hĚ��d���g�p��}���dv��s������ Y������Z�d�=j��.�e'ft*[�0_����t�Iw&�v����B�[�sj�s�Fל�лJ��i��#K=!����D�Ы�b��� T��qޗ�3	��|���PG�����?���.��ڐ���άA\XN��l%�c� S�gꋝ^��	_�N�=YJ�65itx7u|�0�|N������nJFp]�9_>��ЀD�߳p�� �H�ku��/��l����]�ގz)ǔ��jd>���L�Di���}�V�'�����C_ ���N������~Z��9|��,h�5Q��>}������L�m�y!)���AN�	zgq6]'L�}��tAF����GuE�?��M��u	}�t��M_���wiyJ�*{Su��z�gB �*ɲ�Wk��aw��NaaY�,�)�����+��f�����M:��yd��	6���2�V�6��ؗtӃ9�A�k[
#]J�Cw��^�������Y����-���I�jI�_���8������n�df��I�0�sV�t�{�-� YUX�3���������m�ݻ�Σۈ�{̩K�GNy|���8u����9���]ho�x7���$�eaP�)�8Yy85�D��2^B������2��.��e.�'�\�j�˄�eQ>�W�O5�>�~P.p���7�H�B@�;Qi��9�`���7�`���2��U�������$٘����u/���Z��vA�_�]&7�f�ZBn�B�<Hw���'����4.�6�w�������]���H����o�T�eQ�M�4�tm��l�R��nZ��s��MB�E>���=��.��f�<\ԿI\�� ��`S� �ڗ�fiF���w���*ٕ(�_��[R���H�f�3�A*��Pu7c��Ɲ�N�"-��J3���zB�J���p�l	N�T�2�]��&��i%,���n�)K�j7����6o��%0B��y��ѧ N��$��NSI�^�i��ĥ�pq(��4�ٚJ���.�FQշ.���ݘآʦ�����ȣ�zY�1D���6������?���< �f���II�m�ek �]]��A!�WhǍ�`�/i'�1u(��GJ���X:m�J��ƑT��Ä��ӷW���}��+��C:���ߌ+a��]��O���D?\ͶY_���XG��R.*�1�����U���wD����<ǒ>V�Uq���6��+��'�������TY��?P�,m_��\2�����}B(uy�����<��9�4�\H�����Ǿu%��|z+�q�;t�qp�hBv�����|�����|ebS����I��o�[��5��׼[뾍����*���G/�$b��ưn����8BN�׽�-��6nz%16��� s��'��z����g���.��!�~$�˴�+�����MBd��ڴ��"��{�C���tk�,ݡ/�>������K�W������b����4꿚�U� r鯟A��\�&���VL`Pl>&��N��o���->�żu4=x�Ҝ��}
%�<���� ��^h'K��)���k�o��
:9��f�?���o �j�zd�:8;�N{'�D��5;W�'���a}����C���쿃㚪�p*r����T��{y�X��֓�h��D�1S���9�O�x�z�5��J�}���{f�z1��-د��("�V�KAEO��t��˷!h���H�<�ʋ�7���xd�X@,��6��~W�K�m���ou+=���~cF8���ӞԃvM�W�}�P�ǩߛ��K�#)|m��2�j�9��Q�_����M�8�|�0�OP�Raw\fc�1+�C �W�_V�d�����0�RZ�x�B�5�{�%x�t��$Q8��2j��{��D���"��Wr�r���ڔ�d�_�@��.܄�W���&L��[x���/�0=�`�p6�����T�-yBz�Y"LҕQ(�A��68>�`�\M�?���%��ށ`;ˠ��E�4���/,��/F!�m,�A2J��\����J�"Q�M�4b�� }*@�I���}p6��E�Ʈf�Y삇�
��p��Ba��~�帔��8��VF���"�`rb!���6��+,�'���?�t�]�0�#ןΌ��nf�|`,W����M�Ũ��fɜ��ʄZ�
x�å_ziM��������(�ęK�����X�a��e�?��7YGfE���������+k���̳�s��;8)	I�{�}�"������X5�b�A��Zj��
"7�0Ы�X��bB��˟�e�%3����f} =���d�S؇���B6����c��
��� ��ˍ�v�H���e@�,�׎&�Ev6V~?G���^�r9����$�А>�+����;�zB�
��9�%/%D)�~c��H�8�2��E��|b��|$|(�s����x����+�!�;�!�Y
:z�~)F�YJ�r��%@�as%~����GϼT���fj
}�~���Si�Q{�nףU?�:�_�*���3��I�Q'N�&�"��c����U�*8���^��\���1j��*,(h�=!$�9*Ɖ��Tb�8�/|��k�w��5�~�[�T���c�CB�L6�I1V�D�{�KE}�R~aW�����-Έ�R&_�ł�����#|"�Ou+-�i�����Zi�^��U���FR	����)��4�����ID�L#s�]���ފ��b��HyP�3�N�>3�农��Ɠ��gs~r���^���,ujklO���]�
��ْ֮5����
}A�Xݯ�`<Ǵ��$��vx�E��e	��?3#��פ��5��#��&�{&o�^������dST��t����xFG��A��[i�ž�8��衍q"���L}�VQb���R�����	�U���p�m&g�;C_W[a��.����W���.�
�i�k�0�;1��:^�d� ���Q�'e+J�L�9�.u�R�R����l������r�)ˆ{����_Q��7��c��T<k׶�OX x��w�A�����
z�ۨ�,��k�0{�ߠZ�su�.���]����4���#�2�q�?��p������#�a���v��C钡����f�E>�z�#�C�����-��)�oDA �n�џg�P���g�{ �F�����_~���ENT�!��ys��WԺLK��m�?[��)���м7j�}��ּl�4h|��]/��<܄��ͥ���~+�c�(�5�3�ǷQ�%�-'�f��4��T%������~�<; "XC�h��%w9=����^�K��\�OG��V�o8�g�,�sЈv�-W��֣B �b֤\0��A�*u(-� ���y$�"�p�,K�w�ȋ W!J$1d���7$]�2.Ѵ�����pa��HE�ᢁ��;��?'뿤v/�Y�VwI;A��0Z�֊���Ph��5}$Y��	ѣ�=�!p3�ؕ�{
�a�aa��L��b���{�ʾ��n)xm�.%��ߕ��Z �,D�x����-<��Iy�6��I�����4�t�`��6|,+�;9���JS�2�<ò���kԪ8)�~)�Wy�;�X��?8�l_/Ŭ�6���?�,pG��C'M[�O���q~[�0�8�9d�q�Þ�K|�f����GOY�7S���D �"ҷo�����Ta�S^]Ϯo�>7��'�����]㕙�3{�Nm��8���I�����7~wЯ,�������vJ�$7-�ݍ�>͜�0���9�N71~qlR����ӟq8h�%B�29����Ń��x�������� �ϯ�u��_BW�2뷙�W{��b����F�j�ϴ�(�_t��O���q? 
['O�ߴ'���@) z
��Խ�,�٘�G[��ݳ;�o2�����:��ab���$<�L�yg�Tn��]E�@�۸�Ȅ��1ST�l�ȗ�+-� &䯂�?'�����"��8������R�ݙ��֞�� �ʥ��D����
�:��1)XE
�E�Z�YF�)
uD��v�:/��Yx�ު-6�\���4ӹ+�)�Ɠl�7�B��WV�'\b�I�uj~��,�
�*G�͎��4��(b��I�K���SJ�s}<fݡ{��Q��Ls�#ѵ�h��p�d@G}��h0+@#��I�ƾ�F =~����'����B)�Z�<{wV@��+����+?1���nm���>�јxS�?i��%7��}j����5&L��m��y�%V��7����'R�k�4�����F�Q<�T����u�*��r���"u����g�z�]>���4�$*����h����L�kW����Ti�����O$��>L�+�6�P�يD�7�:r'5��^C�d��]pjc���9	o�����z�N��_��y�� �׬A<P���K�_4CV��&����s�a7О�I���.P�s��#r��a��/H� ����n��x��ð5����I�?��� �^�i�
{�/��B׻J$�ԧ�����t�K_����ݚ'��P�R$Ҝغ^��M
�"7��^�(��R����d{U����336�M�X	���^jF�ۘ����W�i�Js��섛	���#"=v!���@��	��V�w�I�:7��̩4wFk�m�t
a,Ro@��񱬐.J�p�I�ju>�̯4WLNm�p/����F?.?�&�(����sO�����xߖ�O��E�`�	�_�Q��o��Ohu�z!Rm��!WG��z)�W���1��w��[��f���F��^ځi��/e�S�k�[�����;޳2ND�P�i(JK�i��\�M�K�*ނ�3>�\��@ ơ���N�m�Q~E�Ui��`�i"S$zU�k��JK���8�4Z��}�.��p>��췅��ۈ=qB�JsY*4 �h*�\�@ ��t�
A�E�O�/��f�&i� �d�5�o�?��a��a��%۔��i��u+�rg�������ң���������ܒ*�XQA$��<�z�7v��A���$}i��W���V~_<�/�м!�Tgm��)�++����)�j�Q�*�¸��W���G��,�p�6�ng��}3��I����_�:�m��~H�E�	쪬K�Tm�Yڴ�w��'m�W�UeC=���ڵȟh��״��$6�r�y�,�ߗC�H��`M^���>�n��ơO�遱?���E� �ݿ��a�X�D��*��
�����"��ή(�%���2�vN�^Z�����oY�C���Wn׺b_ǟ����z_��Į8>���0��<���RZ^���ۑ�W�����}30~��d�A�$���,".�}�eM�6C��4礅��Ҵ���$O��Ŵ7������)��X�&h�(�/���[ʃwCT,O�n������m�!��k�<=JK�w��#`D��Y����Ơ���AhBXf��{��X�F���\�����ɞ��h�~��������H�
��1.:H����	�)�I�S�>�L����p/Ę8w����?  �{��pQ�5i) 1�C{UݝB[�9���y�lY��UZj�NK�����A�F`>����h�`_���U�c��q3�7��x�n������dv����@GL.��m��/{��jG
u(G|����xq��=�6ѨW`�j�/�)�U}I^�ԋ�d�<�@�Oi�8|40w��E`y�<wUS��d�$01�����G/�ǌ�9Ul�OhqvS��2�`�J�;d7Yc%�=�����1|��;�������8�!����fU��U�h��XGΘ/�bH��|W���CW���TScsE�*��L��igAt8c��̑9��h��ε����hΤ�����~�(I�����J�+ϐI���%q���+�#:^2l=�NRǴ ��|�ԃۢeV6>��4l���d���<G�Z�Ʒo3������Iy�Y�����4�B����>�� �;�~�J�rw`.q����G5l�b��Зr8]��9��5�GiKfl�F9�^�TC�`�Wu.��N�4�Z��U5 ���WFKR��u�h�Tk48�8t�Ҽ 7���5n۽��Q��M�*a��j�NRv���ߢAO9��*+���qx�ȣ	RkP~�*ݡ��=��ڣ9wO�U�����Z�-�~� ����io�ڻ�OJ�<5������rA�z�)��Pb��2"tӱ�mM)8'� �����t�۟�Ȣ���nN�[�Si.O����U�+-�)(�J�ct[�OӯuG�Ez@�vx%\���?*s�:�+�"��4/�:>�e�RP��)�@�i�~��ޤ��'U�h�{���É��oH��K0p��d3�-�R@kY	�a3KR�Ij���%^W3��o{'p�a�s�T*�b'��
�n�x��s?�!��1*��BE�|3�O��kmZ�hQ��rIz]����x�Q�w#�S/JF�n�@��xJPdG*�AG��~V�if��Z���{R*X;5­�X�G�6$Y�>��Kխ��2��C�	��n���������w/I�
���� m�� ��T��T=5g��/�E�C�q2m"`(��"t�V-�oW�Bta]���K�����O���<E>�.�p�s�1y�:�PT��(ͫ��r7�:p��h�Y��CHe�������85�����H�!l�}����M��)����i"���V��&�u�/ 6}+��n�&�[�	Z5��eM/?F"|κ)��z�����}K��9��q��4�i��vY��(��V��W����=��.�D�AD���I��+�i�]��%���[i5��7��O�{t,c�����8(�D6�DC�@�ȗ6H�`g�Q��As_��<T���j�=G�ˡuRfD���j���&��)Q�8����X�8�4�9�g��H{j�=XH�H���B��I6��(f}b���t�f�):��̀ h��@}������?^/�4�Y����[��-9�${[�Q��U2�X���n~�L���,��J���갬D�.,=.�S�o��}�<h����	�y���
�A���#3�{*�N3��P��&\�_a��#^b��2C�5�O�g�Fk�\j��D?[+���U,������4�Z��Ǹd�h��N�	%Z�\�����u��j9��O����bta���|�oid�#�+D���-��Ң���֓#	-�����%���(v��H��ZG��g�ګ1;�k�,	��o@�If$�<wb_2C3�{kA��	�_�<��x�D�K0�HN�]��	n���z=	��U���-W;���4y���3�a��od���"�!:ȪDN���Z��I���W���$l����d���z�'=�Y�l�
�{��+�~@�>uÙ^������ip
��.`��9�R���/�K�zA�o�B9I<�MT\	ҸVk@r#�C�M�� ��b-����yŰF�a����!�i��1�,4����5�d���М�U[�<Ǹ��Sι*!�!�<��}���YP�}^)�M&����C�J�V�팎S�v�cs��|m�q��8e��RiU�O)�f^��	�I�<��#�@�Pp	���]ƶ�X�[:��
C>���e��9��uK��rG@+P��&S�I8��ȼ3�u�-&�j���h�D�
��nh}"!YN�+�2��-�zÛ��=���� �0���ۘ����-�
r�8��n�@�b�b���5~�{����D
n���lj
υ�Xy��
u�$��<�M��Lщ\~<��X�f�`!�ŃlU9h��+�Cf��" ����y[��d��ҤI�'��Ƈ���j.<�cko-�4������F�͵��\؞��c��ko0�1�����<ڙgU�Grp:9�Ϗk'�]����a)��#5��ے�Q�Zg|k�ćwM��HE8�����xa+��c���G��I��y�t�gNd� @��@g�I �[����Rc�99��q�Cb���Fo���+��;�,O�u�J�U�Wo��� �����Gײ4�d�A|U��U��>c6��?A}J�Q�)���]?��'��0yZ�;QE�t��`4a���ʱ��2l�zl�Ew&t�!t#v��/�v9*���ǳ��,J3aThՐH2�/t�$#��|}y2�ΜOD����3h�)��Ra��Z��#Y���^;����C��V9�LA�T?g�/�-�_��T���I�j����W����'������e�!��H���#���$�O#J��0����~խ��D��/�P׊0��PΩ�9���O?��ws�hZ��6���Ω���w�V
�nv�@v�pyg�M��s��7�T֊��٩��W	0��`���h<�?�`#�6�E��،D}H���k;�>'��9��6���?t��I��$]�2���q�,g(�����ϯ9zg��|_��(�ˏ�/ZSYT��>Y��3���.[$�],C���Y6��.�o������ f���i����T��x&9����5���_$���m�K�أ~��21�e#cB(S�S䧉�Y��\������!:حr���֩/N�[��7��"Z�M�,<p�Igh/K��`_u��#O��epA�жi�/nJ���/x�y�d����u��w��T|����q$�0޽���p�o�������m�?����nRV�6��>�������c{�s�&'���	[�y��e��p_޸�_�����/i�rѨ��/ej���qa���?��9��0}�}W��VסS��5���Y�	���U]n���B�uM}�۹$"kh��l4�V)���"Y�?���亞�v4����e�V���":wbq�d�64�\uW���`�t��u����A~��R6�����r�!�Ș���S�@����_��(�f�)&��J�[�A�Y8��$��x�o�:�B�F=e'��GŢ ��tTWw���?�Ǖ��eԛ֗fH�S���u}�o�����D��Φ����]uk�=�24��{*��
%w*h�5�#x���ׇ'L�+����ӫc����̄��B��P�T�6G�A�?^��	t/"��,���_r��!@�~�������_�hX���i��O�+i�%�s�L<�j�%W�@��Ժ�H�v�X=j�g*m�//����yǉ����R>�]�U6I�S�e6���L�e,?������ğ�6A�J��Nr-7�z�{6�&�׎	�tv�ʕ�[�Y��ֺ��d���If|�t�WzJ<����w"n�H��l���<���ƓX�̇��ܸ�Հ�=�D����h�O�1��z����+Js'1|X��H��o�Ӵ!�RrI� ���2�ZR��#T�J��Ȇ#�@!��=�:�8�?��W���_�5��~�D�*���&� +9D}N���*���O��Ϲ\�ˡ
 Js��K,�q��c�lA�im��g����Z����m��}�!��Qi�7�NE�R�|�l�t��L�wsb�z�h�a�I����Ic�wѸ�e4���4�	�K�H��o<�����+�m�3��&׉�.��'W�r{���䯝T����?�X�"#��3L���2Vzh�>�?-A`'��N�_�w����&� W�Z?����I���im� �H1
�,��]���Ul������듰B'��E���88seB����1��鰟����L���0w�4�=�܂6�����{8��;�[����w�d�Q���3�:yJ�:�����,�Y���Py�*���5�H	V4��C�6~d�!}%cu� g3��I��r�>@c�pB
�W����E�w(��&�K �噹�� <2�1=7�\'�)�SW���g+`�'��~����Liy#'߆�� �K�X���	O7�r�������~|�p���Σ�����A�#�w�Թ���o�����(�'����r�+X�2�-nΆI��V�U[�I�Z"���p�x��w:g�%�5�'��([Kĝ���5��}���Q�n,�N{�^i�h3H���i�;5t˖�w���%��8��h��W���vh�����v��d���ؕ�[�,�5��Jl�t��8ЎҎ��@���c��X��
1�.S���MTr�@v|{r}3MӺ��M{�Hݎi���=���|���Oi.���8jkX�`��K���Q?�Ƕ�<���v��*��W)�+&yڽC) 98�lb�C
�g{��4���A�� i�h�������gx�Fan��-��?��W־<����۴W?@��p����N=鉝K��WN
�}�U�����zm���)<�F ���& dH�4ae�a�L�y�LM(�q��9Ԑ�$P�$_���e���$��*Q�B�4�װ���?���+��� ݸ��s��8�AL]���ָ��ņ�W:�RX����bNmIL��vm7����7�^����#WZ8���.�9I�a�%�x���#����W7����E�Ag����Z��H�;��J�D�m2�S_�R_⿝�ߨE�}0*8��56�z�`F�)T�����f4?]�������ᔁn�>���b�a��{Y�v�;n�TiO:.vX�7�YY�^�~l�G���ÿ��&u``��ρ�jP�HR�Hs��ý�{��ý��B�u}�]_�l%Ǎ�8'ԝ\�W�_���B}��L�� ���c�ǻ�;T�������Տd����Ώ�C�X�l|w^�l�����2�����l�s,~p�q4Fo�`J�����]_L�aX_!G�F�ܡ�k��q1�I���Q0���XY�X��S��!��� �N ��Z��0S���i>�zdVC+�c��`s�u6�d%������i�eʢ^s�ڐ�1m�ك�qtV�'�_����] ?��Kܥ��`=��ؗ>S^�x>�<��9z*�۬����-'���J�}փ:������K��FYҋ�-����GDe�h���G"�}�&e�4ƛd�!�;QZ�'�:;^�;[N>���/ ������\���%U����˳L��]�Ok�7'�+=����/����Ƿ	ސ��kK�J�B��_+��R�]i�"���-��kop����j��(Ⱦa�o�������|��lj`��FQ7�y�:�A��(��	5Y�� f�����y/���9p��Hq��Z���$�x�?�hE?C��f��n=o����lz�^����l;�)M���$L���m��x�&F������5�X���=)�0��l~��,�+ђԫ4;�=JSsJқW�MV�4��E�Y#��ܱ�c����=���SZ86j��/�2k���Ө� ��fD���}Sۧ\��Kn�����ܨ����cZC	�%�o��7�=�q�AN�Ƀ�{�\��t���Ȟ[�oP ��@�5e�i����6e�<��,1�LN���ݎ�}]k�6�P�i�lHW����G���xP�3W퐔g��wMWO��Ӵ]BqH��V��ŀ?җ�е�Df��R���ʋEiɥ�47�yFÝ8Z����&���MND��d1�X�a�߽X/�1��D8�ѳ��t!m����K2�u��`|V��2����X��؅�x�E`��<��X�Wx�=V��(Uyqjryu|���E�R:޷uq𱌰��`n�L��4_���< %����~f�i+=-∊�'݅�,J����4DxRltd���&4��u�z�����#������Z_Ǡ��>,�n{�í�.�s���*i�1D~��tɈV�}$;��2���IOs�{������m�r��t�W��g������d1��+��(��x� ҝ|,��{)���a����u��q���+c�����5�>�+a��H^�q��z)�V̗z�c��X�e8��I�ˇ��dٷ�jB�t�C���c�yj\���c�e�*��b�7�T����� L�,hg���p&��|��G �p���Dw
SȠu_r8N7�o��s�~������>PQ�YjS�S���#�H��Kȼv�k��_㢇BR�MtF1��&^x�r)�~�6"�c�nS�c�7��傽�����������-+D�&�dm�&���%
���z�,)���;Om���B/_�ʵ�24K8�vF!W^D<��Qʤ��2#r��,�WҞXm�Gq�Q�񷶉xzn5m�̌�t@w��:p�-�l`=I4auj�7��Mt w|H�m��4�6�{�iޒNc!P�)�/��0�� ��0�oIE�1�	[�h�1��M� �ݠ�E���G��t7v^��M��ImS|D�o������Gc��λ�W`-�q'B6��V�c%��9q�fCi³��"�R�Xv�	��8�4���J�z�,Ө����G��;M�>�c��*!{���_���!"��֌��B���l��,Zi��"x��z;'8��Ert) %o�1B����Tu[L��j�v0��X��#���Y��H6^H4��Q�}���Z��t���8�	a#�H�*��i��`41v166��/��0�yD�
`6ٮRm��JN֧�ǩ��w��K,�@i�ԡt�΅�{Hɱ�j������/)#��Flc�+&`��ޮ߈b�kv��ViW�e�'��Iw)���A�O'Z��b�UĖ}	{��:�0!����H�U����BY�3Q���G��[��p�(��w�+N�3M��&����4C8�2���^i��QBByC����*�����5#�3��a�m��=�ړ鞊�-s��Th9Xk�]3��Q.���d><j�^iQ4��	a��������G�Ā	�c�S)O `�@.�� �N����y�R�2G��:>��OD��$���o�@�i�~�Ŕ�_����2`�2����N����P���Ԅ%�h[�sz����Y������H$�ʈ��!�r��+�5��ie��~�|>��n��D�_+/����{�g�w�IHF��Fg�p��!� r��?x��&������%F� �-���#hƿ<�	��;�<ǖ��s���h��N�Yv:C:$]�������N֞z��c�`3�+�eW����;/��Yy>��J.�
E(QhKx��v�W<��>���|7� >�S�K6�FA2"	q�"�HЧ�v�_!2C�x�i�xH�֧4?ܻ�����
��#{Cg>g$%�c�ʡM�+Q�E��i�a2Kli%�9GO�b���KG1��6e���'����j�s�y?�X�[;j�G/֎�{B�igO��3�$L}�VRĽu��3Y���M �����Ĕ�e�{} �lៜ�_��f�>W�ힽΒb,���J� ��"�[�P�[�mg��Y����cN�4�&	3M�L�@a��\/u1�I��ɏj�|��H��N��Ӯ}��?آ;�e����p���"{�S!Q�7:<�c9��֡����O}����sl�I�k+m4K��4�C 0���;jb����nDuvΰ6�*�G����̐�$�-��4�=���ו��"l�sQ�v�+xW�
����n��l2�*����^���u'RF��/�_l;�m���*m%���(s(�^2������h/��/��З@�8 ���*�
ίΊ��Rp�^���G�ֹ�����vT���#rAU�=��vI��B��\]z�T�;)M�.���
j�
X��CdY�<W�\H\x_��*0����JRǆa�h5��/Ys)����j1r �d�&�o������	$<��I�x0��v�d	^��U<��m��5���Ag]�M���N`V��Jbb��o�W�!�)��p$�-�S� �����@�V�����3�q�Ǥ���6~�^�4aF�����
�Qm�i��M�}@�f��g������!��]Vx��to�r]�VZ�(9h�!7aҹ+H:�{�祙���8���WB{H����(5s}@`��'���>d�/N�.��8���%�|0\)H��Q����`���MmwI�
{sT~������;�_�⨮HT��u�'���,�X�vb<L��Ր+^��`X<>�0��BW��-�VNW垼c1��J�+U�N�����'���K��1O�џ,?�nE��>���3�J���@@�H�
c՘��.(`�nOj1�u�p����;�ju��X�k�~�e���)�]PJ����}��֝�L��]�[VʌK�I`��Ҍ`��=X�M��-N�:��S����e���;l�9ѻ�t����c�h�ͳ�wpB��c���R�٫#Xui�d�X���.B�~�I{d}Q�x$r����q�,�ω9݌MiD.C�����t�4��/c
���`�S"7��\����|�G�LR�a$�_�E%� f���U?��oK��O;�'d�=�.
z�Ԛ���k���:�."��f�2�7Ib��̉��j7*��0�~�䙝SD�ٗp#�ĭ�+��3�0.��'&4S��m7=}��G7s����f�g�qM��s���Vz���Si�}���\:��r�&����h��\%rWB������ax�:XMc4el���Y����%�zT�v�K�:��hӗdF+\j5W[�2>Iԋ�3�h��E�_���jH��V�J��S�uj�K�hؽ���FoD%�\jI=��x�^��i�:���o ��!��
���F1��I줅��x��x�4��p�y��$2�)�����5�87�@��C�[4�~j��}��Q�5s�'������)�Av�#O¸�/���%�anK.�}'v�0����N��qy�^������\����Qg3O��L�~�����Ȗa.�賄H�����L�V1�
��$%r�+�_fQ�)��[��:�f�b!m���FߖX1�;�O����d��D������m���h��#TG���� ؓš�+�W����%
 ҙ��E��/��b�ٚ�{��׎�����4���/9e�kٿ�)�j�b�{N��<�]�#�4�?t����I4�$��2]��� ��b~H�?[��t��=��t�\��w�N�?P�/��S	�T�8$%�?���Q�����4�i'x��TԬ�E���]m�h�^��O"Q�č���ԩ������i�i_J䛘�+Q9�Ԡ�G��P�g38��ĩ�b Y%��4�bZ��?�^�M%�JX�֋l��X�>�G{oʔ��H��6ߐ"���i�1#�xG��@)Ju�j%����W�ySڮuy�T��F���~)���_'�&Ikr	�⛑�`�/ND�́16����4��=�ޕ�u��u6�����1��F���
���J(;)W��lV�<�Z'� �KD����ɶ�p]�n@�ek:���w| K��
��ve��ev�zﲅ�ߞ�-��> �`��zSiY2��-x��&�eg5������*3R�P�fm�L�y�ѿ[R��$i|u6�_�3�ѐ�X�|��/��Vf��r��|��"���BG��_�����DG/��_������L}���Y�sV	�t��R�>�%�tM�?��A
��o�#	�6G@���~Q���YF 2�`Z��8(?�����}Ylt�	���@G�E�&
� �ݜx��v�����ޔ�Bi{��ݔ�qՆ�O�q��ZT����)X	��L�b[�):���b����,���D��(���oK��f��t}2	�h���Xi ]Ư:�G%}�|��&gLIjg�yV��6��b��d���T<e�9Z'�Ҷd�H+�kn���;���o�� ��@�f�&:H�Bh��#������-�>�)���`�����YZ�C+���e��M�&���CN��u���7iE��Ti�C��6�{0x���@��'.{���%����Wx�}��U��䏩Z�-�Cj�t�ѭ��"�I�1f���
-�y!�k�9l��ukg�Y��Ə6	Jo3l"(	�~��~�ҥ�1�ٯ�~+c$4=ch��R9-p�H�>4i\ X����آ����|:@��� �Կ�I	D�[�u�*k���-�D�ni�XĹ���/1��1�����5���{B�s	���>����EeZ��� }�Rڜ��j��eq6]��F���C�rH�`����_i�k�����J:�Gr�+ـt�~���J\xU�]2�^I7����P�	7�*m��ަ<��TTQ��zT=B0C�ɯ9�,*׋jI�дL�n�;�B��sl'�'��甹�\���P"��X�gK�I5A����l_ũ÷���.7 �*�]�8XF���͢&�)+-%�JKB_� ����v)-{����m��Q5��)�O��=�3�����{�\�ǒ6]+!2ƛ�^�̢��V_��}�6�~7 ٝ��(�Ȑ��`�V���fԹЈze������	��h��)R����4���!H�RH���<w��ԡ�-�f�����?�6�>��&�x�$�Ə��a�]�xTi�1�����*�ޖ>��C�Q�j�T*ӹۢ�N���x��QaRy[�j����>ޭ��wX���;�]h�X?����7���j��;q���L�x"��g�Bloҝ�%�?Q7-И��� ��C#�d�������֋b=��Z���m�.5�ڤ�x�06�֭�.��߭4))X�����?$
W�y��ܸ �:�~%r� ��O6%�͗����D���ۗ�{��7n�+扚,@���J��ծI����C m�AbI[_�)~.uD��p��� ����k�]��I$�мg&`E�}K��ۣ���{��7*He�Q����W�[��;����=s��.�9	������ojo��3b��(&�OKY	_����i��ˋ�*���X,�#�-1f#y98�i���&��ѡj� +�R['cE���ZYE�2��&�nX�C�wx�ط�g+�/��7��J�N��1��!�*Z�S"�q�&�p�\e�!�L;-�4OCU�C�[�<���v��%��7ORZ�w��-��*l��%nKi�����|���\�#��Qn�Ic�tn�Et{��u��B��P��t�U_�t�i��KL1!��G7��#6F5��3�~M,mB|����]h�~w���OC^����m�@g�m��`*a�}k$���|���˓{;2���A���m#	՘ͅ�b�!���E�ٱ�a1���!vmT�6*8Z�+�R�A����k��hM�cx��x�C�����u�+�:�$�uJY�u����۹�e��n�W:�PA_�;��{Z�N���*�]2�v�.Ne�F�(�ܲ�b��I�C��L_|$��
r��ƁBmH�ECu�Q�`���p����s�);��_yW#����D�W��$��@��ձ��3����Y
^�������W�D^Wn=: 6Z;��T� ܣ�w� �`��p�K�'e��Ws���z�Mǐ��xؼd=F�?���L)cw�L�>�U�Pʻ�r!>��w%zۄ���e���������3y8]u��kdO"��n;�m�ǯ���;����w���!�\D�6~���-+D��r9P058����	풷��?
�E�/�3$�fQ��@{�������'J�>+_Z	A;?r(t����l�+t+r�'Ӓ��v�}� H�C��x*[ސLTa#�%��\	��/�C�~@�3�;c��݀<	A��V4�LU��r��u(m���xO���AD/k{�����jw6:��0.op�v�Q��.m9o4�sX���ٺ�m�Z��]Xa��u���欿	�Ι��nt*�%&.�6��W)���u�����ڋ��l�X��`#erݪ6{qd��+�W�{��:>MU?��/�/����_rq�Q��$hO��*#���2����X�Z�^���}=A�D�Ǫ9n��6E�j{2�ٗ��f0(�yZ�;v���+9^bE)����$��n�F���K��Wr�u�-S5�e�JyH�Y���;�0Q�+M���
��H��ҩ����Y;yƒ���xE%�	��*�e�f��K�ڟ��SnqDW��i'�yj�RMɅJ俇Yu���t�F��as�-��g�0�R\�1�w�k�p>*�j���?I�,��JHm�V�����*����*�J�4j�t��K\�vQ�k�{���9+�/k������	uWn�F��:
lxM�,f�PVc;��� �x��J�p������ڢU��sg�]Q��
�� ��`����������'�O*��}���=�n����,8zBi"D/���[�/�Ċ��%�n�"�:��)_2�xh˔g��ܓ^���؋M�$�`u����2%��J��&�a�Z�MR!�IK��&\�7`��w��͘o1.;����̍$:��~�m�K\Z�>�ĭ�14���U-���ho��#\�7�zZT�3����z�-�4~�w+��J=�>���/�8>)�7�4[.���j�Z��V�h~Q�7��ͻ��sA��Ma)Zk�����_�4!!v}Q`�x�-�D��U\PIi�ʃhk@{��ă�K�[���SX�c�I�M_n���(��9?D	֌N%��"�~��z�oe���c���,�5���9�[��[���3��X��?񑝎ZE�t�w��ޒ2^_&9D�����ɇ��c����heE�fi&"�����jl�r����\��U3�v+���<\�_��WZ� ��E��d^@��n�W��U�A9b�\�)s�-F�E#K�-_$�~T�-���U�E��т��S��&ڤm�N��~ך�&f�1�����1����}~Nb/�	c��>��N�?C�՜{$�dC �hD9��43 80wYLy�	�+���q	�\Kh}@}^4��W��41H�&���f`�[?O�S���#�g��k([籆��}ΰ�eN ���zɠ��+ڍ�(�}�����,�����Ɨ��DD~�3�jt����Ҳ�#Ë�y��3�5bK���4�c�C��aF�[7Y�U�u���8����g-��RڦS���t��i��ۖ�ؔܶh���4�?��K���&��?��!R��ԉ.$���F�S�5�w��P�8����+���%s�%�6ݛ��E�J�|�(�+�ͻfIX�<�o�l���&����f��h�Sq,�kfLr��t�n�ϸ����i��g�0�����u�tB�~V���ܹƯ�R���2���k]���ݾh�6�T���3�`�׏���Mw��.'hK�yzڻ�2��S�euе��V�֐-�(a�E����IY��Rw�Y�u,���W�*�@�O�������MO�$v�m�v�ߩ5���T��?����$�!�����$�\i+�л����	��<�i�8b5����e����g�fLz�^m2s?�@h�)�P;"8e���&��9�^w�?�)Gl�x��x�Y��i����2}�K}��*�8�>]��i�+�~���ח;hz.�/�g�җ8#{Cr|�֡"o Z�g�0ng}fy��k_N���!�Ƴw���k�����"�,�Ȼ����U���_�C��x@���Vo=�m��=o�����@��-Y��
�~�y�Kԇ�r}�^j1����u:��+v,����j�%\!���KT5�	O<���w�dT�7Y����F�a�Q\���DAf(-�����*���R_�U���iƺe���qo�I�0���&�?[�D�Y&4���I�x��"-`����b>=�u��RP� R_a0�(��/��zA�ѯ4�CB��ԗ���Q7c�ZZ{j�Ă҅�D�Ú��O��K�����QH�q�LV�ω�7����C���@��0@�V\H��҅��
Y�4�,�w^���2�O��Z~����^cet4K�\�Fm�)��������H"�6+�w��c��B�3�t,|����^�'�m���	�Nŭ���	�����㈪�d�$�rp�~m2U{ȓ�^Џs<�3��g��
�BB�C���tc���O�U >��17�C���ܣj,�v�ko�@�k�('\"���U�xE������p*�+�Du�E�:":��nf���_a��?�wTl��g�������AP�#�J�v��H���p�U�����@p��,@�/$%k��>�\O��rM@M\Оg=AٜƱT�s� �j�w|�
����/���ǤQ@{P����[�n�?�*�����U���Y�D�;�YH�ԶshA2w3����F�v7�U��p��T\�o5/��Ywb_�\'�fg��c�+뜺f-Q��\tE_���"�p0�� �]�:�$/�����"9rL�a����5����9�ȁ7�2���i��ħ�tҼz+[�f�����U������].��h��d�^,�r����lҺC�P�ʳB-�S��!�֎a�1��wȶ�ZO-N20�*��/��P�`*J�oڎM��j�˲q�.����Nb$�>?x�m�H_���ߟ�K����`L"��]Ȕ3��~�vO}�����]y�������зO���L��=�	lz��п�$�ۡD�h�>����T�G�˲Һ#9�\��C��6��mP��a�Ox8ΰᱧe��e��Y�<�>�ZL�*<l�܊!��1x9����%IJ�5�O�uaZ�p%�%�ɳRiY�Y@�P�G����*���,i��ە60��zY��,�7���ݶ"D#�+��D�Gm��C����C���3XJ_J$i}T�l�� (җT�Α�������[i��ӑ�'V���}�軣��R��b�u`��Q}_��^M.��\b��ŋ�d	S{�A�)�-�&���ڋ|O�5����X>�QZ>���H��C"��P/BLP�YiӁ�k,���>4`?��"w��ϋ	V³L,f�y;��e�y	�E�U�v%|x�X�%�a�o�܎����CB���� b�F�6zj)��+�oIl`\A���-������ռ��=��9�Ӯ~*!*R��9��\�)h��-q�gз'Ԟ��]�]��{�g�����8t�����4���K�1��Gg�=]�_(�u��bRh���d�+�~�sgH4��U�ڛ��hg]���8�h���##-c�̩�'8���6�5R���A^�L�
�q�eҨ�q0�Ek ���"ݡK,o�|�����W<�X�4��G9$����Q�N��O^d�|��T]qVgEW��JRXP\PX����p��������K�ɵ�ڐ��7�Gb����`5ԡ��ə�/cO�35Ł���!���}L����x�啳��;88i�4n���K�/���,L�W������l�LT�1��x�`��rW��фa�:v�	s��qR�����]����'ɘĖ���\&0�a��k�ȳC45�G8��_��žM��Pw>���#΄�q�f�.�-�ž<�q��s�-��	��ħ�|^rC%�0��W��+B^a�e��叾��!�(б�Na?R�}s�At���Zi�7Z��TM����6:��R�lA���W��r��B�Q�>��?�����,���9=�vo��N��iw�w`~f���R�/�wIZ��)]�aU"��-oy���-s���!{O�=.���m�=�_
�t�N|H��d�:(�5D��~���3�N�t"�^�y�_��_��.��?vK]0s�Ie�cuk��G}��JY�	� ��v�B�mA���2�50��-y�#��圤��0F�ϲ	��i5j�<4�dp1}��h�K�w|dU���UpE����?%n��X��nAYMan�y��Я�5+�^�e8?�Z��(���?`#���d�f��ŵ�9>e���V:M;H��	�,|C���&e�'[�*��e�x��9v�@Jh�d��'�>]`a�L��l%�iڔ�xY���ߦ�\�ٙ��8_9�x��]���YeJ�t����G|�z��O�ߍn���)�A�X�g/�?�;���R�]ޘ�$�岞�9���}�����x��y��T��S�����f�9�@/3&�ڴ��ɥv���o0Y\@�ߡ�ظm����9����d�^}$(���Di�,;9@���ڔ��lib�z9����ɡf��et
k"�1G�B�#ҥ����nSZ6:�W4@�wJt�{\	�3//��]�n��J�_J�jg�;'�uoj���>!8 �,�(��F�@ױ_U��G�]��%Ӕz��P�7�.O�|If�����>�=�Fx_iwi��.]�hZ����f�u���j���=xZi)��"I�WY�=�ۄm�G�6�$m���٨�
��X2����o�ه� ����ƑO��Mۺ�P��R�A�sx��u%�_f�v�P��C�}8j%J�n��7���*�ئ/��7Ә'�Cԭ��L�"��L������t߮l��9ZÂn��� *�� �}"����:�W)�=�!Te^��C���^`�F�������Xq���#xK��2������H��gX~�"���ARE���8ڗH��AKm�W"#�7_��+f�4;.���oqa�`��khT{��L�:�B���{_���,r�ҡ�����-�������ќ��?K��F�O���">5Z�n�w��X�Q����Ei�mG6?�j�I�7�/��9����N4�b����U���5��H��l��vmM��1����-�MUY�9M
��H�"U�Fi�
QT"E�*ڊ�VEE>��(��B)�I��c�3���8��s�QGG�
�Ћ�\�@Qha���4�Ji��k-������`��}�e��^k����S�o��N
�6�+d>:����˹�3w�Dc�a$l�|Ϊ��!fTd��<6�&z�Tf��^��q��=x�t�*,�����d�u|]�a �׬Tu}��N��� �k%9�y�'��@RBC�vj�g������2l9(���)E6��n�6Ǧ��(0jޔ���gq#ݰ�6�X:^hNҥ�Cr&��h7��0�h��*�o�r����7����5�5��Eg���C�1�v�lH�4����It2i7���Hc�g����W��#m�q�����d�t��&N���ה4�ԍ¦�'�W�C8�+	�K	o�;�e=��w���da�;?�����F"Cr�1�=ڃ(�Ǹc@t�_�%ɫ���1.1?R���e�7��/��&��f�/0�}�myc�� �;��<a��X;��}��3S��n@S�[x��h��+��F�~��:��D�{g �q����ϰw�����=J�3�3se�z#���~F��/p�Ez���sԚA՟!��� "8z���ެ��$�8~ĭ����>����yř�fE]?�:J+�$��4O�Y��\�8`�k�A*��f�pu$*�	��aU_�����8Xj�D��ݦ�T���|��s��cx�ڵ}��;} _6k�h���QW���;_�p�f~�������g���V�poC �/��B�&�e�JGjf�	:v?�x4���u�	焭I��ج]�A�ۛ�tc*a���{��
��k�Ԝ�A02��*�42�O�>r�'���ld
�f���{��>��955��O$j%�E~�F���W����������=�"�o�j�����DHˋ�'�?Zz�P���#��%'Zu�V�̅�L��P��7�{:��?�&�k���Z�X��w��	�(�2�ʚ�J�ͬ�ay��,��Sο �o8\��B�ϫ��uq���A(�tʸ����~������s�y�Ve�w*c��t�Iu�]bT�����E>���+���E�����#��x�Α@2��=ܧX>�R�~��@�3��Yр��a1�g����� 4����0�����پf�� ����[:Ed��lU�͚hd���śI���͂V�1g��4SGq�EyǺ�S+'�_��R�yχL�"6����o���V|_q�w�6��	�u��⼞K����QC�~DϷ���CI�`~*�@ H{ �2�
i)�;�1�̟���r�Z�k,c���ץ�~�E0�����ex�l�;AT��r����F����Z}4��l����|M��9a��;^^��ʼd��%�S%������X�L�:Ɩ����c��9b�N���|�Dk5��UX����FC��t�ǝ�^󏃹س~ڇ������H?���IYE�ڶ��K���1.�Ő��e��mG�?Z�x�h�V7:�T^y9M�m��ţ��96���j�z��V ��"�FVB{��m�ұ6$��D���]�o3��j$��l<�'�:]l+wV�w[���Hyo�B�/o+s�ﻌ�_A�)$��*�3?����K��3`�1�L��g�$�2{��G���j�>�;����t8@�_�t~'�V�����o��5�3��yS�w���W��!��΀FS|��0�>�ET�~��_�C�8*��G�뤹��F�U�"
�~�O���Ǹ������MWRlrU��ګ>�dw��BT>Ȫ�-�:I����5cm7�D���F*�v ^h�{sM��<U��L�`���cyb�U��D�g�ι�D���c��V@6���˒��T^S9/����l5p5#f�`4�$�R���t��=bqbo�KqS6׼p_���Y�dӿ��W$-�v��;����$�r��x�j#�)9OLߵ����ڕ�.S��2�+G*y��Sv]�;�1�'�
�2^�Z���5�2�r�ꦅ�5�,��GrD�`:��*0{���H;�:ߐ!�nU�-�G+i�7�#��]5^Z��`���E��UG��\/�����~�K��}!u��$l�[ic�����ǡ�w��+�Nz�k������6f(�I��Y& �o�t� N���=?�	���E��X�ys�n�P'�a2H�qñnV@��W���g�,A���{�Y�0��){J�aW1`�{H�D��6���|F����lږ<�Hð�+&,ד_�����Z;榿�~5.30�����&�ޙl{t�@���b��8�ٝlK@����]�8V��Սp`�(?e��_<�xy�1= �ӎ�E��k���Rg��/��x��/t�Wv+�C�C��Ʒ�6'�n��)<�&l��V�o��.f.TOS�����+v0�Z��C/@�N2n��W^���\�qQ|��'ےmg_^ղi��LI�^�h* �( �(��DhZw�Z��a�?ϼshO4aS��f�K�h�u������H���=�Q�d�Qv �,2��=F���r���7;,f�M���=�k��K�j�چ��B}�#�(�������]b�Gܳ�i�������P���1-��oaF^�}6�%�犦/U5�Z�"�]Q`�����%���m�s[�^�Ӹ�~A|�1���=�������G[i����������9���Y2A���b��Ez�#�f����|ٜ���B�2��H���oIĊ���b	��&�"c��%���e����r�����������)pZ
�HMm�=v�Q�a���Vy��|7�0+���}@뉍J��R*w���ԙo�o��)�#hx�E�bxϱval=g���Um��Im�?oo�,G�[�̾5&	*p�����'cۥ�<@�����xp�\�l�5�!�Lj k��{�H�(�	���
�ѷ6���}����!=	�i�R�n_|$?$��Ī�k�X�m�h\�|�~U*���ET]͡��^����;�^|�����rOQ�S��{[~l*8ϦlׯN�G�)�ߜ�/?#0Q�U�_zv��el�Z�����ɱ&����_��H�P��1��:#����cbO����y!�W�Lk����tv��H����(�w�����BڦЃO9�F�\�"���	����w�5�r�)q_�m�3����:�؍В���4VN�i+H9-���= /�������F���l��,��bg�o��~�����"��wc�3^��w9�}�E8���|��{O���)��.�46F�Լ����H���<qk��Q�[�����6O?`��J9IS�����}���T�P�K-_�<ƿ?V\�:^B�E�	EZs�S��O�B.�"N�ø�#���T��ƈHn]��#�C�	���QI(?z��v����y��xu�'�)�1/���a'�$���
����-!V��^�ﴫ�g�Q?�s�Gs2�,��<kN|]�j���j9w�&yO�u]��U�ۄv��+YN���6��5�N�v� ,8�O�1Z��c������Μ&i^H5OψF��_�S�`D��Ĳ��o�7�v��c�y��ƟSQ��.p@�C�@oN����w����:USŨZ�v1�h�"��$ϩ<�t�I�5@�����X�L����D����}�����O��3�ui��3��4�e���T��`�����������9�fW����E?F��g:��5��=:יv��L́��j�I�!�9�3SH0u�=|p��tF"�z�P���4*�]�9.�c��I��Z;͖���k�֏�󲴟�·�ʲ�`p����q��E٪�^�v[�AK��?l��~�����bi���6��ke�	���~}�5)��-^�j$�M��:��_ߤl'�d+[���+�NZZz.c"s�[j���㎻6��=q�V�W��`/���Ms;�M��ݫW���]��جٍ�4�$1��ohd���6��a���U0X�Q�?S!vh��uC���]-5>ǯ`Q5x�T��|�
�.�#J��
��xAʊ�  v����h,J�5s��;�8���HB��;�٣��o��O�����D��'�"�=�;U�[�K}gv�^�1IK�8s��u�1MK��6ߘ��%�$�}�x�"U��)������w��
���w����}�>��g��p?�}?�-�����C8����Q֕�)����䙡]�-Xx�N�\
u*���YD�sR ዅ��LQ��É~�����܇0?l�Y�H�13˘f�u@��ŧ1�8���駱�4��9i�C+�1�m�]�8�M?QdD ���jA�'�q�VM%��<��P���;��wa��b]O4�c���妕���Q�ST�H��wS_�����븕��dR�n��a�ôr`"���&0��}�9�@��Ԛ�4�)۵{�ӌ�tㆬ@�q�l}V���$mpS�,�j�HTe�8�ԓ��Ư�|��9c��9��w!������-fY�Q��I��S��:�D��k�����V|�����_u�e�z�Pl�Ҡ��^�q<�1�m����d��=�ct������n��W�´WW�Lo_��JUk�O�S����$w��S=t��I�*�YR����)ų��y��p�qw�x��ob�_�&Ɵ��m�������:.:�w�gqw��h[:�բ֦���i��yñ.ȫ��+o�iԅ�x�,+jr�ht`BFZ��o^xC �hԅ1��2��$�v�Z�kh�/����n�.b������T&���V�*���}.0?T��i�]�o����K[���A!�J��8��$��?�N'����?�������󅸇S����W�V?�k�P�u���L���?�:.��?p@�N�1ŃL�!�l��>��y��w��c��H�lQ��1���wE�OeAd�~��A!m��E+!$����G};��H�B�d�>͝�A�-T�����7�a}���k��~*n0������׽�@U�������+�����a"|
�(�m���ϵ���T%�PY��h�hnM�z���&�n�5Uj�W�s�I��)�:��!�N��:F�H9�Y��q�π�^�K�@p�����j/����ic|�0 �&X��Q��w�2Arl���ꇄ� �R�r�F�$*������eҌI{���P�����gΒK�R��P��J��g�}+a �Ÿ#�C?#��-G��=��!�Y�8;W�u �)��i�����PSWe��Q���騐B���r�D�f}��<�����n��E�3��k��g+��<Az��4?�}�O[����������~H�u�@eE"`��^e���H�Kdx������Oݴ�Gg��n�_�1�N[:r׫+� �2\q��7�&�s�M]�^'Y����
}�ϔ�&H�/���;SRx�׀Y�M$�G�}��B�'{S,�	(e�9Ul�Ӽ�(�y3�rh����Pp`�u9� �����}PG�+F�����`�u0��[SY<��'~!A���P	:�.�U�N�);��E�s�hw\��K���,�q�)$�҉�?��wB����"�<k����C"sE���y�XirG��e�]�p��<�6��]>B�6D�y����٣�s/��ϒ��G_�a/���\G���CS�,8CY2�O§7'GT _��^�ɦѻ��4�H��^�S���3�F���g�Y�$��n���V� ��sZ	�e�T����|�꿍7b^c�.���hv�Ԍؚ��{M%v���~(̣�GC��m�2��3�_��B@��>#�+Z9�<�7m�'�g�^�TNڰ�仱��{�u��PI�5ڔ�Z홌H�����5�`-� n�~Ե���asw���{rDzE��z�W�`�:�,�+j��7/�|#����K�}�f[���J�>E�4x)L~�'�ci���$7�_I�� #f�5��f*[C�*4+ܮ=���a�Dኳ9l�ޢ��]��^���˷�j�T�u"��]�I��ꐲB�����*�+ĥ9�Dx%DbN���?p"�h�B?�9$��m���\e�ԊS�I��𦼔�u���=:lM�����l;Ґ�M�}��͕���_�-BÚ�#ln�=XL�o��H�ٮ��n���_� %�!���j�@�{�E�]S���w�S����6����N��m��8�����PuW�W��y5�]-��k�w�9�P��w�m�oS�ޑ���%�����P���y�iڐy������n��wO4�R�6��@�����3�\DRT��9��șm��W{��j@7��pK�Z{QUe���ؗ@n�9W�#�WU��ǵ�'Z�*�i��9o����;��U=��.�h���n��)�h�\Ѫ����SE:4'�X�0sh��\�4;��h�ꇯƑ�d:eZy;�D��h��0�!\6j�r�w��WD��NX�̋he�(�*\%T�;�MQ�	��(�� �-~�y�:Ҁ,/_F��3S\@��VT?g㪅K�����F������M=,�Z�+��FU�ʱ�j-�-�H�Q$���REI���E)��dL���\#I]_�'~�('�Q@���*�<��+�����l�mE��bN�n�8�� �����0?��*���|�#¨���Խcq�2�m��3��p���nA*W4��r�S2AD�H����t�4M��l`��կ��gN��$���J���{S�Қ��Fx�V� ��(��|�z���޸v�+�Cـv�$��k��9� _L�YCe�C���u��<����ՇF)mۏ���+}Ǚ���c���P^���ɓ��������fos'q^9h�6�h�o����d�6G�]\d��mK�.%ɋ��3��)�{��+�Y#�����A2�C��}m��`\P�m�X��q9\��q##��W{�p������ެc;	�yu�`�М*�'��}pE����l���'��/K9w#�.��L'������aj��U�3f:쟵��;h�D�^�ߗ��j`��,�A`X�8B�i���/�}c�;��4zb�p*`E&m���N\{�s$�  w����#Z��N�;o�(�I����0)w�v��M+��Z,��%���F|D�Y�0�JE�T�4.TΕ�R�����һq6<~I�u�z��+x��	c�=�qF�B�Z����"?�:O�}z$)�ԫ�@_]�{��f���C��Au�|Ǥ2g��k���l6��6?|�Os�����R�?6M`����iF\H��T�	<Z��Fڴ&�T��H3n��V5i��j�x�Rؿ��h�i�T�y�Wt����&���1i��h_��;����:��!��m@Aqɖ+U��7]ji1���x��0�-:�uQh�?�����x�}')���\�S��Z�_u�-y�"��8�,���D��,��i�]$���5�_}�����&'�o�t��$*&+�X�}FQ�Gz�R�P�0R����T�f��)����K5j*�C�A�d��|����g��u�f�4w��Y�]L'o;ُ��U�\��	�ف\�# �Ւ7�;4<,o�����1,o����
�@�<�y6���89A��w�0 m��%���`���kډ�e�JM\*¡+#��;�t�@�5�S��/�$�CW^R.�&� 5�>���=��%JY�v-!n+��)W��B�Q�`,qN�Il>��z?�	�m��l����}fm��GEM�#���Q��}�$�8�쪣N3b$�/�'��ح)=�B��7
��
��RU�htx�&��)�"U�����^�[M�xS���R���#��J���i^�s�."Z�6�?�4;��<����s6���4k=hJ4�IzB�*��U"��V#�`s#�F[X�4���uFU?�_J����� ÿ(H�D��Sf�6�9�a�r�����#��ia��!º�'�iY(������.�����5Vc��b��7�%����8�3{|]e��*'2�|��N���:��`�$ꄹ1L;�^�c�X�H7�&^����j74���`��3A��̇FA���=�ߝa�Y��(Ɛz�1��^�5�3׮Ғc�l�H�Z3�f��f�2��V�m��7��o���Ƒ�o��cJ� Z�����w*`�T�?�q���/�^��c�A�ߙ�ڭ����S��@�hH2��p�m0�J��W#z;�ՙ�1+s��
ه���E���)���i~Q�Px��+E+%IIԒ��Ü�����ȳ��D]dQ�`�0&�����R)��&S��ڬ (�34Lk�+���ک���c�c�1硫��������̔ qڬD�Bsx]"�9��w*#�5�K���K����h^㗁�2\u����n�
@6�4\���,*�7ܲf���]�/�������_�X$��<_���"u	`J�~qQ÷	�23p�b��S}d��1�]B��Ksf����6=�������w�����*[�
}�a�H��F,��2�a�U^ti����R\G����X`ܛ8�!,3sR��'��F����/�`cF��M��9P/�O�J��D�� ���NN��lbz����ɱ��Z����:��C��&�s*���c�8}�>Y�f��	QE��p������ť@42�tV
�hW�q-ď���68?亷7Kx��+�ո՗��v*3���L�Sg�-uf�s�Ίd!eo�>�-&M�n�����T+���&�c��ZM̀��qx�DV�V_�����˜��`� �����Q}d l��t�*JR�Ҝ�t"|q��d^(ʽ����=gP_�g�j�@bA�l�n�v��gT�c�y!upA�u=��J�-�q^���Qh��#ј�Wŭ�(S.o�*I�&�F]*�{|]c��P�DY��UQ�`;U�hBe�jh�+����A!�a���YD�_�J�oH]4�&$�|�u��?<�a���Ҿ��q�N���g�.FWpo/�N]}條��ya�x=�^�;VsfK�C�2��	��q��ͩѿG��=��/��+0g������O���H ��~�+�O<;}���J!D`Jg���)��t�������`|�.t�O�	����<�� ��a����)u7�+�P-��憾<��O�܌u���~6Yx\u��E���N����j���5�7�0�+�*~�����,�+�vJoi�;�V�a���e�{Zxg�q[���*��A�?���Q�F�(������\�"�
�������Z��������r�֘>D��Rc��3�81�$PW1����O�#&��1�V��^R�b��Y� �`����Ȋ��}��Y���*Q�>_�F�g���
�FHr���W�9P�/:�����:��-_ר��M���;�c�2.2�5
�g�u�j��	˽��{w+IG��.��YP��n^��M�9�Ms�m�YD��>Hc�����q!�45t���䱒�d��&i<�cM���u��Yũ�����YZ��o��;x �1飩|��m1
=�8�� ���޶�d�1������tByr��p�����7I�Nl�,�1[�Hu����R8_���u����� U�O��a�+L�C�\��
|��'����MBl�H| L\ZF=+���������7�0[�]VK|��w	�4���v�!��R�>k�^8^/�������C�6����z��$x�)�S���c����K}��M]�?����c��\(����ϓUݯ��P�Y	����I���2E谄�M���i�o���<����ȊB!9^�v�����.���T6K����{���m*N�/�%��k�8����~���s��������ll��j��X� ��g�XN��=+��X9i�H��>�4R%橵��R���q�-���$m@�2�2�J�s���(�!���^�m�SS���u�� B�H�K���0�-쑾/`�+AZ��<�����ȭ��h�c] e��aw������@�΃�Wߕ��1CR/D0uBE���ŻyK5+��_��e��<�s`�7T�����e��C���[�I�@
��.U%mU�
��*�%]�>Y�4�~I߹��z�?�ܺJ���@���2]�l�U�ج�yĴ'��D��^F$m=U�/�oO�o���+�=qzB���I!�f��"�V#��=m$���+�	Nm�9̎�������X��Fs'=	�l�A�7�7A���̵	���26�{���1�B����B�e���B��;��.Wa�[�����{N5�1����3^e����ن,-��x^��k��ޕ�(~�b^�G��q�Hp��:>^#Yq<�ũ������OV�]{\u�X~�:�����v��-��ʮs���@?��S�u��J$�m�:�z���O����?��B|YP4����ގ�/�>�d^E�cw�;���;���������tE��F�����	����KWn��j�[���m?�F����~C��3�y�3g�SW����s�|�c��7�ַ��Ch%��)MX��d�$�zq�$����(�?�[HR>6ʴy��h�,���6o���1׌�zD�w��A��;����}b�8B4*	�~����1���dxd����ڗ�'�0��^��V/*�$���L���7���Z>f���Ws�\>�3<����P�hJ�U�1I���N�z�M�����s��*;t���� �����snm_���=����ŕ���R�:G/�h6�ި�:�Z�����Xm>��ӫpN17��ݾ� ������xh2}�u�s��#��߾�ֈo���������I|��>ߺŷm�M�K~*�9ķV�-E|�k��9X�a�A����H��sxx�(V�$�;�v���K�_�� ����TD,���-j�3ȸw���"r�r9����\D�嵕9�������9U�E�=����{�bM���~�j�� ,b�C�o���!��$�ݴd�ᆷ�1QB�2/:���#XD�H��W����N�E�&��BhxXc��!�b�����E��=AT��%��4�y�y寏�˃���ҜT�3*(^��wH�N<�'��*�wo3_e����=�|m��\�Nd5��,I=��D���"����������L��'9Y�?X�-�!,����>�Zp�u��������B��+��<�+�N�k_���S1��b�ϋ�b�_�ǿ���e��9��aӖ�8/�+���,4�ER�@�C?W���K�O���ѽm�n��??�� F����lZ�������?��x���ֈ��~�#kx�w�xK�+!�i���m�g]�ڳ�Y{���n��q��Ǹ>���<6??�s�7��x,F���XJ���kj~j�S�tT
��3�J��l�0�YB����^S��g����l�6+&G Bh���`
WT�hf� �b��1@~����he���$�!�Z����H�-8��V��+�+ne��jE��H]�'C����?F9a&c	�|_�0�Q����P��"������'���@o�J���N��U	���I�'�!�:&���A/ʹ�]vՏ+��-��=���gl�FcqI�{hR��]�M��|a��y;p��bW��HVw���BUk�8@�sS��>uX�_�"@��ɳ$i��nk8�i�2�5w���|�OU=lܙ�,�9��N�~���F�?�M�k3C��K����>I^F�O���x�Aj�-��7�n�ʡ��|v�4*,5q;6M�1��B���q�XaQ8��;S��NE�@V�����r��7���s�2}�I��~z�749N��8�Ӱ��rH8:�*>5������K@�I/�V��8騠�1�<zs4�6���`�s�&ӱ�;���O���6�-�������$�ue�e��0O�SBo�+�J���?zu�Ԩ�?sd��	M!tJ����T�߰$>d"��X�!ņŞ��X��۟M�6�ۤ�n�ʺͽ`E,HWH����i�Eف�;����`Ħ�Y��q�7�՜j���������Q���N�z��h�|E��d��>W�.P��\��}�!�-���1�	�r��hRq꒩�Nb��v��R�;�ÎZ{�~L��w2x2\u��U�|�F]���a��""�	��8����S���>�%�}�G��CO�*}�3T�G1�H�o�ұ�c�P��	~�@x9�x��(>^�X<g��8$��KM�Օ���Uj@͏�c���|��	�J�X�g����/]�]�W\S|���_�eEt� ���Ug��lT�e��c�u��b��������|���~���|�b]:��^�=��e�@�g	��l�������|[�F �ck!q�~Y�9AG/i���
�Dz�y/��X�sr�v���̷�83���I�	��V�ǗY���#*B��&G�-���/6~Wޓp�d�e��k~�{���F]u��tʆ��"i�`��;;�\ �<�/�T��z�hݿ5���6�Fʲ��%�'ct�IL�{DLhhP(��n��ܙ�d��L���t��s��	_%��Y�]��m����O&����y�^�Pp�����IϬ�FϿ���8�)�"����'����=��k��n���6�lG�Z�0��1�Ѽ���a�D���8��$��e8��k������W��w��W]��[B�͙�̓���e$�=)d��RFx@��
m���Ks���i��&5y��6���(Js�+�<����x;���X7���Xđgp6���tg�s�A#��42ٙyQ�X�w�r^���ӈ�ʊ)6�mG
OW�3-kF�P�z�!�8��K���D�J{�7{���	�̽+���@T�������;|M��͌fj*����z��N^�ŭ	l�޲V5u5��U�����+�x�̞�9sl�I���U�D�"\ʙ�I��b�(�s�rY4	Oy�_0;�9���؅$!�N3N�9fi$}�/?c��vc=���s�rl򖫌����W�i����~�HO��rv���;,�E����+v��U�`���ʇ��'���Tw��{Z�G\u��p~��d�v�q�Z{�#p���9��<F"l�p����)��j��=��3f�b��b!�c�7IT[��|�Z��PK�@E=N�1}���cg��%�� Uk_˿�}��.�p�q���a\uɄ����`�F^~?ًӨ��jO?�i�C�x4p�� ��hKh�@890��c���@�|A3�V�GX2;����2y�-`��$3�(̍��Z�̿�zX0�U<a�-�e�-�xB�T�Y��h�����g��?�eR�P����3��m��'��c2��ڒ�AD�`�����k�v(�Js� 4�hV���\�4>�.�˝���;!�i"�#IJ�O�o�0?��V�$���|OS����ϖ�@y�,<�)��3P����ʝ�$�'��=C���m��Q�:��y�z\������
�u/�y�UX������W�� �9;N��ۺ�2e��H���V`v���˳��@\X("��絕;ό#��)��m$p�+w���3�N�m] �	��F�1^h]g�0��mSW^e�ۙ�����۶5��Q��4n�d�#Ld����p�޸B�	������kp�)�~c�!j�������}�&T��7K{ �w�'�Y��8� �����|�<�^$Z��E��0#з¤��i� V��w�F�ڙIjm��A0T��J�8��3��V��o�3;�����v��V�4�����ߥ�v�A�;0�I��ی��zG�hOO�і��Ω���v&��^��E�z��'��-�:_�=���=�M[芾�z����6�z!��9�,����C�<���)�	�j�׬�)u����7�B�����X�p^gT�>�����H���'��>��K��^�?E��������rOh�}����y�B��B�J�3Xy��c���;��1�>���l����i��L��L��?�Z��w�Ch(]��7�u�C��_\���x��ȴ���4W]�y~Jh�Co���C\��-6����/0����-v:K��3 g��3=�lK�����٢�Q��2����97��'�G|�	'g<X):�h!<	�&`�o�����2������w< M�����R���A�r';��pt�v����F�V.��R|��A�����MV��,�|y�{�S�,�Lq�/��8I��r�&���r�ۗ9�eX����Q�Ĺ�-HǺ�e���Y�D?����M	�>K����Gȕ�� ��k�P���� 
��X��1;E�s�L���=eu��vr��|5���VM�_�9�e�gZ�.Ƣ4�m�X�ny��r|�N���]j,J��ȡQ�3�i�������N�Fj_��SE0'+M�����B�]����� ��4�1
*V�,�
"B�C�T�a�}�F����(!t�l�}Y�����v!d	�$d|R���n/�MK��>�J��t��FA�}Q�Ii����0�l��C�v�����J�rH�X/vR!tJv�N��RRuاu^M��&������*�6O�����5��c2I��]!�1m=#���V�#o�n��ˑۣM��K��Fȶ�0�^G�e6��������f�3��8��NNU�-�5��̬SŻ]�#�JB�
��i"�|H��~�-���}+"Zv�8н��9����l�n�h�Ҷ��^t�k���rK'FF�(�r�8l������klS�.��-%�"M�-n�wM�LS/������1n�.����`-��:�=Vڳ�EpRc�4��a�q�|Pi�iO���j���v��d��I�����m�oke}�@}נ���﷨���
8��*��ҪG��"�x�{�ە����ɢ�2�|���_8�_�-2��a���l����o�Sij>�`����4e P���dĦ8jm��V�TJ9]�p���!O3��eO�t��5��n�9uB8�f���d�+��J��e�?��T �p�ƫ���$��ʘ��9`/���[���.f�2�X�_���X�"�ޓ��tW�\��6�9��!�2[�o,s�`�H4��I�P�ݘs�����Q��pXh-�CTOpbp�x��o
�'���Gզ�j:mR��k�!�B��:W�Ď �y5��^��9����0����c�92�÷�K�
E�U��ӱy��,tov��S�f˛�]@=%t�4��]�g0���b?�J"��F�x���*�a���Ǖ�ۨ��_Ɠ���=��Ā��h��w�k#Q~->�Y3Ns�
���z�9��_|��4��7)�u�%>����4��e���zS�m"��ș��K�
����HQ��#׿���\�S��E#�f��T��M;Lf��Xs��� 0!8C�;́����G��0��*=�h�cW\{�MK���|HA�l�-!n9be9fM�����m�$#0��`2T�"$��'Yq7�����hy��o4�鴶/�����{-� g�����Ms��t��9��QM��~f�?���<�Wܭ�ֿM���.��7���1V3���/��_�����-��3��Tæ����d����>2�
�R}�d�cTp�RuWŝ������4:��+��\��G�����_�����������z�96�H&�ZI]�Po����C|�&���ʼ��|�K�pu�����#���y5�$�ɻ(K��q!m�;"�N�^2غ��x��F~:ߑ4�Im2�)9��3�ݟ�����[��������fn���)����Oge�0�|�[?�+�`�_�u�S8j�X}|��Nˬ��V&�C9�VX��I gar<9�A��S]� ����^��/Y�}4H;�&튠a^�1���<\�w]�>�a��p��f�,Ơ }����9M9���f>>�xcj�D	��NI���U�AL��;�Oo(;���U_�{.)������j1�����ug0=Xwl��o�T���ݸ�l�S�6�͵i��@�7m[�Z�0���m�5xc����I�j5o�C50��G�a\=ʞ'5UǣD��B�G�ղ�O������:�{���NC�w��\F=rxpF4�%�"C����u�D}]c��ja+��Q"1�3^���������������_��3Cm�(�t#�����>3�v�V*��h��*��(����zMf�O��Y�@*F�_��%�:��B51/T��)��}fZu�ފD�S��25	�L�^���lcyo����JZ�����3�q�R>D�]u0�W9��\��K�Q�{>��%�v\�&�*�:�Հ�w�Pk_òP�O"�*v�]�^
�����Y������X�c��8��Ȋ�r�L�n���>���M�/{#Qw�vn0(�Ò�U��i���b۳���UW	�L�ji$��E֦��
���5��}��C0x�i	�y[��Cn�~�3�g^��k�	�^�۸}����?f��C]�A�.�����y��}dg"�2��Xx7?�=���>[���#���'����7'�sj���d��C�����Т�&�jNs��_���p�;��:Ǥ����GmBK�������HRBLJ}�����.h.<��7a���N�DŦ�������:+�
�h^0	��3��``����n�<`󙊻����B� }_�Y��6�s3�]��J��ȶ�~�CNoC
��s0q���az��"����K������ד�np�>�������q�èH1nK%�I�4�Cg���*ˇ:l�0��oK�Z�Ç��w�N�ST�+�_ݻ+���=i�w3��9CjE:T6W�\-�^=l��������Ggd���Վ�h�'!�~D�U�HY�Mc�;��Y8�J�l*LLab�%"1�.}V���^v��x�9���D�p�^��sPȲ�'Hz�,��^�+�C�GO��!���a\���Z�!c7���qC*פ�q`S�I�������^�����;��i/UzOF�a�<���������;��Ţe��z�P���u9S�i�J�!�E��_S�)h�}�[�>���������6�g2����2=��G�yې�W�KY�n�.��vh�f���������*'0���t����ݘ���.���G6�88�VY��Z���5�õ$��;L��郔�n�b��`����C�˜y��m���8�4�gޑ7L]���n�-��4���K�ݪ��I�#ԕǬ���f�\����S�e��]�z�+�:�0��J�����yloӈ�J��Q_Hѭ߼��@׹̒e̒X,��aIi!��J��{dt&��'t[À��R���Z�G=��(��H b�����{�7�&��|^|�2ӣ��T���rx�lb�Jz-t��=�띜�5��t�^<k�h|�����p����b�HZ�zfm�4)�=�-�Q�����pݠ>%�e��P"%����y�"J�n�߶�<��^6MQ��C�2�붋�5�bsZ�׷ M�t&MӢw����k�E[;���� ћ�{����S��A�7�_�*Yߧ�˲���J>�Sb�,1%�A[����j�X3���j��S�\.	�鷧������Q��c�x��,�}C��~�������U�(� ����t*Z�\)SͲBT�n�5�����O���ɂS8u�(�H��K���mm5�>���/��w�>����y:I<��ڻ���>O�H�D�t\Â��S��@1!%Q��3���T��%nD�_�)�,�䵷��}J�������ӧ��ewG��k�Q�ӧ\�U�.k�L�S�l���(2Er����`Z�B�K���|��Dﲖ��>E� *�JF���>%~kU�u��}�,��  Z4��O�Y��X��}J\h5��6@���U{�Z�<	F�7?�x�#�b�L�#�[��V��Sҝj��n���w���w��

.g�P���QġGPW�7��|q�w�� � ���/T�c��B�G�����	�ڻ�[��xZ$�ޣ�u;Z?��h�����4��c1�0�GGF�x��j�~,���������]>N����q�:]<=���&����������';������U�K��F��}\�W��im���Ծ�;�l�˭4Zz�s͈pit�΍U�u�j�v�)�e�}J(��+V��>%���,�O��vp�w}��:�� �yշ$>~�c�D����n�4Ρ�#|:�i�xr4S��V?��9to�4�����(��g���VwY���}J�������Rm�2�w���3��W�>��U0�6��M���>Y��4���b�4/���t�C�2�\@�U����K㼚�������c�B���"�UF�Q։�_�=�1O�*��'����güi��e>��j���/ϷiC��L����H������VC4V�z�xd�I�i��ǒ"�G��l����.�OO�CAf�Ǻ6��T��@j.|4נ����>��}�`<���bYbm�a�����[�X�<z�^S�<�_M��WCg�}�$Ŀ�2!�}�ӳV�f�M���#�9t�a՘m=J�_�����0ы����s>�$��A�_A�f�'���#�xZ��$5�,��m|��:�ʑ�$�˺�mH�}���$�iJPx�i|Y�d�qހ����V>K]}<%XN�x�11r(�&Q"PI
��#�׻�Io�}٣n��zd��KU�S�͔�3fB�uS_^Df��g�U�h}O�2n��@Ks�.�/n���s�E~������f�g��-�a�F��Z��k���F#e��鋰Wu.f�fFOE�<3�����]���Ɍ}�;���ہ�iXx��Ieo���|޷B��2m���o��:����h2B%b�B~�g#K]�����P���n5����㈚U�ȟ�
������TߗJ��S�[�D�i��`�k�JN+�O~���է8�ӊ�����6���:�h,�i�Eu�o5tG���&��"5p����6SL�ou�d�.\�i"�|���;�N�;������(��ز�7���9�o.������(+|p������߳Vߙ6O/u�r�7��̙Ƭ��f�}�����  mғ���h6�ZZ�\1h��5]<n��K	���B�g����y��"y��R��1J/�e0�c=���W�Ӽ�Y��zS�KՏG����#{��Fثz�k��U�|�M}�������3�c��Ҹ��ʤG4�j����x�����yr�/�h����"���sq��U���&�|��"�,cZ�~��V؍3���LE�^"Sc�:KCu=��O�D�n@�o|��7�:羯R��j��5�j|���ŵB��c��Tu�v����h����XA3�8��~l&%��Y�\�����V�j�����&]�Q���?���3��푂hD�@݋<�v�z�)iޗ�=���hC%�o2��x���u���jm�X��a��þHTo'y�`�q��kH���L�#$���\w��J���M�j����{������������v�H�{\ȋ���|T\�]�3Y��e����li(�7",B��g��~?%���"���i57�Z�$���.�>d��s&xԀΧ���~�z��DN�P�����d��XI"��߲��.�/I����(�Ǐ��#�71�!���P`�co�>� ;�`R&2�a|�ẰSP����i�Dw���=��]�\_#)QĠ�!Ơ�dEP8�-��$�	�n��QH@+�yϰpY�(�g����龉�'���!;�4A�����i�!h1C�ȍ���;����Q��P�jWyZ$����C��K�[R^��ӜCd���'�t0Q��µ'p@oZ1:�|r4�f[r��s��
9� l�Qq��<�����H��e[�k&g�({�g�@E΢r��*ճ�pWG/��a��M���P�HC�Y��	�dt(���Ƴ-!�5�d��9��Pۭ��d�MlX2����o��qawju��kJ�����z}}h@5\{|_\���
_}���r2�ՕSQ�<׀x��&Uϲ˻?T����i�' 穀q�� =8��OѾ�A������t�8E�ؽS]�*/dx��~�����H�U�oZY�̠��$!�ypi4�`]�o4��+�Y�9ʊ[�w�:���[��MF���x�X� �=�az�#�O@|A��x�N���;���f��+K���z� E^�Y��^��bv�A�Ӑ1",`�Zt�j��QW2i ����܉�tǯ`�?��k��;��;�iG��\��C�����FA��Ϯ:��@5����"]�/�D���$T�o����܂�c�|��$�驽��<N�Y�z⹙4;�Yn�
���p�_.BPP��������F'�)ԇ��@}�i3o��zdn��,�+�7��t�F-��K�c�E·֌~�q�5=�IG�4��.a7��hq����������H��&���=˙����,�>� �.��4���qw&V53S'�����L'���f��?S�y��-�� ��Q�e�cy^~WH,�R9��7�]X	��)'RÉ�n�oʉ�dS��ޗ�9��-G�'��	�އ�E|�#������`�����:���٤$���}�+ͶE��Ӝ������� a+�ϋ��Nѷ�T�M��P1_4�=�bv��N]��٘�óݐ�@]��vl����E]#��K�)�B=�F8����6X@o'���p�F��I]�h�"aD���l����>���­9��5�(��'/au�����{���)Q�+��H,��ʓ��}��ǑL�"����B#sD�sCW7\L�2��r��ʰi�V�Q�@��\i��(X�ղ���&�̔�V'���˩f����6z�kWt�xL��3����~)ϋ�.���e�+Z�.Ǖ���C2^�A�f��X�S0����N��qi�����4PW1�x���9��V��{ ɿ��޿�$
���4��{1�%���X��ކ�U��ǌ��]`��{?�{��Fc�1?�3�z���i���;CE�3���^�g[���i|̛<="��ubg��9w�h4��>�ܜ��<<F�{*8Q�nڴ��!�\NZ(�x�xI��k3`�_^�sD�|������_B"�[��������d�m���Fy�o��7b�G�E@�4�օO�p��(m�=!�Z����~�+q`£Ns�����!����	�+�'FN�k��LJ\Q�R�<Dr��*��aq���sa�u�s �E�%4��^���T9�i�I��7n�M�$�և%��T��<�ƈ�x[���=~�`�^�qJ�\�WZ��>�ɽ���l���6Z��7��h�hd2�3�v�q�_��g������d ,����Lz�f�B�����9��	O�*�{��c�2�gg�y�g�ˋ#�������&���'���� 1-d�a,O���1���-�_��拤���Ԥ�R���x���G<��Fl_�u���`�<Kô=op,m^�P�ieH��ؤ��.� 7���˽K]=Sa��._]�k�eK�.��S��!�pE����M��,v��(ؔ�&[��:�N����`F�ġ����{ �3�)m����$H�{ʗO[�p7-�����@j����$�>T��4)Y�c���Vt���ڛ[M�⊻мi�X�xW��"�X�~CaN��G����{�9=��/_�8� ���X~����YRwa]�L��A���$^]�љ����o�0��&�C�M��z4��!��bO�gFDwK�s���ރ�5���|�$��x�|ɋÀ���8�*Ήx*�j��~�-���F����l,�!ѓy�Γ
T�p�&�GD���Ĺ�*R��L���!r� �L٨o"i���2u3�^��()����B��pq$�	�g�Ğ��w����](�D+��`~F�F�BJ�����VPU�'0��H��0bAz�IV��n�}�Y�q���#�6�;�d��>��ƒJ�����|J�@�)�~��P9���Ysy�
��JP�&�fc�ffs�|R̦9{�4�im�RPۈN+><*VN��]�ӊ�v*�;a���b�i��VP�Y�������K����d�/'k�1��m�׺�s��/��zzF��0k$���=!�������:_(�����|�5�>+�:�eT��Y��<+_��,�7��	y���|�z�R�V�8ֱ��1�A�,8�C��w���-���J�x�����V�\Fr9o��!��B�99�p=��:>5�֞R}��@-�w󣋿׷��iL�Y�J��`Ӌ��%�W�7eD�~<��턲\� �+j��.�#i�0���"K�e�<�C>��|F'�y!?�~9��ꕻ§�߰����%E!в"�s8X��-�I����lm��%w��Xz��Y�֟�+.����J&J����T'ē��Ȼ���F��4:b.�S.h=�./)� p��ף#����_�W�F@k�9�;!���K~��ǳX���]>�;��q&���h;]zQO41�ߺ�H�h���E�3�=�D�$	�>[��'����|{o�h�b[[���5�H�V_�*[����d�������
}�,r��y�ଘ�l�?�����G�@�6j���z���Ȳ�J��%�+�í�:S��k�	�ZFeDW_�C�����Gx"�N"aFs�^�694�s�lY �2�o��^��tu�:5��k%�9�HS�ꉁ�w�G��m����}�Ioϖ���yU|ƢP>m���Z����i VN�0~� ��κ�����F���m��r>s�U�=�9r�l����'��V��̙i/L6+5�G/L�g�V�7*����?b���yP���p#�Ь�]?�������h3^����@�BG���3�y,G�b|���R?�����3�W����``��3�?��8�R�J�ug��r'	���5s�^��D<Dז����4���4����C2�#���o���Q[2��72�w��K�ef� S�*p���v�����`��ҋ��\��������w���<��w6X`aXdŨ��4լ�Ou�&a�T	1*mm��S��B�g3b�C����m}��+& x����Y�B!����=������~>Jvgg��}���{Ufi!o�)��m�m~6MzO_J�m�-� ��"��L���������B�m�LI��1���Y�e=�Q��e�ui�(�A��
A�VHB�m˰%�H�ܚ�ao� d�S��3fi���Dt��.\�$�9~�D�N��	�m�Y>����M�����;��[���g��|����0�A43|�Eb1;Lx?��>��фM./�%�RX��� ��vճ��S�"B��t���I�^�\j�6�8�~������aT���}���L/�I�&UrƑ.*��.�/,�D��D�Qm�����m�_jId��=�W�Eo���[4�g{G�k�q�q.<�Ș�m�c=�/QΩr��8)����3���c��_���;7�'�8ۯ�������ia�-��e�^�s��ЗB�#������1=��>MG�����������ӎ[K��i�T��Ku��,'M����ӿg��<������zҩ���FA�Y���-5~T���3�K�^�Ctְ�.�a�-H)#���V��I�v)x���Y+��rY�1����M������%+�����;��U<&�!��l��3բ��yf���g�>u+P���\��bd=���\0��ع-�E�t�E��2��Ŭ�Џ�k�i���Xq�|��7�>e�������aDyTL�<v�aQ���=b��%��?�d_/�p���8xi�??~T������r
Qd�)��s�IYů�qh���9�$�#���Ԕ"Y��+�F���C�,����:��ß�\X ^:�C1��PżO.h�x�|���&M
d������+b��2�]ă��a����Kl�\�4���iz6=Q:��b��j���
��	�H_�'�E���8�&��h6<���9	I 7�5.�]#�=�8�-qh�w��5�\���/&�d��|���2p���izs�y"3_��a�����E:-�������dg�����
KxJ����NҸ�}� ��)e/~<T�mI�>�^�;�@`jd�q�Ų�$B������m�lf��� <�D�-���V|,���Eț��l3�˵��D0[Cw������b̟���'q�.19;��}��61!�8M阝(��"��O�y>�T�*�Z����|���ڤ���"�f�?� !/h6Iq�-Q��άy��֧zL����Z$����mW�kG��ĥ�g�u5CJ�ds{�B�&5����^p�M��n��,��^e{�ˢl(K��1y�D��B���C���&?�B(�@N�X乲2�ʐwX�r.��b�~�VD�vt#Y�)[�ӗ�q�B��U �O<r�q�OZ]��׉�r�J�6��)G�����lmZ���s��=ܪ���;� ����j򠴰W��j��8���G��Q��!��.��"��0%y8=�j�]�]��d@�@�����;s�
��7^6�` ^c�v�Wѭ�by�Q�u]�'��S���3f�(����V�����?�1�{�K�]G3[����z�>v2�Wz���?g������jW���U9��^�l9�E��XﭦK�^m�>=��J��!j��N/��s�M���}�=&���ȸ�Y����� 
+k�l7+�v'��YS��6���mMv�J�tE[�����GOl͘$�{�����v-$��W	��|ץ(��dN(�oP.@Ȋ�'�w��q������ȱeH��f�^a7���rb��	|	�Mz]�l�{9�A�#Zm|�e�6��!LS�ڀ���h���X��ӧ����7h��ڴ��\0��>�~�b�|«]�6�l������E^�!�� ��>[�U拴T�++|�$<�}�$?���r���C,�x�ē�ʿA�u�k��tuX'���F�Y�!�����W_cnn�p�c6�{E��oz��ȇ�tW��K��0&�C&pZ`�>ǥ}���+����>�v�3�DiS|z�+���J|�c[���@����>�8�q=zE��¢��`�Z3�$_-�"W�"Dm��0�t!.Q�n-��D"�<�%�x��&�l�#�G�|���t�>��?H� /)�c��
���/��rKI�_�~���@J]��Ms���=�?ݓ�:p{!��^�? �ne�����1ͧ_�r*�Ro`��r���sIx����םC���g��Ssh�7 J�䕪M��~)G��m�V��V[99|�^S *�$�ۊ�x��2�]����x?"��}�[e�����L.2�N�Г/��}���v������z@����L���Jwf�Ds���6��^,GE$C�Qp�ج��jR�/S,����3܋չ��fz��QfR3ɻ]�� 3C�s/��ݜ1��1����{L*���r�_޼+S@��c�r�R �v.���������@
��X;��&�H�Ħ�l�ic4LC!'yoe�ÿ�0�3u`�A ��nx�VT3{U�_��ѿ���$m�ƶ���Ms�Um��׶P.JL�R�䦳&h۸�ۤ��*�/���#�l��O�R��߶b����xk�g p{�b���k �b��-�0�(a�xv��_"�i����wh�_��sx' c���H�G[�E�^)2�fo�C�?Z;I��V�@�4�rR)��Գ��"�!�\��#�/�����p!g�5��bL�O�X�f��V���h�V�L IZ4(�i�}jN�Bd����s�h������$�\���]�d�Z����$y���r�+������_y��O9��:���M	��6�\�}�J����"�y�PW�~����� F���v���zQCju+��exA�?(��H[�d�9������M��l�Q�e<r!SM�ܹw~w'w5�c�T�J���h���;�Lα�����c�Oظ�d���'�򣭒���%Ri�k�l�����S��"�-��ʰ�u}���o_��/$�#k��x��F��Wzuq��j�Ǭ���E���H�Wďj��x��'�PrN{HPKH�*�D�����T�f�2��8���C��[���������j�)��p����9����º�v����`CӉ}R��z=�/�W�#�ItĶ�3�1�� ��r�kt��%�b\fgK����)���/����4��貿���4dm��h\�6ճԮa��IT��vO8��XGCUF�NT(KT|�v����@G�0�*+�WX��kB��V���x���������}9�߯��*�����z�g��dd���C�yu����y�iΫ�V���>��f��H� ��%h��Ċ:�F��h!���O�C.�u�[�Qx4h ����A$�f�����ym��k��T~�El��j��[��J��.�3ބ�?�1���XS�Ӯ��z�B����AϚ����Ⱥ~,�F����)x�ﲽ<��uR7�bѫ�u�g��rikz;|F��:��d�����~����ːvI�ĵ����Qֺ��ܡ��K���~E��/�K185����~�rM�T�� �i�,>������#��rB��ma�g�1���;ƨ�SF�!Œ�jY݉!M#,(v�yF�1��
-�*�w-��X�h>Z�ڕ��kL��h�Db+�T<d<("�&�HJ5E��e�`�A��x%;j����V��a���ʘ�.�u�J����Ԛ[^����E�\ΦTH�W�'E�H�CQ/vȫ���m7��˿���8�����ۨ�df��]�V���_�ƣ-vk�*��zХOA9�p(;h���y��6^��A�[�:�@���6I�u��'�<���+'��^�2�ɨ�ڭ��*��3�>L���
�E�3ͩ��x��e���ɂ��u�4n�'����(Z�j��A�����6R f�M�gc�YPO��Չp=ҡ���؄(D�fkǓ:�V����\��H[�K�a��0�;��{����Q��$���hcOg����es����q/I�(+�֥z����a������-���T���9�
�j��pEk�e���Jb�(�Cd�r�~b��O �f��P!��T��RՉ*9l��j���TK��1�<l�!W��L�uy�_��\��؅Up���x6񑕟�؎���ӈY���`֚!@�@9�P޲���[�^��r&p=΃7pФƨ�j�T�
?�+�!��FK����f�'�(�^E�9�
�}�*���5�K�!���5�Z+/-�r�1�J7�ME�!W�P�)���<`u�[5E�
��?B+���6)c����hu�,��>u_��
�Ƽ�y�k�Yd��:�R>�r�m#�\;�͏U�DX�>ZVFjG�w���ñ�a\R�,t`EX��,Ox�X�#8@��LDo�q��H���ŏ*�~�~��M;�~<�]ƭ�yk�D�[8�?{Z�p�۸�t�����|E��(��D�%Z/Q*`�F��ӕJ�c�(��o���O�?��ǌ�/1��0��$?\jԺI�ꕄ���A����5��g�o���f��k��,	9����G�/��t+R��Jg�#�������PP)v����N翄��}P0��C�SS��۲;�	*�Q�`0&n?�����?\p���AG@�K�Hm��X��:�O�>A.Ϗ_Q:�j��D����2o{��5�k��8.\q���$~6���ӌ�Df��4h�~��K>8$L�)�A�w`
����O�+�K=Y�H�g`��X|�G�����5�؟�Tպl�Q���>U_�}%��2�2Q�N�6QG�K^S�Di�2�i:�H�����cj莈e6:Y1���@�䯩ѯ��:��k�J��{��m�:��k.>�N5��W.�������������qp-��q5^ފYP��lG�q�ȴa�Q��evo����t���<Z�u�:�2'�2�ri3�;��%�/��S47ބ�1��}Y��
��[��o��x3ol��wg�8����36��2G��ӑK�=��s'Y�e�k�w�HXͱ�ͫy�UWrvށ1tn�g����Q0��b��iY&3�On=�	��| 9z^Tf��Bn����ё���$k[�C�g��]"C���!��9�����§�2q�*�e��{��-R˷C��a�"�ts��Bu3�-(����7���ÎDI�D�AOe����=ԇ�C�<�aȳ��a��΀�{��)
��vS�������e`mҥ�!��/ձݟ!
=�pCf������mMQ�ul�i�$�+��/�X|�%&Ϟ�	!j.��W�\R�-^��'��QWsњ���͔1�F?���1 �j���,�t7W�t��� �Ǎc��c�;�!m"�Fm����|V�=��EU��K���$8*{Y��՗�B�7��}�o4�ŉ�l8�>��U������Z}%!�H�c��r�iP�P$�lR^>��p��,��6ӡM�%�js��e"�m���e�5�Ae��!���ﯙ�����-�P�����[��5z=�>���Dnb��2h.��pgi#�`���d�M6�uƪ����0$_��Kɍ�Ĝ5��?�z�y���gق⭴��F���!�#��=�ߡ����W��s^�Y	Ƨ�U�#8����s���:�6�A%k.ġ�ғ6�����M��
�X`1ֱiT�C�-�_�fp����A	��E)�A�吏��F}5G�L���T9'+;oJ�1���)j_����׺(�+�<�u��~��~�}���([<��)�CQ�Q~�����'�ȵ(������\�Iq���L�c3���g��v�3�������$RŽ\1
P\_�>�T�AW ����g�A��=�^�@{
�x�"4��H�֖�T�?��A,��j�հ����~�_��b���ES���W����R?(o�<�G$����Φ���?��)
���Hl}F��"��sLQ�&��5//�7�|�A�q�7L�!�ls��I�8�ǳ[!�$2,5���XX���ѳg�������<m�.����t���1��VT����*8��"~�E�v���n���~b�-�C&nնcE�>�Y��h>/;�@ژϸ{}O�(	iA�����.&49��!�&4a�	��8�U�L̬��$&�ޮ�Ԏ��<��i�����"�E���@Zn�v�>�D#��)je�D0�w����N�}G�WD���-����E������2ף'\����}E��:�kqYU+Q��d�.�I-�@��mAxE&��DD8BN��q��ty�`�U^(�(��mg��z�I%;�6��2� ^0��}����r�2ؔ\�"F��}oA]i+��FQH9��c@�V�anli9��`I w �6�Qh��z9#�����G�H�w6T��\��4�!�W��H\Y?�J��~+�Ȇ�{$m?Q'	WK�!%�`S���-{�W�d$�ϐ�g��+��=��KN]�
�n���pkѵ�r,�!f4�#��t��ؓ6N<ir\��o>�ۢk�3M{dg�E������Nܙ,E�~QNK��ڻ�������h]~���&}`�i��.���E�D�L_$�2 �,ދ����6�ٗL���X��t�����/��l��k+ɗ�<x�YWv��.EI��*��N���fH�/o�tA��@t@���L�m���>�@ �O�h'�4��V�IE�M���ޢ	t����V9��fbJzլc��u�3��>U78��]��,�O��ItE��E����z�U0�yG/u�z�;����[V�YU(b}�u�Gd9���I_��jv����g�=�C�)�RR��|�z��9�9�u���߃�=�C��oy6�ۛ�� �U�S��pW%ڡ�r��&hNGx o^s%}�c' y4��c�f�L��	�{�(e���t���Ȱ�'@��N.�V{݉%C��H����Q�������TY_���O�'D<���W95�38�e�yڐ��lVҐO�ňh@����Q"�T�vf���i��Obl{���
���k�B����S��)<��S�HFEx��M�& |^$�g#�$�M�f���᳐�k�mt���P&�:��\����ō_@��:��q��T�8o� ��q�k>-�X�i7+ba;�_�� B�`�G�8�e�{�D��H]�ʊcr�F45 �D��0@�t�����̛�Wn�b�Fg�/ڇ�����=����Ч<�wlMc��?VB��r�￠��ϴ#rS���(�5T��h��:�ο�M��&��;T}�5/)�k���/��O�rW/�y�x�s 跽ju�͌�E샶L�hk�D�}�)s�q��ς��I��"?��E7��W�j�9A5�fs�^���a�;{��'m����yh�#3����O�I,�����xc3��}f�jd�]ȭ/�~�t�д?��ȩ�q=|����׃��w��k���hC��}���tk���u�q�[����ᎧqoꡚFK��f��#�4c���#����f�n�u���V����֖�$���7�|�'mV��3�m2<J����}$6���6A�63f!�l�B}��k~�6m����'���g�sc��va[�D9qv����#���'�h�-$�Z%.y� ˸��긶s��*kcKML��]ہa�j�8q��G���á��1̄���z3u��׷'",7��c�w�'�<K�U����g���	���T����Z���e�v �U�($7k�пɏ���������$���g�%��Is�X|�z�'��J>��|5=��g�S��H?�E=�(#�u	�'@z}L��j�����*����;*�W�J�~�$���"�soF���ֱ
v()	�[���_޷��8j�%�J~�c��3.���{�߽��["B�*q��g�il{�'ݠ�u��Ѡ>��]�� .�tj!�"2"�Q?�n��<b,�y��LoX?f�dKV��?�ԗ�l� ȧE{7y�� `���j�e$9�.c�1I��b8��{^ H��'����~O�$�ZPr�S�C��I���7Zz3�u��~���5*ߡ���*m�5�N�إ�1Bt%�!�/�Q�#<��/���"�#qv�y��p�%X�r/5���R�g������e�%k��qK7���T5ζ����V�}���abI=i+�[k����[����+x@�G����K��GsN�zYu�C��1�q��a���Z�S����͹[#��[ʉOt�ׇ�9��iKZݙ&��/߳N���L�v\�}�/mE�N�~�M+k3˵�
mfUdB�>ӡx��"V���ܣIR������u�Cw��>I8�$m�#Q��Qi}���.'�5sr���$�^�����G�����nFջ����f�9��h�'�
��.O��hb�d�,�__θ��$�F@8g�9�1Wz|�>�/�G__.��M�F=��rO�ù��}2Ǡ$ǟ�?�y5���Y���]��z�ƒ�x$ׄ��M�z��m�9�}~^�$k��t�C^S�Uf�S窛�����Q���ʑ��>���)���3��W�:�IIt>����ȧ5�h��u�f���[��6Skԗd��ӑWtu;E�ȶ�;#Yf��Vە�z�[��P�1*�>�P�r�^ԯ�ٹ=$�ov���o=Į���X�(��B��f�D�G��G���dH����79�i�%.��Qn[㎌P�xmk���G�p�2g��B�� ��&���3�<��b��@3;�ބ�QL�/�$J7o2K7�k��~%)ҟ��A�h��B&W��f��f�].�S�W��[�[NR�)�]MN���/�A{j��k޼ؖ����h����ne�^�)��[֧͍wD��f|Ã���g&��X��6'���A%S�;9���m����f�¡O0��z�>�G��l� #_����sي�� 0�^�V�)�x���Z�@��ϭ&t�h$�����c{�#���o���.���ʒ���rS<	���Fț��V�ȑM��E��Km��l4��D43DC�yn3��cYTB3m����)��ǾI9�RA�r1�F�W�1�n��8�M��S���@8^&����UB�cOY��8cl�Ce�D^��Q9� ��3$��r��^Aؑgu;��&�Mϓ'�
�y�O@XsMJ�����AR��������� ���Ag�X��,���%���|ql�y��v˲�ȴ|=y�O�����re �L�<�Q{�+DoPd�F7��]CY�	�s�P�����E������D�W;���Q�u�I���+\��:��?#�G���,3�ϊg�O,�6�]���Ԡ�~�!T�A���CJ{s�8���@ȍ>D��@ӊ���7y�9 '5P#Q�>á6;�-\�vs���9�6�יga:�2י�-DJ�U�	�~A��A�g��J-��D�� q�]%r�I�f'��#^�W���tm�vX���z[\����^��ǅj��l�[0�{w3��gL���-��h�G3��3��<��������F&ɱ�[çi���y�4+`��vt�Pa/�L�o�*��C�a���UOҥ�Y�������Ø��[��h�7��I�>2���/y�1��b+]W3�#�5��F����M�;F�UU0�9��u���+����$e��i�n���hN��8����]/,�S�[aqh{�����UB�ahe}�E=jsP�$8�E�##�� �?�ʕ��ޕ����2Uܐ�|�f~Q=�"��Ĺr�c��*��;�A��/8,Ǐ@�*�G7M��o=
���R�*�nd��-5�*\LNᯓ�Xd�W<��x69���'"ԛ�7/�_ډ#��&�ΗZupNpo�ɕܢ�<F��3]��|��Df��ɳi)�Lt��~B�'$�6cC���z��N"���l��O R����}��kԹ�o�=^����U?��m^�]��/��Dk	t�q������3j��l�{A&^��3��RkN�~���iFJ
'/Df�s�aO����r�A�gҐٗ�j�{�`�ܑ�E䠰�S�e~;��H�R)7�����^�\��`)|�N�ƫ�f�B�����{D�!�e�Ejb��x5�Am;ɥ+6���'��#?�$�Wm��C[X:k�h���F�Z���XG!RK������^&Ķ2qܖ3�N���H��:Q��U����]i96{�-�Kຐ���f��[�$�_I�^I>�c9�m�~�c�
�z�PP�����)���(����=���ڡ8����L�P�~)�'������B��7�n�(�;��:��i8"LЏ@g`�V9~�g��0h'�v)��Yt���N!�؉�	0]���l��J?/�㣅�D��m�/1�u��
I��#�?|JǓwa#��D���	�^��ѹ3w����՝�}k�@4 ���p��q�����=��C�]���L� &9�n49��_pW�C0�?��b���'�;ǡ� �������OM��j�!5#Y�3V�K0
���0�"yXi7C5������\�e����6��@K��9{�i�q�.U 6�Eu���y"��<��I�^���)�h�V���]�w� ^��f��˞�2� ��x�F�7*l�׋�����3B�l�4��$_����l��J�"�X�nOz�P1L�+z0���H�K(�4�;0ڔE*,m�OKr	��붴��:�B����aǡ?�Vw���K��V'����>
�	8M� J��Dc�^�Z��Ye\�$O#5`���
�R�m��V���=-��U���y}���b��`����JO��Z�8Fh�ӛc�´��ܬm��fzN>���~<����Zt:v ��������a�lu�0\4آ�C#���L���ss5�9�}+���lQ�Br�T9�ě�0[���c6�#�62���d�4x�h��DQ��,���h�G,�a����y�7f���4B7�����!$�;��b�tQ���>;dr�Pa�����n6��_�#�V�D/Du�tt)�1�gg��~��9���?�>p�؋ӋL�1Y!���&��?>�%IL��K�`�f�9��.=�ΰ߲�S�5^�kVΡ�^�V�XJF�-��($%ת�6�:��3��D�j������z�z��"7�5ַ��Kݶ����0��0cSގ.--*�.E3>�~}~��kziѠ�`� 3��$�D�4�Gx:X2�4�%��tj:�������G�ha����(���e��]:����
�Ø:�Gt�BtM)��?��>��o��ee:\=|<�Ν4���5�����LSf�[�z��pM�:����q����RPwB/x�οy��U��Anڠv�㨩�ݜM7$9�v�ah��Kf����ɽL�4���|)~s�8�V��N��
ԩ�D�S~76�{�vsR�8�i�/������"-\>�n�!b�xc���_4���"~%��k����pO$W�!������$��Dv��D���'�K7{ �=eI������ Ǿ�Kr4�x��㣠8<�e�2m���af;hЃ
Р*�"W������K^�|�;��@�=��<.�)���,U�s�c8<����?ɱ����v�G:�H8�`��K��Vk�M��I��A3K۠��X���'8x̵�K���-)�Ѧ�%��>�9&�����8������w_�/̎ۦ�A�}
.�����oxv���2ق�3� ��������ӌ���4��W͙N��=}�6��h�\L���Gn�' ���G�B��D����i��@�9
�#�]֞�:��JR.��6}(�����IF����rS03���|��m���M��*���M��P�q�{3������Fz���[��0���P`=���h,��[�j�Cy��R�<�E�.--�Bn�t��#�J*��TfJJa�(�-��i��Ʌ`��C/�K���-��[�^)�?Xѓ=�Y`��C\0���Pb/toX)�޿��X��Yl�~�O�[�Y^����	��gikC���yӵZ�v4ꓫ�M�^��V�r��w��,��ezF�5��"��`޼[�=�!�����'g�wk��r�dW��1r��1����r�h���6�ռ�/�n��H��NK�0�v�A�U�U���/����B_��&J�;ٲǑ1hU٦s8�1��0��|rl�P:����i}V�>�?ȸI}}�'��s<{�dVI��j�̧c0W!�PN|��E��5����eZ�f{����Z籽�K)��=�������:���A���
��h.3��O�`k��M�tV���}CsZxk���&qD�/%#h��a�֒Zq��1�|��3������x���F�IX�1	+�=�H�"V�����e݀n�@��c��d�����W�Ƹ�=9�qC��[�������xZ���x\������P�u��N�+V��������a������w����_x>:W8�|ٻu�@�7�o�ڒ�ԓ�U���Nɫ0J���5��G�M1ò�Oܬ��ՙ�����f7?y1p%:LI{V�naL�/Wë#ǼLZy����3
?��Cqk���������C��ZE�>ͧU����ZE�Q�M ��%��=Ӳ� 9�'��^|.����m��H�ler��o���������ϡ��!gX�nק;�R � ��v	Ag��\�frS�s�[~�F��̑W0����-�?��ʹ*�	�<�ɻy���H}�Y��f��B���� B>}j���ث;��yzءM�J�Z��]�ԠvktKأM�a�6�\giS+��O�Z������z8[�Z�s��\=T�X (~��?Kx8�B;�}��L]�KR'�3:�ʝ�7`0�D$�_�O��(;O���b���v���>����f��,����	�[0/�i�V�ȱﻙ�����w�{@L�u$x�F�'���O���w���!7-pk���(wkG�t.-�F�Yr�bY�|Hq��ʱ���עߞĤ���M�����a~�Cԍ>?��ʁ�a=����K�	�-$�ui�k	���ݬ���,b(��
}��\�5J�iH���?��<�hec�x]j�9���{7�{h@�I�.�d����vj*�)�ADy�Λ�ˉ�4B$�|c��V�o�x>G�� �x�������V�!N���Vҧi.�¡���Od��C������QK�\Ր�^��C��IG�l�3�������H]�-�oQ|�K���1F��8�6����;8������O�}��݆��0W�|�2
��l[���F*�ը�$%�Wx�0+�"�����
���4{l�)�%}T{��/i�{=�n����K�_J����0�i|���#�0p<�H�A����p_���_�~�Cw�c�uڔ��:̼T?�V���\���-蔨'�ҡg����)�+sw����b;R8�\�0�l{$�F��o��"�2;�hy��%[�%��zBoHn:i��Mq��:$m�2^�Y�=ĸ�3�cf%� �mMF�קF��O��z:��B�,vJ���sh�)V�{OpZe�Q�Om ���`��>�K�v�"�v�G�?��'�Ym?��K�O�����+��n�R���&q���4s�vȸ�� ��BlTҏI�����n+s��.S��H�䢶��xd{u��O.�9Z�)��gJ��~)�?yW���P�^���x�,=�+�dJ�����r�g�M��1�A[Y�M��,8q�`�iud�U/v�|��bg`w���V{��x-��j�ח�t.=]JK{�^����K��5�-�8,�kۈ�v���N�qC͗:SO���M%ѹ��5�)��J���7�6�9<)���䛳�*pP��d���V�lǄe�P.�֞aSΌֺ%��S�@�QQ@�.,�t2��n	���@W�T�A�*a�,bW���p�!j�*~P��QC0��|�p-�e��{pC�14���<��a�P�d�rW�	�b"������uΏ 7����x�d�"���Τ-�)d���Qm�[n��ʮc]g�^����r�q�0`⿃���+ߧ�b�H�F�b_Ȑ��� $UE)�4q�׼`��vr;8�`��\�����H��L���/k�AUmZ֛��Y փ���IAJ�8s� (�����r� KE��,y<�J`(����]'�ab�l�/vX!>�Lm\�˴%/��$�G�@��v�[ǤC4E����J3��Ь�/��<J�c��/.?[{~|9;[�M_@N�q6���w�����V�-ԓ���h^�����3�����U~k$�~ʒ���ՠ����[��G����*�c$�<�z�%N[y�
�b{�بӑ���7��I�˥���#����j�V��I��u�4)�r"�s�޳�r�0Ze��	5�8m��$8E�9pY�#�B{�S�X�a���\(n��^/���a��J��M���-w��e�s�b5�L~���ɴ5!\n!�� �G��.ՊE��r��c����K���y�L�
P�bg�f�˧VO�Șl�B�Up�d3x��d,�5�Ə`�ke�ԚF�9.+yU��1�(;�m\��]y�����w�!�7�GM{�7h�'H6m�;Y��CÚϵ1,`��ְ�2��?�����03��y�Ȭ��:�p^$_鋜6����R�7�U"|���|��1q�yԭ������ж۝��>�S�ob����Ny�`����'4!�e�$C���c�ޒl�����D����(�,_�e�yG�������u���K;��6,q}b��Rq����:�k}�Ӎ"�~w!�A�C3�&���G���cO��kwv����DQWy4-��r��A�M~��_P �[����Qd�`Y"y\ě������VT��#�8��T�������'d��^q��\1[��%��&�&��2����(�����	O�f��l�^���Ncֿ_!�.�˰�0F|�k�q�4X�����9��v�NӇ �ňs��ȥ�OsBҧ9��ڔ��I��T��gy�6�|�)C���y�i�Զ�DJ;I�u�����S�5�=��m�q���]��.L@/�#�����y��n}��rQ}F�E$ b�#��zgQ�����~;qC�F����e�=q��8v��aS��һ�����-q(�6�K�@�(mo嘠��u�q8��-�]��LƯ�p�Β���'�C�VԃK��CR!o�X�5�߁rJmp�;��:K�c~������u����O����ڝ��qm�)�]���h�h�	]�6�2]좝���71���R*����r���L����W�P/�f
��0*�T��挂n�d{�Ne{�	��[rު����hb�g6�{�Jb<c���6A�3(�3��]M�r-NI"��.ʯW���m����*�����/�f��P�?ў����ը!��&Rz�B^���b�>B:�#��sk�a�����3p�	Ua�M s_}5J E�,Dc%1��"�y������,<�j�;;خ�����3m3�.��$��]V�>���Q���i,�ٖzB�*ǖ@�a�`@|�@|+�}�]�{AE����n����dKk|���Y"�Nsz<��8M�Pc����i���J�$�~�C[P���Z8�O��<-,X�\�nCx�Vj��۔|z��z)ia�cl�0�iji~خܷvz�J=����'�Qe�Y�Wο�c����5��p�=����'���HK�)\=>fY�ܴ`��"A�h���Դ��+p87�
UT��	����0� >�]�%g��B�I=m<�>�~j�^��Fk3m�KI��/ȗ���Ug8k���Z��ո�����ߞ�{h��-t�� |Ѿ�Ct��{��B}JP^��*��~#�M�ߴ�u�,���ѧ矷Y���m�xo(̷�|<����Oq�}�9E9����)����}�)����))��MUΖ�o�^�U�6PǊÆ�N�-�5G� Y�=F_l����n���`�r��ѳ��K��%7,��y�W��[���G�Z���L"5�OP��'���	��������Z�i�$=�0��x�����eԗ�P	�J{Ceie�y�V��U�2�w�
����/_0_�r;�N�V���&��a��z�š8���hm��\@*γr�]Rl�\�>��;����ԍ��}��N僁�8�}a��3&�^tjЙ�Dsr��^��/QI�@�Vr������ X��O$30`f�#�#�ѐ�*qV�%m�5s>$~�?ֱ�RO��2�a�y3G���"�Y#���;S2����n;��(3������N>�����CB��������M'��M��u�y�եY�4�{�*yճ6�_��f���fD����J�%���U.@�cE`�?e��g��I��/������D�N=]ӈ |<��xΘ?��1�Ŋ�o%a�:d������;$�5��{iT1vCΰ	��! �n5���R\4�XJ�+oӺ̵bp=N�C���A�q 8��s����"��E�ɡNU�8\����2_��WK�n���f�y�?�8��?��h=�n�g����Hb^��_�90?�o�d�.����D9�łY�a+���r�Q�J��~�����RF`��x� ��Y�-� �kX[�������	ݿ2�\(�0�2�/f�@-M��ߘO=��5���ˤ}\d�L��B#�h���� !{a:ͺ��4��L��pq�'�0�V�+�T�j9^J�i��������+qǆ͙�F}6b{3�[T�" k>����:�s���g�H��*OM��8<L�a.�8�Fs�\�^���įc�H�^���U���� KR�[�vk+P�9�+T����"����m�����w�M����^����m��n���m��(<g6''H�/$�\��-���.������G^ı�j��A���L�1.�$�5�
�/���M9�%'&n'V����{Fc(�-,_z�]�&Ǜ2�8ݏI`�Y�����q����m�~��-o�փ�*�%�ZKo�3��]F��P��U(� �~-\�L�5縚����4�F�t|EހWp��)/���������¦�=��f\U��t�r�6^����v�9� ~�%� yOOO�͞�)ꧫ�3l������|�v���?z���I�����@�o!m���;�������D��Dy��}�{���?�����!hG�j�����+�q��k�URZ�j���՘�@cIG^���iڹ�P3��ر}7�p�N���Ui��e�{X��e���'��i��X���C� ����r�I���9�__���\�r����`(q	�K҆.��'3�$+�3�S�z�������#v>ųF�H8�]|&�DXJdݟ�[E*�e�����ށ�P^C}i1�d5G���%���n��&Vsf�ցNs���F�ҥ�kH�6���d�'n�s��*�@dqm3z�q�5'�|��U,H�5���͸H}��a�8�59���k��U�z,z��xϴ���Άk��"A��L���M���#�.�1����]�s�sD�%x;���aX�{8U(S�q�������}�`�p��+��"Zˉ�4k�N���׋����T�N��g�v����wX��_���(�9?T��t7X�c�f��RoA�|_����_�󅞀H�/�x����h���\��MX�eiN�+��\���~��M�&R|�;����NN���D�D��[���;���������#�EZħ��V�+$���7���9�xus�Y��%�:(qe�*zp����N�� �-��rp��G_���E�H���E����W����ݝ�fp�ß�VE�4/)�3��Ӳ���1c�5f(I.!���P�s�+k��6��bMi�w��?���8��A+�3d{a�GV���U�X���Íb��{\~u�9��!wY�{��7������9�z8�Ů�6vFB�,�7�on0�/��p���؞Q9�����:����C����&�]w����C.�w%	����r�k��o���Bc���h�~I�_$Y����Bg�B���x_d��n��A(�%@ɽJ3��a��ދT��5��g�i]Cy�m>��rD��J��~-�q[���}p=�ߵ���Ē3_�ʢ��7������=�{4e^����{P|�v�P:E��ș�t�\�J��C.�qA��rH��*�&~V��p*��r�`�i�Ro�0�Yz������237�թO��}�����.�����ف�h��.Ǡ+�6)�B���ye�߆��R���?�|�����;��j�%bK�
����K�Wc���&T)�g9;�d�,Ή�Y�z��|���F{U�h̝�|$����O�Y�P.�>)��������	|7�)��b�>Z��G�=�����!Ç�p���0��{�Oϥ��_Xk�����Lg�]�����G�wM���%�����tᅠ�}S�R��zY�x�9���cetMc��-������#߲�
�rI�(W�i�Զ>3G�s,�Q����nv�C`K����NA�y�����h��b�r�Ѳ3$.+Q󖓴�(<��[��^���e�����>�cçvg����f9�m&{n�5�r�n�s�eH���QY�:�H�վC�.q�"Բl)�d�Mq���%�"�Dȧ���?��f���r^U�Y��P���Mե�R����&������A/��,G��^,�}�[�߼��zY�>=�=+u����$9~c_�?��Ǉ�MX�I����fF��xK4��bn}{�v�Mi1z���r�қ���K4Sv9>�׊)+�t�M�]Rh[u{*���3�{��`0���BT�zҸ�=nI��CM���L6a�2~ٝ�wH;�`�!"{��?F}�9=�O�؅pCk��������Ͻm�'�,6�&������	m ������
�T�^�5�FN�y .�I�L;�`���|r��m6v�R� ҡ�N��2�|�ć��/���ɱ�~���Q9~'�c_�	>/E�k_7����k�c�s'Ƶ��h���r7U:�)7�FN-7Mr��sC�nM���/�&�C�.�����m��%��ҿ�3}�~Ǉd���hp��Q`�|H/Y^�������}s��~}R���Pe��IA|�D��1<�e�ױf�����$�9v8С�k`-�
݁����_'��ay�L����%u�5�L�NkX"_C]pGm������0���-��ƱM���̕���rZ!҅0��=� �a�.=O�4�?7�ۂ9�֊��e���xM���mW�9ױ��ѷ�1��6�mo�$��'�d�I~m�O��������<9&�����-or0�#��_�P�t�tk�\�r�Iuk�	`s�����Mh��V�>!A��]��z�?�Vi����&���z]�1�/$iN`�[�L[�
/�~=�=�ْ�/$��&�.&����������{Q��T*��g����H�Hւ;l�Q����_�ַ��Ǎ-f�ȡ���פ��7����A<�v\�q�Br�w�[���O+�Y{ǧ�HCu����I��d�<=����\�|�z�6�gĿ�%f��-ރ�8Y܋x1�#�h�A=P.���w:���6�t�_D�Vz�5S}���N��|�3��O�.K��~�q�~���k(����ه��Z6����U��Vd�p����lSΗc=v<w4t�Q�H�s@D�1��-�J������lv�oţt�e�<�nf/��ok�g�I�
��rR!�����̀��%�^/B���~#���f��U���:W�Ao��4�%0e/z�n�%<?�(aS��U ʷ�ˡ6��M��u����NϰPe�=Qw�0�C�2��m6^^c�Q|�I���H7T��v�T`��r�\��s$��r����ē	�5-Z�)�ޕ>:Z�M"�C�9�$� 6JEubԵM������,ro�����o�v;2��@�t��/�N���kڪ�M�aڇ��H�?p`�F�q�P޾�0�����&Q_�&��DIfz��c���i&V}��C���촶N�6��UM#�1Ȕ�nv4����rl;������	���"Lh���=�,�nM,m.���:�N�&`\O�e�A���mמ�ȿ�=x�}m�-�c�o���3�G��I�$<�lb��-���p]]9Q�#�V���\Ɍ4�݂\f�ْށ�P���Gk��"�=Xd�a�O���'��Ԧ�������[��m^�5��	߫�l�Y*A����/�B%�@s[�8#���	u���[6�Voi��G������[�f��Ō��lKɻҢ�~՟跩��z^��a��R#���߭����G#h�ň������o��:��7���.��ns���'�ľ��4�O�R���lV��;oaE^�2F�%E��#����f��NV�9~��iਨ�HdT��R��_c��<g��R��?�hiP�\/7����%���~�_�5��޿f���'���/���6"�`��U�,��2!��~;nK��I��
�mi�C[Z�z�԰oN���Z��;�iR��? dD�BH���6��o|E4ȵ��|����>m���p�k��c;8���W������̉�	3xC�H<fK�e���ڻ,!��C�/ ����L;��s2=K�JK��f�����y$c�3q�(l���O��>�iP�r@�(�6�z��׮�H�~�A���ʹ=�xG�O�CM:���u�8AX��Gk�v�d�%��~c��/X�YF����|ƫ=�Q�E���(7S�}�c�.��po��ű�}��c~nWmv�����#�fHtɵ���!�������c���Q7�G4<۩Iw�|Oאָ:�N��������x���)��
L�t�����h��N|o޲��.�	��T8��j��e�lٟ���ny�t'C|h�Q��U.s�*~����[��9C�w�բ{�n��⡜O��i˕�"��6A�,���&���K��C"u���À��8�<+�I^_\�W�W+��s��~��~�M)� !,��������Ma)��v��o�ܴ�e�Pi+	4���+�i)U~��T9T��O��i����z��?R�V>*�^�y� HY�[ˈ�h�f�b�E�'x>�.�B1�����M��ݯ[�S��LAh �sz��?<^��Vw��|��t���n�1Q�fG�^��J��&��-���\S�9o{F�Dnr�O�����T�/��|�Q�WQ�K�K����p���%p���n�5����T�� �0t��^9Dq���ìъ�Ə?���~��G?���I��`�:ʖ@ZZJ�����~��D�)
|82l��Q�/8��}�+ʫJ�S��B"gY-��u�f5��!&�q����ߟ��s<W�j�"&�~�$$�ۜ��I���$��a�)}�g�{��;�������B��J��@���Ӛ�V�E%��Cm}�{M{���&7����Π�����%6�ξ�37�^��9�����=��T��� ً��k�f�9��S��+�c������B����yq7�m lT��B�
��z�R��/ƕ���|7|�Y�1m���.hצ��D�=l�0;_�B�R�� п�MDR��ZAF��U�A���D��;z���M�K'�~ٵX���� >/���"�����Q�{�!I�b�Ӽ�Y&�h���n���������\@���E6ih�3�?8O܀�@ͽ����`縚eN'V���M�N���m�E��6��������¥6;�#�v֨H��ސ��aOJ��lΦW��YLʝ����S�i��4t<��]JC��t1��1�����h��=�օ ��?�e#���٨�˒`����q(�����l}	i��޹��H�)F�ΰR�l�s�e[�Y?�2W3�)>�i29#*��H6�:��"estI�i%	֞�����ة��f�����F������싗Ś�[�%E6 �K�!�B�#:N^�]��Pmti&v�b�ESk�i���x�wǷ�P:����Tk�|�5O��#���~�����	��Ӡ������!��bq}F�0�և�ܟN�-9�#����h&6=5��Na��ǫ����Uq�ݩ������b��#�X�����!�1#����%�i�y�kH�89`�{h�<�7���4�,D9ԍ���7��O0�cruL�������hƉ?�VZ�F9���$��K�z�Vm�N���-�Vג��)c�#
S���nl�ß
}jҖ�u��"��15u�w�<IB���a=�*j�o��4~P�*)�j4�^.B�x5�X�AMq�{?��+�Ж��&7ѧS�;yշ�/$	�rj�������^��/����0��z�?+VѶ����F򱦺�P����É[�?¾����?7MK
��hqݨ����V5�e�mZ�,P��U��:溟L�R��{w	��{Q��t���t����m�p*���"�z/A�������y��u�������9�y���I��uE�MZ�մ��6/9�4VN��m��c&<��:��?F�M�^�"+Sm�(�5�E���=m�0ȷ�,�� �/!�",lҷp}o���I7����g�!W�_B3C/+HJ%Ff�@M1�r�tx2g,w�]�e��c#/�޲k��I\;�����f�;QQ�yC�"�.AOt"���i����4�0l~h��E4���P����ޠ�kL���{��̯���H;�cVt�3��P0��г�}���eo������Ԡ���hw8��F�������>��6��ٽlZvrUO��u�z�>-_����cy�kX@���ڵ��+��Ӣb�#<%`hH�H�m�]�3C����A�7�Nr;a�-���][����k��x���ƍ�tL<,�4�fG��[Sv����D�N��4+�&"��>�}�K@�u�RZIO5�ˋ�ӟ�ՙ���'�>YqiJ���W7��f��nm�����Cy��eto�:|Z�?3�_�i6d #,�	T�bRy�͵�k��|}&�9���1��nuC�g��\�B�Df2�����ة�RԨO$;��`��k+v�p�b{��I&0�XB�n5�(��
����TT�s�^1�d��#�vݏ�m/������	�A��Q>�n�%��Wy����Ebܓ#)4�ɶ�J��j{3�u���{İ�zԵ����B�d�,U���*��e���`@�N�Ȥ^��E�nQ z��S}e:�S���>Ge�x��T������Z�к��h�F��8�?t�{�N���������AS4�5���_Y�\�`#1�H=ϫ�A]�$�q�>X��E�v��g�����+�c��y����s�Ѕ��(l.n��]�K�:}f�(�i$~�Q`��(�Rh�%�:K�/���ĩ��|X{L@�f1���d��^�9�������){�U����6z�<|6��xYBݣ���Jz�7�����
Fڜ��J�I��`����rd��v
���sd1h���x}��YM}I˵�d���3�E��y96 �vw�Oc����Z$���%s�$�+�#_ٷ'!�Ӕw,����p�3�!MK�k���n��O��:��A�q:�����0g]k�,MY>�-�Ac|�9�ۿ)�Q2 0R�0!x�����ToGY�g�����ga�!LI����T�_
����u�e4��	N��t��y�b@��!�G�<n���)Ts�����^:b�ź/�(�z�1,=�����䋦 +P��T��Bxdi�<{��ܪ��BQ�v		(��;}��������Cj�]�t��y�"�H��&�?/_��Ѕn��.kx�������
���O�[�zȤ6���(����0_�"���a�|�����+�x�*$���q6u��Am��&%{���1c�y�R`3��!��� ��� �h�܎�!��%�X��-���G<�������س����$>ڶw�]�u�D �O��Z���
�%9L��t��ޛH�$V����G�}X+_���ӱެ���k~k��"$�%�̯cJ�!�hJ��J��Ť��m%W���l�ܒ���_�sNc,}��*Bw�1`�c���/��m��_2����@���DrSp~�����-Ӹn{2��^7��L}�(H��Ћ*?���4Á3IA�Dd@Y��W�B�9�DmY�z����B�WP�z�U�ڥΜ[�:`�;X��'o8�ݢ�9�ڰL�b�j�4}�C9}��!��x��[n��Y�m�_��!xZf��z�I���!u���]~���o^�h�{����z�[�������[D���O��!Rȴ�r�g�12p�4.�#6Mmm�gU�izY!�~nN&�h�(<�0���_����~���f�vV�N+K�2�#��i��Iu��ej�qOB9�;�M��H��w"t+2�Ֆ�눂�)�(?��.̼�`�m�v;�tG�ԅC��p��9����H��/'�@�4߉������i>��{DfN�H�^�v��QOy�&�_��>Z?��wzU!�^�\��,I��Ȫj��ZW�#a�N�,M� <pU*R'H;�
��9p��Q:����7��ڕ~l���+'�?��6z;���&��e �SD3SG����K���i6���������M���t�p��kJ�?G�Wċ"���9��ٕ�h���4��
')���R[��u�i�~x�)P��doK}3W�D����ffI���u���ϊq֥���F=qa�փ~g�L�7g2��[>�x�j���Z�bWȍ_���W�ȿR��p��jt��C�LU�_�_��]���{�|[���+���>���ȝ����Z跑�����B��8��FL�d*	�_��qf0��d<��v$��m�%j�B��*Z�����V�5�v�P��>�>����O�1đG�B�X2���yg�sF.0oe-g���OJ�|�iR�vȆ��f�DƘj��E���E�_s^�d���UFt�\�n��� ���F�p��)lrx��^h���X�Q�[�2�Z�E����KR�p����r��;S�!��ʔp'2X��F�Z���:20��Z��;���</�׾��)�.�~PVK�<�o����Q����'s�B��|��??�����ؤ�d��DKv@��R�V�%o9#n1�r~�FqM�#���	r�>�?x�(��8�e]�Em��$G���Rk�ů�rġ�h���K}e�����%�>|�Fxõ��o���T]�c��⥖�	*��'���if���25������MA��B�Oh�Io�{޹F����r|�>R�~<<�?��v�`Tz�B;��A�U��P��?���V�%��3�j���⭺]��{Q��1_@W/gݤG�T�"C�! !��i����r/TZJ?FU�~���VxSG*�afdwA\�kȴْ��#��3���H�F�	��Γ�YƂ�$k
�a��w���r�g]/�O��H�������Ehf~�e���j��	�&�ӝ��*�^��b�iA����dW����W�@?�,���=�Ί��(�xf܉�i4�=ki��rǙ���b%TQL���Y.��/D�o�v2^-@�Xd��G?�p��7���)�[4 ��3�ϯ
���]�],촙����I�(������-ח8d�B4����8 ��3�J���Ƭ1M�<��+������Ww��S_�X��h�5Ϟ�{�\}5rF-3d�DƢ�ڐ\c��T��:"���s�"��l�28?���7��I����(F4��G�禚���ǭ���uG���Λ^��¯3&_��&���	9�����F�?6Q���|�1|��H]>2�G��
v�x��A�&�w�
O�|�vG�ȇ���l�90[�@�˶DR�<��5������ݰǃþ3�Z�@D��_]�f?��G��*�e�$�$���gۜ�ʗ�X�i�jk>.�TC��݋l᱑}9���u�S�W�C<���i+�S���?ݬDP���+�ᄹp�Q��E�<Ժc#2���d�g�� 7W�g\���M���c��?� O��"[1�ʟF�@�o��K�?u�\q��=��4z��Ew��^<b�������4V����jŜ�������J��+֗ L�����Fgj��"O��z�5���g��̧�OK�P�*��v��i�����DL��b<�$���#&V٠be�t�>�*���ݚ��� �/M�i|�L����+�4?(:�?B���c}��rC������D>T�w��_��*I��Yy���m���z�V���u�CV���u��������r�9$~�����
�<&!�����x&�#��6� ��!�Z�$��jz����*�<Iŉ|PK���*َ��(A��:a1:j����V*��7���i�!��!��Ә���5S�T��iH�B5@9�����z����0R�5���A$�ҋ��5�jE~	m_�����m�w#��^��ک�s��\�����J�y(�;n1ˤx&҂��m9�3���ڣǦ!M��*�����"���[nHaiv�ɻ���%��w��׉�yWB�7uB:{�9�C�E4N3����2�N+�0�Q�#��ڗٕ�����B�uѽ(����8�y}�|^��茗�yiT��%/�b��n���7*� R��"e��x�B��i,m��p:N4��,
B$��m6��c�f"�d�CJ��
��`�9M�N�-<�����`ݢ�bv㝲 }Q<0ю��KA���Z ����٬4F<�� w���� ��I������B�����2�B��%���(�
�c�u��oC���@��l=��]B[(��G�R��s��,x���d����"�^̻�߭��~���8�l�{=�Mu+��\b�F�}j�Y��F����9Ee�LC�kh�ҁ�<`L�x%G��t$4���7��6c��h�[�<ܜ�D~�b4ſF��k^�a��V�7�����O�J�����ؕ{������R.ʔ�W��qK	���/}�x-�1ߒ��rTjˍJ��H�ẏ��������CD���f)ڡH��9���w�|e9�����4W)��[\d�=m�r%Jd��T�,�&B��˻�$���)&�>:��B0����<�'��~qc���8>u�R��R[�@�4�'�|��&�fX��&�Rl���E���dEݿ��^�����wr��_���z+�4�����uO���`aV������|�p5��q5��\��D�uy��,n<�Ű�]�*��s"Ҁ�5����YM

��w��o�!A]�F�����HbEu���Eړ�EW��p�9�mL??��P8JYH
�f���1����[�������3Z-�᱿��n5�����J��$�ů�vE��D�}��<	����<���-��_�`ͤ�;�y���ҫ��vl����@<#�'1�Rm��]��T[���Rm`�|��(�����Ɯt��@
����2��=�l�Jo
�=�"}����2��[5mڱ��'.�!�/����콲ݥE�Xb�mi��e�ͭD7��I��N�b3�>������A��v���?���^�q�2�q�r�z�9x��vz���Ŏ���9LC�&y��_����GR�H�s��7~�~�jz��������Xi�c�ͥ56[���՝m,1+�4U�D��EĨ�Ju��7% �A�d�F����d��b�����fؔ������C���Y�M��5ppܱ��i��ֶ2�)5�D�\���T�5��Ks��`ڏ���Ƶ�m�����K�-��ֳ���m^8���U���;��x�4ׅ�X���n�xv�d�׋����n���
r���;Q�SA���K��̍�LR[+&�h�;��_?���߅~\��e��`Mmw��vl��h�"�͘-'iZA��Gs|5�� d
}^�P����$z���c�#^��h8��ud�躥���w�h2Ս���Yp��g�'
',0z᳼"��nvgZ[��F��$�Q|��c���Y����XA�6���y^-UY%h��=x�ӉD�Rm�����,iQᘤAx�$d�A�0O*r8�Vaoo/g�2�n�x���֮ˎ����Z�D�e�B�M���߆���f>ZpV�{�e��^҄���HBgI�渑��6
����B�X��qb��b3�/'��7�xm<Ӗ"��:�n���:m,�j�e@�gRV|o�T�C��ED}��#�J]d8�N���7� Kx��Ӭ��$�o'�x�={u��^jF��X9�L�ںC�( �`���a��'���'�ءI�u�ڎ'@�y{*����W�I<���'٢��}[�q�rY���l|C�>��O���m�w׮�8���Z��E��.�O��oR|[xZ�s����RX�U�;�(�,Nnف'��Nk	�����Φ�/KMJ�.q������7����m�/w}0����G�fn���h� o�dZ��w?I�`~#��9�"^5ϩ����ټM�y5�K���r�E���!�(�WWT:I�M<�HDVV��3�4���'���`��Z��݅jtIw�����ʉؕ�t-M��!�]�Y��9#��؈Q�ͳ7��aR sW)#zp�=���C�ᖧ����h�����g�:.�Z���	l����i����Pu��j�{�Iz�?b��܈�_����;u%^9�xUz�÷?D+�[֊�ѽ�����V7 &{ӊB���y��@^�|1l����Ht���>]�VP"#�e}f��1����4�;O�[]��"'ucI��b�4��o�X�D�c����0���G�ڌ�uH�ND:i l.l?BF�@M~�8�7m���l���`�ў�&�ږ�?̕�F��w~i8a].O��iO��_�XF�-̮�Pn�����Is�f�W��v���������5q�T^2֪�ΤK��C�������dlo�%�jK���:�;�x���o�v|)�Y4����9���Է	R���ݺ�¡���B���W�_�GA.�oML�w/�A;�7��X� �	��k�N�CZ��������(��7��Civ2���#'� ���6��AӫH�4�#c}���4��$��O=�ʾxe��;�Ə	������K�ȭ��b�f������az��4�h����:�|�h�������6X ������=}��|�n���km�Dh����Q�?r%I�Pף-qr<$��/��H[m���Q�j�ihN�iÖ�MP�V84��s3���b3�w�����QQc��&8��q*���۫��۫��
�品���ȮR��v7�!MtkQźՀ$Z+�Wl<��9���*���B�S�F�D�Q�Q�%p��y�?ċ����M��.�����FK����V+r�
e��*_�������~���|bx8'�;��xԚ�`�WU��񑌌�j��f���qP��#��}ۜ��u1E��Y�+�'��3|2�NKb������R���旰���|j������$8��8�|��"���#�h������~p���*�'��S�3�AՔ�8x�	�'��H/�&�=&tz�:ù|��'"����<�:�]wl�$:A��+Z��B9�7���^��fv��5�Hm�9	����K��-
�#�.�!�K�J�6����N���|���Mj�f'�wtQ�m�
�:�x���"f���Q�仩:<��ֽ�.�:,"����뮻�"B߳�/��?:%gf��GSl���d϶&�ff,�6��?��9��=DS��ã�&�#VN��oR�#%��iv ��mIFr6�m��֧��Mi�k��
�Q��4�����M&&<֤�W��?"˻K���6"�.ы^��Lq���b�u$x9���=�y]UVB�xS��A%��5�WH�G��}&<��<���	A��j�il�y�?�1��i�Z
��K<y���H�בA}�>WO�2�C�`{�4Og^gӎB�p��X*C����t���!h�"��EE�E�P[HU�QB��B��g�����5�S���OH�����2.t[팈��I@�镜݁��G�I�Gf���x�
V�⎹2��a�oe��;��������OO�;`��_Se�@O�������35^�JS[Mf+��{`B��Y���C����}�!�IR����ޠnt��Ss�>�S�6E�k1Qʇ]%~X8,��
.;/4ؗ7�E�٫�c�/�e~x��U�1qQ>�^q#1����o���1� 3H��4�#(Q#*��D,4��${ʄ��t\�vAN�>�l�(���]u[Џz�GCI����*��iQ
����!�K4�1�8�S�{��6�F����U���W���Ϫ��D�2ĺ�?�~�x�q���H�RD�Z�;~�փ|������ov����ի���g�&y�`��wg��(��On��ȸ(�3[Q�کV��*峧���%xa{�<�u1RV
H$x�UY��(�,sh��]"��EBg�n�%�rBsV]�iƥ������0E���.�B�{V_�F�u}-��T�`��;\!����X.�b�G�Sc_A@�W��	�)�13��q�����:�Ԓ�[������(us�r�����(�뛷�G� ��oPf)����3�B����	F�m��_�����ʝ�H�P���I��p�(�Ϗg^�N�:���dZO��n�s^2wg!�?�U�����Y"������h�N���R�)�O���4�p�j{��g�6kRs�x��_�T��q���������o�iY�Io��腣/�lYv#��$�'-!�Tc��J�vV����R��u���l�)Rk�a�L���H���;b�	+�b��w���,GY��V��x����h�/���-=�M��a��D�<�@r,2y��!P��="�G7����m��*<��K�ZC��/�������Ӝ�8�t�Q�Kj��tV��k���4��й��?��B�^ξu��H\k��+kݵ�{M�'�������E2�RO���{����vs�y�Y�4�},?��l�"���A�ʅã5���{����#[P� !�&�+gI�*A��&w#��O���丌e8?+�ox�a.>�8z�C�F��A݊|Zu�/�9����%ִ��}��n���uK�a7q]�-�˚��g�X]��C��.ʓ�����7Q��O2
CV�w�C�^��U$*��R�y��@@��X{a�,)T[j�H@���4ݓ����#�����O��f�T�
�e�vJ;��oFE9��kA`;UzP��q��}�p�Pm�3��#�����z��-C���ŗi�=�;.𵫳{8��_�H	��X����!t*�r�l/a���m��މ\�}�����>>F��b��>TgP����ͪ�I�t�R��݊�@��;C+�E�/FҜ���j�@+>� 5.��PUjE�"��e��0�>�����G�ix��l�"�D5ϿGKㄴ�2�x)t8� ����D:Wo�Fz�.d�dɹ��/K��1�&��EB֩7I啽��Av� �nVN�}�'/����|�������}�1���X�H[�ښY*�[��l�����*Sdj����{�*��P^~S�i���5���6X�u3�p��)!�r�pJ�����NQo�D����T���p���l�1.9�O��L��4��-�o�˶�}��`~���n��NL�eiVZtye�5��A�G�9!Y����йaH'�\�T�:.w=OKN��j��7#�~,�V+���2�X����:c{�.�����D��J_�ߵ)�!]��s3��g�s2�#�fgI���5�_�$�f�`�d�&�c�KD�2�6B�&�]tΰ(o(���=�x%[V;��H�_�e����e�xm�ɩ��/�"���ʈ��@�-�N|�������j�<%)�b�A���tK��Ͷ$T���7����>���|S �����J���~����	�R�yaG�B���U��BZطkz��_�֊�p�]{�C`m��-S��Q����
jeE!'����Yz� ���L��?Y��6e��+Q`�ߴ����� ��s.m�?j�,Ul�,�BE*�̌��Y���ؑ���,I|N?�F��X��5��\�����4V��x����~e�,@}S��kR*`�=��Dm	,Q��ݥ�w����+��4���	p%WP��ߖt�e~^{c�7���((�3A���C;	��H}}4���Y�����?f�;��^M����ؠM��1�(v�����g����j��P�e�4z{	x��,GQ����Q@&:&�<Y(��lR"D+�B�"\�bݏ(k�^4j�&��q�t����gH^pr����O<ƞ
㯯[�U5I|�k����x��-���c���I�؃"Il�!��j�>�c��;;|]�^��]�������4����Q��$u͏ņc^/�kk��>"%Èm��c�h�l\8����1�ɑ���`K,��8;��]B�F�=��% ����o HT���e��J��1|(t1�W�c6B'�9N�J0�+U������MHf2�;�m{?B<0u8a~9nֺ�����'�U��.+%�KV����{r��CBV��҉�z�6�ƍ�:��X)��(�+O_������N�Z�W���:H'P�W���5���\����ݦ�3nNX���'�Q1v�8r�:z��6cVO]�U���h�q�LW:���vC-��i��b�C)�Α�u�K����o$��{<����}N���8L:w�O���i͹�d}.��\��L	������YN�c~8<B�
���Eo���K�"v�܆����~R>���O?![G��~�ὐ9c��l}�	��Н'a
E�䳀����6c4���߂���<�|%�Gd�D�;[�G�ex�8�⭟��e"c�ᙹ����O���䑜^��4��ױ�~��"}�(-)���~ߙ�ߡ���'�Q`ՅvX)�a?B�Ehd}H������6�i��GFbC�}�a_5�:��ƅ=VYO���>gu��rF��}3r-�0�S�#G�F:����k�g�4
N�E��*ѭQ��B��~�:=��q��$I�@��
"�^Jv4�>v�����H�=�[��a��H���Y��c�k8�ד�l}���g�>�rl�E� �Ӓ��x��LҔ���$McO�<�s��u#���+9���s��@g��ڞJ���6Y`P��t����;�z�B"a�ȉȀR���ZNZ�I�-\��E Q����&��v!O�ɐ�.��N|.D�r�u&�޶nX-��
�M	�[��6m�y����{[�6E�����5V�Z����a	փ6��^����]�2�t_�ˊu4�J�+�ڵ�k��$�H�^H�5�q�}����$"���wU��J�����	~�������E�ClT��LאҊ@��tWn�R͖��8��}�f-� {
����m�ķ�ӡ}�l� ��L-��u�����˙ ��KX4��f�H�B�J,C|*̉�G��}f�J�-t���6Z �/pz�q�-��.e~�L�W����@��r�ߺ�f�6�ޚw�y��1n�<4��-� Y�;}�~�&@,7���������ZY�6�:��sű�н���5����u�EY�u]��ԡ�:�r$͓�`�	����I��m�\�/�x���΀jJf���{
�7�i��Hs�E?��k>�mq��6R�H����CaoG�����Rin�Z[������&��7���ܛ�n��"�<G'�^�	�3�����5��T$h��&��l���ov��о~��]ٟ��?ԋ�5/`Ԃ`��~���x�
ŭ��w��KZ�U����-��Y�)Xi"�1���'O�K�{����.�����r
 ����&��'�Z]Q�/m���9�
}Le�Z�T���@7��@�
#�j�R��O�ub�l��a5�
h�:P�Cc�z��t�)S��a*@bK[�tj���M����
����|8�#24�����j2W���]�>�=�����Zi:q�%�0�r(�׮N[K�6ڮ8JJ�V7a��'����ӕW�Zox��� �⼈
�ǰ&7�[�.��7�km������%<���W)�~<G��n�via�6�����*Ι� ÔcudH���:s,Q�a)dOH��}�[@�o��r';M]�w&�!|_����Y����f3��-1���a�Z�bl���60��koX�=��uB�k��$���m��oŊ���Rhy7�M跠������ڠ5�Xm�N����@����-}�V^*G푡R�Hy���y�ڭ\ZVþ�!�z�|��u�J���7����g9Ƞ	��5	����Z�g���ӷ�u-ZMs��Y�;�LI�h�X�����4X0���I\X�kk��32�d�b�ǶI��u8��.�{�Q�z_����g�#g#��ԍ�
I��*.e��&�N���r�w�������Q}�5���;��r�n^L�Tm�5��*�Gĥ��z�z�k�0��4�u�"�N��r	F�\�#�!ᐩ�� �o�Y�����+BH&�����ľ����R�?Q8��H���:��)�qdP�c�C{J `a�6釐� R�M��D��y��Lۈ�fe{?�%��=�6���"��j;��PbxUy��3��V�1���h���D�2xF�ǔi��*[h�~o�v�0'��謡�WzhQ��!ͣV9D�ծi�k�א���(�Gv���|D��HG|��:ķ|(_��_/G�X���4�"aH��8?��V�}���X�X��8d"$V~�X!���v����'�D������!hh��rH:�4�$ӎ!n�����^��7�f�Zo��^%������l�N7�g��C����?�"bE�A{	���"���hB����y��O�;�	xC�孵��a������m�/7$�u�t�I�JX>�,�d��I��*E�[�qߝ���T�ߞ�;V�zbc��q�#�F�����{�����T��ݦU����`��S�`/���_q�_<0�� ʁ�20��SxN�V7�r{՝m��*j=�-|���Vsq:�W6�r���7�N��-���l53LP�O���`��k�Z=E����Q����J�DU��m�Gx��,�+��vG䠍Tc �6��
%{d-���}�n/�eGɁ��T�6�w^��o�b%��=(���ٓ���k9����!1l�0d�B?g���!nC���ɇ�z�P05�7.��t�Dt�:ijXDb�����. 2VE�2���
�ą��,�,qy>���}Np�%�iEt�/��z_\-�7�%n�LXg1�~��yҰ���w�����J0XA�f�ߎ�I��3.�S��'�*����= �VC����+�$|��!Q�Z��T�3w���t�Yi27��ӗu�i�
��&bv�ZO�ƶ0�ϩ�%gZÛH?���[_�Y+��Mh��t$D�8r ��E,Ɔ6/�R���/��+�e.]��T�ω���o�-R�	\�^�҃}�ub8���Y��6�V�rt����Y1I1���Q6��_����6�����xҘ�L=6A�)�Re����	���mjK[���Ⱥ��kF��~
/L6�it�6%t����0�# 74<�i�d[x�~�~gn�x8�i�˾"���M���3��뵙Y�oC����Ni�F� �o}c�>�)}&�|Пs��״�D��v�^ї#{�W�iC�!�~h�#�;�%�	�����nz�%��,��w( = �@����J������NlL��t���9+��Ǎ�`���v�
V���)qçmE��k><K߈5���櫸p�h�S�S������D���:�ݤD�2Ezk7
1������]o���}����G�~���w���!�u+^�����z��#�A�5K���w�!o�?�7I��{��
a��Ι�mf�9iğ,�v�E8�ޡ�G������I�@�~L紓� tc�q�ew@/�=$����ˆWy&��t��)�w��T�e��H�h�-�����t���6���H"5�Dn�P<g����k�+�ԗ:��OCc�Vf��('�-��}��w�,�|�� �gojHM�i�$��d�ʉ���r4l?�	���p�G5��-��VU�%�����N��5s���<:(�/�������}K��S�E+�������UhP$<�7�[]�+Vb�(��@�r���w�9��$�2����k����E4�w���B�P/who$��I@(�q�����a�U}r�ij�X7�r�V+'�'+[t�\��eV�qr�Ca�i�r��9��b�F36���#QÛF>�Ɓ��#$
���E�Ü'�/�D�.��3�evz�K;�_�v�[[���Z�5���/Jr���h�%5]��ȓ��h�B�>p��$�Ҏ� 3Ćj�_�7��7r��&�Oz�ڗ�z�v
x�r)k��"g⏌iB���cC���h��[�O2(�n�Z�b��Dk�R��3�x���	�0'h{N���IvJ��c8x�-�/���ӽl4���պ�X&Mu��$��]w�oS�=�.}�C;(���9`��2氓!�
��NYy�9�!덟T$٩h��{z�3�r��e�rq�!�-�)��ಫ�e����J|'�!�͉Q:����v�N�~it�N#��.�
�9TZ夀��v������J7�@\�	���Ü�P|HǑI�����DqiuYo���8f`Y��.e�`�`|)�`��U�Ľ�dkR��� }=��cY�O�(�N,��_��J#���ɞ0���#������%/��d[Z���hg���y����V��4Ш��=�ꓻH�f������# �Љ��b$�1{��m8Cln���s+r�g���y]~v /7�J:� �U ����YL�90Ķf\.��r�.f��bv��l�O����q9���_br�u7[�F�%1��u�vh�&wPD�Q�I4��H���d}!��L�F�&'Ě����[/������섧2/���#�7n�e��ϗ4�-��.~��#;G2�W
�T�k�7҇"ߌF?�	C�͟H#�v���־ �uO[�[�B�:����)b߅��II���߇����U��C�;�_F&;�rIɚ���e����?�VD"4��F�k��Y����?G�Ǫ1��W�v���e��%�O	�}Y�П{�a�~S��=ƪ%��?[��kߵ�#��}�Ru>�7��hޟ�O�C4��x�7�DO�����pGݦ�͑��j�k�2k��3#��|����q	����u�4G��^��!����y��¿��w����N���a�t�7�k��&�6�w�'����ޮ2R
y�x���,�H��[@������u(�-�B���T�Q��*¥��E�^QAR�F��$��_��9��`l�S�F�I2��ؖ�+֧>Ю�=*ң\��͙y�%`�N-(�q+Nq�a�����~aj��,2g���+����\�}�(�NE��f�?�7۶q�v��K�~����v��X�+��]��"JR1/6�5�~&�5�y1�eu������̗#/�H�1'X���	��@#�/�a�֕;x�纥Ȯ�{3⎇⁊	<�x�M�o�&Ł�#�\��=X�EK��.�],�&�Lit���#����ki��:kK��ZA�.V�p�uG�����ۤ�`ٖ�@Nv�U�CV��ʸ(5a~�*ڞ��LG�Z��h���E��8;�GpU�l���y��mK�%�����a;w+�v�;o�>���q<��T�x���a�di�u�M����ek�4G	�Ä?A�&����T�g�A�����[l.Q�T��ֶ���D:1������W����"X��79s|�M���$�]�9|��S�����Ֆ>X�qEZΘ�J��H�T�EV�}�	�ѷ�گ����|Q��n6�A!$\���h�Q�Q�&��W�E�74w"��j�g����]���W�������H?����+D�
OsCC5����4wPc�?�ik7�}���r֡�.�e�UH#��t���c�F�r
v�5cܙǯE���-��k�ď��A���`Ɗʸ�
X;���ѫ�G�^��ELP��PR�d0ѻWҏ�.�(��L�}gk��ɠZYQ��� ��EՍ�/���*�v�m��"��+~O|���<����k�M�#N��3ڰ^��"`���Aéj@I�n�=-$\��v��yl�"�ր�X;"N,׳Rq�����mE��%rŢ���]ap*��؎K"F�^_.HX�?t�*-��uɉGGd���~!A1es<�����ɴH��X��Bt��&�o�/e�˘��nc�xQWx&�!2�p�G�:k��p�
?�cؿC4�(� �&r�L��K�Z����
Z���D���UZW�����j�b�\3��Ӑ�(��O�vB��E��}�GsT,�nP<E�z���q�F�4�UG���4^���΂���2���A	�C�Z/���/_��Uc�������������d%��$@I(���nTp��f�I�,qH��s�j�7��|�o�h�W_ј^廗]��J�ޭR�}3W�U�t���;�!�`����#�;���}(r���y���)N��'5�Zܱ.����N����U_�or�;�����~Z����3Ul>����۸��ghc��E�i&h��A�Ñ��L/ͮF�����W����������Z�g	�v��:Z����OE��'i&BZ������6/�28�!խ�b�):�9���w��w14����S��=&��-P߀���b?�N�)7�� �vS�#�V]6I�B��5<˳�cb�^�.��EhzN��Y����"���k���Ɯ[��]l[�Qѯr,��}sR�0^+��JDRŹ�nu1��vR�aGIS�a(9L=P�*(Wϔ��)2�D��34%ㅰ�.=r�;�z`~k�<���>!	�C���x�w9F}ϟ>SP���
��z��W�_�F��H��$x��`�
e�֣�������54��h���U�2�̳+F5G�S���GQ΋DU��f�z�p(�t�=J��go�65��n;:˦��]�������`c��Nya��v�������jY� ����=���䤬����IWG�z�{�u�D��<]{�b�t��)���
�a�M��G�e�x����GS%�}.�މd�6�el��3��.������eVt����]|�_wł!2-ѹ�~�H��td����vd���}/20>TGǮ�J��!����c�[]̳7������$K��j�����e����;0]SiБ\�ͻK+c˻�GV�S��-J�6��{�_�T�X�L�C>�?�������lϤ���hI}�[mw��)V�}¸k�6ݐ+"�Zal�NK[:�`b�:o�c|0Ar�zqގ(�6���e�C����٥FDAdA�x��i��r��,J4��O�F����#0�/	5ůF7��9mјp�N"`Q�#�����y��D3}��M<�r�+�i���X��7}�&��cY)���YNh�1HEǊ����1AzS�cL�h<:g*� �����{���b��躱|iq�	���:� ���i[�����g��VhРҡ��y�|��M4��B8���� ���~-&E�&��cVȑ,��1Gc#�W	Qa\��ę)���ҧ\M��*��:�G��*g�"�����߮Z�bm����Q�d��ߨ��3�E��f\}��@E �C+�i �Jo���?�"8��ܥt�Ott��W(-�Wly�g G4#��'߸��!)r�L�ׁ�����5�뗻m���#�W�d��ʷZ�Ϣ��g_��0}B)d���\:�������]�L�ܪ�T�?l����][��� �lα��MK�W��*�2����H��}K4�N�ڛ�3����pUu;�賯o^0�y���r5��,w���;��^�Y�n��!ձƦ]�_��]���QAb{��4�7�Ά�������m�C�����%��lǚl�)�bϞ����-I"2��s��W���3���Z
&����i_c�����W[6[�i���\�҂r)�jz�?uˑ;��������MM}J�9�}���ssu���k�]��������0�J���xJ��a2�~��%i��U9��~�_�z�wI��K���;�6��"���V���ڲ}Y�������uhʑ}���1������҇��}�Q�Ҝ�~��ݴ2���r���*���j�h�~�:v^i@��?�E��O�"��3�17RQ�B�^� m0;����*���S���&�7I�n�N�~��Hv�#�x�,�4��
��K����P3�ٝl��1C�βtEx���@�'�v:��bZC���^�T��2@����ݖ� ��l��A�X_�Z��Ԓ$��_�s(��-�	����[i쏲���9e$�����T2Z�xyD�3p$��a3��d������H�-u����Mê�t*����𻺰���א���oq
�oq��f���i��L�s�\
Mw��jlE"�����Knɴ��"�n!w�Ыж��>�Qt,sw�q��,K��6�;�oVt�C]�)�%iv�e�K���,�BW����IRk��n�_Ki��W���N�y],��;lf9���w�O����|�s���.,O�{��O/���}=[���9_=�ߘ1��<�g�}�G)U�H���L�o�C�B��K"�\�3��{�2G�¯��K ��ĔJ+k���Rx�a.�;����{9��A�(���[��������m�5*�j
��2Q��W�_�1�p�##!K�2���O����mu��h�z�w�gn$R绍��H�x�JF�M���C�]<��3d��.�t#^�K��6��x�5ځ�3ӌ	iR�
E�S(���]3����u+�YƱW2��o���`��L��6�a���~c��7�Q��6��6��Xw�χ��q��.��iS��A�ҠA��oV�;�B+�64�y��*�,)�񗲁���.6����ի��sʡ>��&��q;!CD�Y1��,�<q�O#|NG��-��b
�چ2b�b����ド5��h���Ǔ�
'��rs����x��"�/@SjAb����w��
�yR;e|�927`S��?��/fC�*���Xh����7}��h-�!�.ׁ��n�}
J&PK���(&-5/�,*u��ǅ\�6��w�%am�$3��������u:=����Kud�i�r]��6��8�smZ�W�"6��>��Bk5f{�S��w�\�ߥ��m%�����9+�d����	v1&��TNݩ����i�)n"�q�6)D}�h�=� ~�PE�u�h*��^3����M�(�A܄�����f�U��dz�Y� �.s��L"�$�����i'�(��Ӎ�cs��!��S��|�5Z�|+�X�Zi�>?h��d�F�Ǆ�t���և�?�ۄ4;i�;*A	���k���l�"���g�!3��F���L����V=�֟F���G�������'�����q��tEP�۴��U�''��$z},g��xz�o:,�/��nƹo�s0^�����j�PI� �P�w�e~�E�|HQ/� _�ո�(;��� �^�s�<��J2��L`�|�D��n��;�P����A�4v�!���T���B���?dޱJ2�iם�������i��G�<7� �0�󒌷dk��t�k2���~TM�Y���~���W����2���gl���7�g��NIx�v��͞��3o���?� �����3d=f��,���3��0�\O�J��ؾZ,�sW�u����"�T���]ݘ�E�½h`�Y϶=w2��c*.ob*��mo�Kp �.��4��g�3q%���Y{9�ٺ�輞�Z���Eb���i�Dh��T!�{'���e�g9r�-s���٣;a>/�����+<���,�oWP��;˵�pD���i뛙���33�9��Ud\�U�����G�(1|g���1D���33��=&�u�����K�gﳐ����<���/�g�g2��;��ޞ�l�d�GD,!K�����=VB�"�S�������S�]����ؑ���fx�4�U��V�E���� ��t����ƍ��+�*'r����u�o�F�J��y���A�FѢ���r��|Z[�K�,���&�"���L�,#��m{���
X�Z�W[oȉ��#ׄ��N�eu���~��u�\����{>-GE��3Bc���g�(�ϥϼl
0Wf�V���O�W�M =���W�9�[jz��a���[}>�&��IᬆR@Zz՝��)��~5	��_����U��aְ��֐��^���-���]�e�:_A�82%��k��U��7��/g%|F��:�(���EV^���kZ�e�i��Xv���f��6���zY�Dn�k�&��jM
}LY�ڂ���.T�ǣ��jjtf��M7�$�A���e�x�O6�ztw�;��diU5jl2)����fǚ�6�g(S���l@�Gv�M�j=3��b���U%�b�濆8�����0;Y�-�%�䒫�Q���컘C�÷k٘x�CZ��b<�9}n�VZc"��X��I~w2!J�T(��z�Z��`���2���^�-i�7����&5�m�[�F�
�������^���{jD>��x?�5�j b���/G��8)��;�� �e�b�PY3�m�&K����,�b�/�ʼ�u@X��$����PV�F!C;�F�2��ygㅛX���W�T�_ecs4k�c8ƜB�
q{��(8����H[Zs�����=ˁc@3i=��A���p`�K[W/�Ɛyqs�������aK1%A��]�eq̥�fG�L�&Ũ�ˍ�-���.ґh�QȦ��f��nΕG��)q!�\G��2��,6���y��׍Q��� 2R_�(��_e^��|2�x�y�.qrHnѐں�S�,��mӞ���Gt�N�ȓ��͑�G�� 9�-�Mշ
�V�|��W+с�%�B!R��݋��=�?!������K�\��'r�2��ƀ�i�&���w���=4k{C
<;D�c����T~�m,��M%�:���2�F����5/��*�㡦���k:����`�_p�r��(a.��)8�\�GOiK������ϡ#�
�"�jժ2�`�j�`����:��i���Zi�VZ����F�m���x�wM���H}^Dw���.X�U�����[W��;�Zn��j��pWSu�2�a<��;����C���� �>��H�W7�)�"�aO���u�H��")��I���2~x{�.���I}v��ɩ-��;}�p
�xr��S	f:���U�+c�@|Ra�%�q��An�̔�
�iQT� ��6�)�/�^uH�(`�Z���3}l�#�U��B=\`T�5���mDG����=�؃vl�W��^"��I��2�^Q�'p�<k����<Osw��]N.*g��A�N/�%�NZb�
��x���nsi|����g�s�Gw��4�Ӯ*O_|�`2C�4��\6R;a�Y�.`)�]��t��e.�(;B'j�A��$�D���͖E��`�,0�z��A5Z0�{��� ����%ܸW������l&�|,����!°�7J���I�6��Łb�,9\����-Ӆ�\��ȩ��hw;ՖR7=���G&di.�2��E�Aa2�޳I��q�ݦ��|5����������7���x$Y��]�. ��%�9e����ã��2{h��1�Dq�ȥ�5�!�����]@z��M t m�f�K��'Q�-�:d·�`�#�\3�	����GX���١��w7�s�D�ڥN���6�Z�v���L��Be�%D7�����Ae9���}����|A�ݮ>?/G�A�'V�#t	��59)��w�+4�X:K.��9�ܜ�#����X���Z�B�c�k:� ��]� ��YZ=cx �WH�jZ*�y�t8�/���d�����������U�z�U4��$�~��(�d�|�Pm��r��u���_��!X8�D�VG�M��y��F��A�ͼ<G���J��+�#)�t<$:��.��E1��wgs΄�4%����^W�&ݟ	��rp%7��k��~f���ez9k���xc:[�5�1��~�Y�~\M���H��)�䞡��S��/ȉW�x�3�)�;�0�pȘ}��s�/^O?��|(��Q�����4�1�.�V<g��8!rY6$��1!Ḓ�'�"Ө���!��D�|�����a�*;�̔؏�E	��Fs���$��g��l�mx*�?��\�+�Ƹ⩳	Y����GHy�(�[˫�ͣ����4t�x�nkSO��� �6�̩/`J7$�'�7�d�y!�:U3ZDA��ˢ�ҙ�1Bʴ�{!K�h��1�&�K��ȈgЙ��ZyP���ƾ�$��+I��e[帡L!�r��	lHM29��rYIp36T�K+π� m�7y��,�
��U����!����a����8�4�~p��-�Kw@v�����]oM*����<�מ�k����Z�`{�:j��F_�J��H%���s_�`�C�e.�50��,�S��"Ϧ����N���N�>�'lq��6���m[u)�O\QWtەdU�Ki��뜃{i`j�@���ȱ�D���vY���I��0Iw<gs��r)���Y�;~���8Q$<��Y� i{�d^	Y:�έ~$b�j�-��ɦT�8�����ʂ��N=!wb=yG��L��,e��^4�*����	�N;�c�G��L���P�2��$zP���3(sl�x���c��m���O�]n����h�[E��uc{)~ﲚgEe�"a)��/���`:�pa��V���q�1�x���,�;V�����LY>Qa�Y�n�F�̮K�&��|�,���+��0C6�9-�lr��f�~59���L��UL��B����W1ũ�]9I�~+�'��shI�ؙ9՘��`��D�^4Q\C�$���0!n��鸠9��3��~9��!���Eź]�W�L���ѷ�+{ΐL<%�,#|2����i�j��'�#56Y�pKxG!+����82����8�،�7�8��i�l����g���\�����!x��թ<G�d�Uc�ODA�4V��/�ٵ*�9�+_^���BJ<�W~Q����"��n���� �±����%���A3ss��!����F|�9�W��Mz�W�L���p�3e�[���\Ы<%���y�M������o������M��!�Y`�����jԨ��������B�HD��棒V��J%Bpv5�q)m��Z���ֶ�{	D�	���K��"��!�5�\���ϙ�$���}�W�;;��s9�y��>�����ݽa��kGP���8z ���5�!��'�4bΥ��?�?��ǩ�T��{>�����a�"N��C悇��9�瀹��x��`�n��"� �ԤU�����E5J�61u�j������vY\� �b���BQ�Y���S́O��>��0
��3��꒯����G����FƷ�Td~���}��̱ڔZ#p���>;F32�{j��ߠ���/o�G����~��N��xJ�~m���1�h{[�i`$^�Y~�$�<���b��!�F�֝f6����y�$գ��bT�~&���,}n��E�Y�*S�w��8��Q$k�	������� ō���g�Bkq4�s������ѻ���%��F�lz���K���ҷ��Ș�F��Q;s؏;�&v�>�zy,Vk��.Gb��*��1.T��Do��6|l��y�֋e����9��Q��:α�ƽ+%YO��c��w����(u�(;9c�7_n�i�����j,��\f͏ޫ*��o��u�	}/�=8�9L��.�����29�7�c�9�����AaCͣVx���MN����!���Lcq�u�LJ�ٮe��}�U�5�:;ukx�5-�DM�W.��Z\}QP�����ۍ��" j7g����5�UpȺe���խ�e~��w}�~{���dU����b�zWn_�dK����$a'ٸ�i0ޔ�h�0�������R�}	�~�X��Ȋ�b���/��\���V�\�����o�i��:�2�í9������K�U �X�$�qq,�`m#�y\�w����D<6ץ_LH�*�2�u���;s�p�0䇬��&�U�۽�3�c��.=�E�d�X?�#�[�'�}�Wѽª�0'�"NY�Ǧſ�oT��uo��~��Q�ċ�}������宦�^�B�D�
b�D�U�4q���y<۳�aj�`Y�ة������u�w Iϧ�]�+GdW �%�@&'�_��D�� Ç>%z�D��UҦߗ�ŋ�0+�җ�� kh<��?9����IC)����0�G����@l'VX'$M��,% T+��.�q��Q�{5�������q�-|�e1��4^����1���ͱyj��X�H�/�0�X����᪡xlQP۫�w�s�Ѿ�Qj"T��Hbw�n��^�#��*�ɼ;f�/�R��-JR;�E[�P[g/>���U>VZi�r�Eyǻ�6��A����"%��_+��U��ڪ �y~�ѳxY6������	�O;a�;�p�e[�υ-�7��+k"I���j�t�h�A��z�ڱЬ��J�]Yj�r��������dƙ47���h>�/t�ږ���FO�X�gC��?�x��Żk���{��}��xν}%S��zR0ቬG���"�-��g������D+����?�ü�gY�����e:g��RU#�݇f�XI!]v�m�M��뜝�X{Y���~�����:u4Si�}���;z�cd�J�򺚡xO7������G٣<fi3�<��Aa�A����̺��ҩt�Qމz�K�p����ַnsS�:��^ A�'��9��ORI�ݴ��>A��VN7/�':P}������LA0�I�W��z�HN>sD������j���L��߈;6�
q#Xy�mZZ��z�s��Gm�w|�|V0��ζu0��No1����Gi�{q}�,����K3-62�5e8��g�����V*T�!"�N@�zn��s���@d�`�Y�&u2+Y6�]"��3ohV3w��R<�,�K���<��n�{��E�#�#��,z�P�X�JK������� i2�g��W�9������J����4g����nb����{Ŏ�Xُ!Y�HJ.����Hv��"�kx���X�����c3$��=ʋS�K7�|�����u~:�ܙ\lI����^�+c� ]+�/�����> s���V��v�{��	��Ĩ��r�ʂdW�sQ�O⽿���BEz��<�RmԂO�Z*�ɩ㉺}�2�i���9�����i�F��2e�ɘ9��7LQ�Q���p&4�v�&xr�`>#;���I�����1U����g�^�\�b!1kd�jW`��X��y��@�h��ά�2�4��>��,;W�7����V�A��[iz_��AT�.�(֫F���%���3-��JS6���8|Ti��X��X��&,L�2�OFq���U0(-�s�����h<4��-�N�V_�^�Dڜ����1��L��F�1:���#����ӆ-p����1q�J��紖;  ��u<,�6�}�'TX�7�\�5h���f�b�J��c�M��i����5!��`zo��I\��j:�{Zya���$ji��=W�s��\́ �X�Vʺ��3�H��ܝ��:�Wd�[�} n^�'N�E#l9Ay��28�<5�M�~>b��R���(v��?�ä��#��#���8�n�!�A땨��!96K�p�
�������-�.L��s=̽��l��{ج�ҁ��d�;�Kk�d�w�.A�曃�J['�l��^s�g�s���Y!��x��A��*��Y��D\�O锠R���5�tZ��D���f��W�n�H����#�Ԭ��sD�x�v�0<xͿ>g���,p�cu���	����kK��hӑ-a�K�rkK�#�kK�	�hK<z�W[�ի2�%zU��$����ħW��%�಴%Yz [�fg��f����\�`-ڀ�� ��x�c�B����_��7/0,�Hoj'�\��\~�AvG�Ɂ�Z�~9\9O���R�!�l� �l?@�.	�&}�K�T��ќ�ww_��$�y�^�W��K������ܔ�M�m�[_���j�����ԭJ��,N�+�1����.�ւ]�9s�L�=�}��N��r�Vi\���6ȸ�=��{�j����4�l�=��PvL��0�r�ǡ��q����0/;��BjM���C	����u1��+���e��M?�}$��|i	�}D���<�I!��"���5�%� }�%l�(	�V�a<�ˉfg���kaQ�F,/��<#$G�,H��EN�>�4Y�-dݑ��j@+�˻�j�<2��5��C����;�-��M�H�V�Ғ6C]�B��$!b��%�ͳvx^HQZ��F�ڙT�MW�������f�3I�>M�I�4��.�8C$���5���6ݭ������հi��=�ukU�5���m��^	��O���o�O�!~AzJs�xN{�n�����Bs����C�iD~L���yvF�=�lr����2�9�'F��=2��4���n8���Tr�a�g��w�`�Jq��e���Y�N���o���� ��e��N�J�p��:�~2U4Gt��������,� �M��+���o���h��bP��Sٰ�k���Ά��d��)�=�<���}oR8��x`J|fȗ`{�4�8��۴t���{'��5`In�������S�±Z��ƃr:�����.�c�j�_{VbD�Gq�Q��K@*�����oo"��nX�L.�������T��a�u[�����i�麈 ��tm/䡗�)+87g��4�
TL�����x�����-�}��CD��ә�f[2���`�$�aL�/<L�Ħ.�o4Wσ�������D�t�m�g�ߚ$ˢ��{W���I�!���vt�\@�=6^(L}]e�uU25�.�7��+�K�UV�o;6�V hV�҅e'abCe�%|`�ae���v�0l������U�~LMns���Eek.n�eI���e4������D�L�BKצ1�Y��}�*:�����V����;�F��g6�ަM��s�M|.�YB����OGVR�L�6�N6!��1���o�l�v�{	��XM�F�~�*��SX��<�b8qJ�B�VMn9K�C,BӖ�iߜf�Ǭ�Fal�Vo<(�;�c=��b�t��N�m�(R��Eb|W���`���z�*�M2̼ѧen�sqj#yM�i���;=l+�6{�G�v�,ֵ���2T_�q~�P�,����-��g�b���g���.,9����ӺB�n�K 3�=��	�H����f�p�����>}��`����d+~_�>�Ɣھ1H)�`�*��a�G��5��[D�Q:��lDE���S8����_��i�n�ܭU��������D���ߧ��;���}峈��4��4?���X����҆��^���~P��2����6Yz���*`1v' ��S ���ʨ4h⎠Ί7HZw���&��elBy�N�#��;������.�!�}�c���-5�5�E�I�x9����>�s��):LZ������X����A��|<�L@�6�/HC[&�-ߥ���5К,�Ҫ�6_>�wj	���<�����ѫ��zu��W+?��>�7J���>�B?	d����|���D��r���7�k���h�O3hf���v_;9�
��>(�+.�W����Wr��ŗ��M�q�?M�`ԭ��d{��I�F�f�R���tN)x��G��-pL�p���Ѽ�x-���BA{������X��Y0O!(Rq�wx�쀾�L_���,��QI��h��$֭l\�����x�$��qA�:uvMt���W�;_{���8�C����),Çؾ]���R3��ok;�c��Nj-�"�j����
�R;�+�yV��r���]�����)p'�ܑ	��y�z�4���aN{��x��
a��c�vY��&�s���	�9G�SDX���4S�M��$��`1���ŬA���Hh�=�'d�M�dbʭ�5�N
em�/&�,s���N�?��P��91�ï:�휳�nכP��gԔ�F(&�𢯊�$�[��>8��p�>T��M�Zx�^�_�֭K;��*iN�w�߆^tp����кq���s�"�{���������;��/p+�-O�	|�1������6�ڟy�q��AVv��U9Ȯ���8vd���̲� r��eN��i���\K<{�jLP�I����Vd��W�sC[��K�=!?��!,]�`b�A�k��kd���Մ�]I�;�`��a���	zyN�����X`v\�l '����$�5�3IX�'�ʬ$�ײ0E?C�t�WZ��Z3r�b�C�`�ò�nN�DO�04��^��q�r�Z1͔��Ez��^���+�bo����%�$J�Ҕ����Fm�ҹ0�,a�$RR�q�53���;�U�54b��E�U�s6!�)J��ɒ[CNtg.#e��z�"y8�6�'O~��y�HV�����E��xj�p|#�:O{�,a>
�Fl���an���)�n��H�U��9�?#C�R.�Q�~#夹f��\��|9�T����8�C�0���E��{ɹ��a�Ɖ���B}��=��2����9��?��괷q)��v=�īmނO�G�r8| _�����8�"W�%x8��N�p��-ӫ�1�Kg�'$��rS[�6E��f�5F�E��)ʍ�ug�S�@b^j���J��{�\�X�V�~A�п�RX�^�c�ű�����
�V�R�}�XO�K˿�����I���~��0�֬����0����t*��f^��Qօ�O��h�񊋝o�,�!@7� ���+���vi���V;�)Y3����\v7#���Y���ͥ���ř����R��J��9@�\]r/�Y"o.n�<D�"��L�^G�Y��c��;|z5�7ie�wu�OuX`p���&��Y�?�C�iϲ��M�����9t�T�=����<�*�K3�ρ���m|�	��ߕ��qɜR�l���}���ԧ�x'_X�tRA�x;}C5X�d)-w�h��g�D��s*�l�5��^G�$3V��Ow� �m��ь�C���صNmQ�(,D�= @&}`�MR��% ��d{�ć���S5�+�f�vɇ7�C���U"�%pGX>F2�a,͕�@/AI�\]r�Z�E����n:'�ŕ���W��&+ɃE�N%zq*{L�\c�G%E�?���/��8-�Wdy+����Kii��'asX6������N�x� ͉�R�gLq�2�����'�5��8�N�aYZE��8�z��e��H[h|�t�8$�E���RA�&hJd�D��'`��I���DzNǶB���4�]��QV��ym��=1�n�l�z�=����J��a��,Ib�#������G�?t����wķ���.�a7�@+2�Tz�*�lV��f�}�	W����X��Ł{��G�tE�m�u�!7����T~5�KLE���:8Ǯ�>U�J��~�_��e��څ賕Ň��^730}Q�(���vA'��_�Z��)�?JP�"%�5+��l-r$܋_`q��u���J���qY|�ZL~��h9��������۹ Sw0�= ���љ�ugw�~���]�l4�#����i�_�OZ���}�%����T��8P�%D,��b���^}����I�|{����j����ꉢ9H����S��*����4��[��x,$��z�-�9�B�Q�C��}u��C԰�7��Z�|��F�m���s����L���T��D�%�K%c�"cN>���q�0an)�$�(A�<��+0瘗N��1}�p_r��T��tܕ�ޝ���)�B<!�,�#�o՝q�7w��G�PxC��3�aW��C�x��P|%�J9` I�b��'��i������#�����bU5���cϊ�3�}/�ê�Xzw�6M���E��Ī`�'~m��j�Ca!"�B=ۨ�p�krE�<�6X�A\����Cq�!�U���}�c�^�"�/�u����䔹R^�e&�ׅE��1�-G�/��^�eG�9�dzl���9!k`��S7bAg�6ImCN�ķ�Π�mr����1�9s��Y6�*��8D?��8v��q��8�]�D�D�^����7��>@��s?1���-�e
�ł�︵��Xn��Va��;��	���@�!5��G<>Αj��Ĵ���n���+�Ȳ��hz1�/HQ"s&&�<Gkq��j���c_1�e#l��|���*�.�?wh�k϶B%������R�l�K�9���X�d����yR��c�����p��.����i�_��ʆ�NaAT�.�i�J��j���
�2��Iq��0r8����J�;zНPE�p
�Fi�~�C]x䢓(-��NiQY3ͤ/U���G�w���>�d������tS���(��O�p��-�;ц�cp-r�z��s�q���`�Q۪�ح:�����i�9.;�~���|��d8+�����uG�J:мZ�d7W$1��b$_lͳ?g�"�+�� �`[FĈ̛2�d�c�aޓ����{r�+���R?g ��L��e��p�l�v�%%�-|�l�G����V���B��6����Q�,M���ɧ۲t%:�?l�k?�O\)�����/���N��O�l�;��i�%���ԕV�
Z�Y.�i�qN���C���0�����5�N,�L��h+p�������l�hh6�
��rB|������}�Y
��q�m��q��h���d��9ɑk������Yi,�hp�Ԡuj%Y��7�+y�P[l��9S���>�v�iK!����#^~G�q������c�p��/	+��U����%2��
����T`����X;!
�:.5����)r��>ZU̵xj]�hP�>aK2.�W�i�EtSW�!�M��P-@l|$zDꛓ��ՙt�g@ݫ3�bW��<����΂�*ѽő����d=a��@2�̿�}���Q���/r�p9���9z�7�/�m&��%&��Tz��,x7|��/�~S����|��4� ��q娖cc�Z�_�����M�I_4	r���Ts`��p������}�k#l�U���K��y3~��$�-Vg+��=��q
��m~�c��5�y�������䶙�Ǚ7�1�:*Y���1���S�.e6N_+K��O�b�B�Ώ�B�r������K(62��j5�Q��q�g�V�e��3,�`���P�|G�N>���,�eg3èbW�j�&^a\����2���en�[ĳ�F��2"qN�I~�G%3���r��b�� ��C����Aw�#t�(s�\ዢqV�hZ}M�?�&�j#Sk����|� ��F�ϩ=��xW/�����G�%,�)8Bl��o 9[wYl����Ğ�L���ʸ0�`@x��΢��
sK%�J�����1�F�z��(� �'9RMvrtw7��Y'*舗!!���[&5��B���g�f��䴐;?B�<��������؋��'�}_(2j����H���k�E����+;�G+�bʮ1�K.p9F�M�A�c�
T�+�7��D�,�Y�dM�1퓯��p�t��9��P.���@gy�*����]R3�`��2�7|����&�8�?b���gO+M�����^��1J��`�����39:����YW�u-��YG#ChT���u	��>��y����[�}��Z��J��b� +��U{�<.~�J0C?�#v��_%a�s�Q��4>�C��_��t�] ~�������q�8[�o�dn:+������㨡.�$���î̔otf�t0��/�-��d�;���r��s0Cp�k���{����x���6,U~����Q<�^��]ƏlE�(N��I�C�ջ�@�cƝ4=��m��pT=ns�:�	Cr��f��{?9�����Z�1����|�h<!��$�18�Y���x�,t����8Y�O�j�Ih�k ˜��X����V�z:[1���_�	�#�,�h���y�R�h͇l:M�h���ٰ��>���1��(�ҷ���B�Q���CU��Q�Y ��|�߸�����_�o����>H4{�MN�>%z��܁�����gR���hF�Є��]!%z3.,��W�H��>S��A �<��!<�BB<�̀aK�ǣn������9/d�{�"���n�^C� [=O�y��"��#co@{��X�ߐ�j�H#�.�!��0Su9ۢ��}9���Ң��"�[��4�U����K��9y�1� #�:����:�]!mQ��yEt.�	]ݯ�慒��|mE���z�eǘ�����-����V�cuI_�')I��sw�|8�:U�[֫�Jd�����/�V��o�-+��4��l�����aBɶ$�+�C������Zi��R��p֧����EX?�Ԟ	���<�*_s8�B[�z��q�
f��p�~�O}=n�:��y)�yc��KX��o�r
|�v�.�QD��9�?��gOW�,t��.e�HtwW)�	�����l�ؕ���z���E]�\1!��\+���}A��M,�m�P��ܧ{؃��m��)��`�ɔM��t�q1��@1˸�b��U�	5��$P���GG�M+�^2 6J$�!�)��ֆ8��Rد^3)����Do�"�]kLq�BI�O�&�Z�5&�s-�^v�%��ϳ-W�q��S'io$
m$����3���8�R���{��s9J���4+eڿ��&g�n�L{���{�N��ٯ�v9�g�U�6��!r�g̀/�ah��] p]ޞ.���4�۹]���ơo	#	]B����H��)�j�諽+0�ٖ%�<I� z���0��rڬ�*��Aoχ�Qrw�� �,'-50�Kf���R�f�'	�}n��r����e���t���7�A�B�ʑ�磊���k��y����<?�K��SI�9(�b��P|��`�%�q��P�~��U$ST�rZ%�*8��c��0�".�b�O�V�D���\�ca�T=:4}0�u<IZ\�7C�CoM�'Ǐ�����2�SGV����C�t~O��QN���=��HM����)����*���O�x[l��&�!�!�u��d���C��U�8���+1��HAM7�u�͈��i������1�t�VO��V�稼|�|=H�oN�Ou�������(��B�v���#��E��c\�ސ-r�d�rg_�<�q�9���-�s�\5W����)���	�'��C&,6]u�&uf�7(��#.Ė^�gʒ������d����V6�1��Y�o��~F�p\;\���)�����|*/Һs�W����W#�n��DA\h�Ѷ�>B����uG�J�L�֗d �����WF��͐�-��9�@{)6d+ٚ6?���"�K�t���������D�I8���Dp���4OJ�	�>�(�&Q�������R!���b����Ğ`�Z	ʆ=;�UXy��)���i���R�'9Q�C�����O�0I|��{�ee��0�m|����$��A��ƻ��=(�����mI2��b�)�����LVD�/k�%��ݫ6�}t:�T �__J�]�Л�N�r&S��5�P�u��bz��}��u���c�XY���!A�Ӏ���{�m�p&�Jo�zȽ��)]�~S|��؇���d1����ɢr�=8�cX|X8-lB*��&�!�Yf�6�@����|b؊���f�;�Ѣ��x���7_h���C[F��.Ů��R�+����z|�_ә�aLwc�iD:�4���	O�oҲ���7��,�S��6���=�WE&��v�ӺF�=TY�q��D�^N;Qv���;�o:�,� ���H�����j��$⭓y���_s�|�Đ�/S��e�Řo�s
;`%ŸDb�Mhd�?����L�fl�F��5C\~�m�?@�~4�E~���ٷ}�[�J.F���E���;EU��q��')�՘Z�r߻�Q�^}v�>vw�VԜFh���6��4ظJ�>�ھ�v�l-���n��`�+���K�l�+E��Uz)�#�3[���_�ٷek��1��f��k��9}�}�~��.�1���'����+���?2�+�E���P�lX;]�rq��ʻ8�xv�Ѹ��U�����Ph�q��g��YF�Df���U��QT�x�*b��ǩ����U$��|Z�o�%>�������g�G��=���!�Y˝z2��J���JF��t��q��m��o���&&���ן�"W#�_���G?�]��V����o����Ks}ʦ�e�,8j Z��&�yU�#�L�����5&���>��,����Fl���:mg��Z$�kxϤ?�iz��_C���V��Ixd��ι�)���ë褳^l�K����P�����H���ҸohL�ٝkᨎ��f�ca?��.��K��\΅�e#���s���e�?�� %�̝��0oA���1m��6`d�1�k���_�<��^���s,C��5���j������d���c�u�3���F�D��c;�P�� �za�4��-�y�R�����KO�w�2�>>aH���b��u:2n��f-T�a�V�Og����^}��,�4Jc9��{Of�[*;Ѵ�z]�H�.톷vY�A!-�Pk����"�^�������0v��ɗN{���d��oY�wz�PP�g]�Fs�]$]�]/��O�#[���Ӗ�3��[��'m���O����w��y��宰���<��{�<ESāa��3�<��+Ki�vߞ�l�1E��f��67�fF���p�,m{h������}��8�N����V�$#���3�ڇu��k$$��Mԟ�����9e��8�8�Nn?I�X�	���2RxJyqg���#��[��zg쀻Fڿ��`�ل�?�d"�q���d v_��ߵ.6��z-�<��1W �joZ}Zy��<����~�{�n8e1�6�K8�{��B�wLՙ2����ޤ�t��e��:e�a��խnO"�r������V����}��
�a�9ӹ\���0a��cH �?Ҹ���π�_��k�Zbv�àK�M��$=�P���}�}l��8��.��v	���������qm�_V�)�^E�|^�4}�7�l�dj���rݓ��uŠ��'��`�E ~y�K�e!�6�o)��G�� b#�\�󔖒$N�w�������%��~:����o{5����>)rm럻�zY=��abW�#?[a������!��+��u�;�7ŭ��s ��ٮ/�.=[���t�C(M�"�D_�]8��i�P\QD��J=,�*�b���B@R�
�2��2�ڏO�̦?0��O������-\�w�c)�ǁ�fGV!�u�h%Y���n��;Mn_ ɧD� h���?`�y���GD}�#*���c-b�C��~���)E��^�6o�گJ�tf�J�^��L%�:>2�5;�>+�X�#���������fw_<�t7��$<�YnB��@�xt2w���>Շ��oWҖ0����࣭����l��F�M6 ��f��Cr"�+���d��P��U%�mme��K'�w7�x,4��ģ��`[sչ�'�d�����+���Wۖs�ʆ(G,�����I<��\�*9j�x+��`Q&�^�P�n��{Kte�n��FV���.z�:>g9��Al�lۀ�nM­�]\�a�:9�P�\�1����չn�%���	���}z�X�19B��M���Ӝ8��'����o%�vp�v�箑��q�j�峱�U���O�+��6,zmH�$AN�nQ,���B���	��z*p�fj�{�ډ�y�D��gL#>/!�L���z��F	���Klĸ���=���8XJ�Oz#�8(�(�E<l�,��z����a�F�Ա��d�Xf~�i<1 {0?�~$9aG� ��2ol��t�}�5w�:�� ˻ƅN�K3e�z�+�5��k)+@�Q�}}��v'}*��F�'����f��,����c����'7�ٞs�������_���O��(�3���2C�-x��|m/��C><Yk�þM�o0Ex�7Hݖiׯ#.�:�j����{L��J.d�IB�Sm�ZP{�9�U�l�P�/�J�xz:�HdMQ4z��	�[�>����K^��P��K/-2�I�q,�1|�0����!�~#yא|�X���&\��φY����t�Ը "��ٴ�y�C��}���?X:�:Z �]���:��(��tf�u�#�<1�z����"j�[��K@,��+����Q��Y��[y�+��k���?ǫ'�l����^�v��,��T���J-�������{3��L� } O׵��&���!�8��-����6Z���ȵ�[]e.߄PN������>��gL9���~��?��/*�$�B��|l���J���DjW�V��
�d���0�V�����ѥ��%����)�f%�e��SX�ѯp����q�?vb'ͽ�I�/�3�ZN���kl}!}D7�v���W��$�AI���tIa���Syi��5G����J3�,�[;X[���(⹚f��l��7��<�8�����x�%���S�hE�w��vc&qm�����o\��3���}�����~���\�P?�0׆��Nw�â���u�&�X����Q%!79qb�=�����ҋt�� <�λg�w����t��h�}�8*O�F���&9_����+f��	�`>����Z;�N��ᤣ 3��j�hI =���h��zk)�����ށ��n+b]�9�tn{��@ȥJ|�+�����(�Y6�:@��*}t��Q�'��h����}��m���I�p�qvs1�-�ڏ�um^P��> �4@�}������w�Ԙ�����d���rj�D�j����d)P	q �B$T���w�9�9@yP_�� ��~��ν<�D���[���2k��̚i�K�˾l�h�>��A<;}�b+��1WA^��;�r�X�~(n9��<'��	-�Z7r5V{HMU�g�c��>���X�����\97�><���>|��4>��C����	����Cun�F��5>���so��:0f���2!��ܷ s� *��z���p�ų�N&Lz����Ĳ�M�!Ad�[ԃ���ԭ�ɫ��)�Z}Btg��c:���X�m��گ����u6l��r�VFwʅ[��'w�O=�+~��%Ε��&���Y�#�f<�C(��k��Zq����eқe(�v���l� ��I����;���؅\ .h�s_� ��A_�J倬X�o�� X��}�VD��eU\��O���=��	�2�*:$>��.(��h�̳��+����YJ�tǛnpjXΉU��y�O8����".P2��q��G	4rS#=W"[�g��'q͞<eSI�e�;Uڔ,s$��c��N��z�[+�K�T�Ɉ-4���G����O�yG��1~O\�u(^��7h�H�*F����UT�F:�\��R�n2�Tf-0��ů�_����/ǱE4g�r?l�8r��hV+����j�Ĕ���^,تl�/ֽL��G��]g��`����ރ$?��6�2Qypk�.ʦ6(|�9i�<a�y6���{�g?YZL��~g;�>�Y�?a�l��%�q��Y�\*��,6H� !t':�����n�-���I���y�g,8w01C�&��@M�Us�Ϟ���Qd\E�`��|U�����g�q+0�T����:�+�`D���YB�񐟧�rTp��-�>�rj����:s8Ճ��J�m��)�_� �jz�Y�z�j�q�f�d3��]�z� y�~�Ky�ک;���ͥN{�3��Exn�=�4�P����ݍ���Ӓ�L�-7q�d��&PU�z��%�!��9S^R)��7!��OlҬ>i��c��/2_�KC�N�m�)��2=��)�7�fg��I����>����Mʧ���L�'i��ن�D��˅��#�-��lv��m�sdm��\[!V�����XHSZʲ<�vo�r<�ݖrBV���� ^o�N�Ug�h��*1�;;D<��`2x��Xv��_����y���z�<�3ʽO�`_l(��<��O풾��g���1d-�*i�A��v��V�oCR��ED�%��Nй����m(�Y��%�x螺lͩ1׏�q\�����ӻ�q���E-����8M��'�
��m�������Ӻ��z鈥�/�+*w��E`��b��P"W��}ҸB��D��&�MSiٝQK���إ{�yF~��p9�y�`�}�u�M�x���H�nf��FN��E$33A2*�~�ͼV���W�S�wњ�墄ʋy
�b.��g�a'�
��F�w25�%M%ִ[�ow��G�7u��?[>�x��uY��n����J���V`��HV$7�<`<A-��XQc����<j'H��w��^!�?��+}���
���x�-!p�+��gs��E��p��G5[ۖ�滋]2F�s��K樨�G�q�����ُ�<Y��^ԥ��3{@M6`�eg��n�C�Zڔ�D�֪k,1Y�	���Whf��]-�uz�^������~Q;��볢�t�+tLO��a��@>@l��"Bd����h��	��]��z�����\mde�7S^�u�R�5��q�i�����9���f��x9�9ta�Q�&�v:/ioqEm���ZwnJӻ,F�v}ޒ,��,N)�J�1b�4Q�;	<�����˝�e���z��ۢt��G׳�͞�D�\�n����6��[��&焇��Z�q[w^�T�CK��m�&|n�(=�E!~=.V#v�K�{2��j�|/�V��z� �{��QO9����'N��B�[yG�QW�0ڦ��G�+�Tȷ��Ql�bu�sV3;ȣ��6�F�9�Ͽ��R���N;ь[���r�T�@!����laI�C���E��=v"`�������'��Ӱ��y-�"�Cƛ����g0޺��Vqq���^vON�r��-h�e�0]����MP]=�6>IA�Rc]�KJ���~f��m[���T-�WF�m��ԥl��_MT�F�J�ʍ���/�x�Y�炋�ϡ�
W�
f�^#(nZ|�x���]]���ӥ��"��>5 �fg3�n�m"�����>J2��w^W& z�O�G�]���;�}�N�=3?μ�+=_*���;|Z�������a⴩�����8|��o=�%UC{����?�k����3!{$��<[�`���Y�w�=i��<r�	�f�u�C�=�j7[��Z��h��(*k���n��~!��r���Y4W�|���]��J�<�dѓr����k�H��Q��^e�s��^ �.	��&���Y��U��X4_��o-L�Сq.ΜjO�%<j���\�x�,�(��%�8�x�i�����1(n������%JO~��JdX�X��u��A4�G��D~(�ɲ�݄��jI0�b�JU4c�_i��&**��V�����_A'��/�Τm�ri�����W�=Z/n0[Pe�Y��UnaLx���"��	��Q�c~�O�11����p��8R�a����oz�d�a�}���o*�c����ծ�2���a�`|�p97�'m�H�֜�+���_˔�}^8���N�A�'��VˢG�Wb=N8�l�Ǝ��o�d����0�5�@�y{���u𔷵�ԍ牝���k��j�c�GЕ$]��:]�/���JkQ�"����)�|��m�i�K�.��R%+q�^⵳��dh�$S/ɤO;��3��f��>��Op{���%�1��G��?&���b�,c L=���bn=��$��.6^K��R�)�? ���>�L�=���R� ޓ2�'��5Ġ����ݔ�6�[���2�A6J�k��o���ч��F}�y7����I{-��N����uM���{��1��&Y�):�?ͅo�p0&�d�������ڢj�~�5xS�S� d�|��	�8G����g��K����p�q�'������NL�O��\����t/�>��>���O4����[/b�6��@��(�骢��>�'��ja�ƷO�ڝĨ�B@�b�Iޛ�(��Ǧ�p��#�����Sb�n���x��tX��ns�g#S	��k\���oHnʆ�#sk2mG�ߤ�d�}�D�)�w�'���b�	SLp܏��YCK�!l�X��//�s���\~r�����-��u�K�!��bQs1����~���v������yt�_p����V?�fm+�>�8Y�k�;��h��s$�)&)2<E�ʹu�����sV�">V���G�-�\�3��o/Z���/�8�񕤳�%䯋�g�z11)@�I,4d�ϊ#�[[����Z�/��i�\Av5��s�en%�۴eI�e�(4��<P7�m}���2�[�L}�����o��IXSZ\��T)�\ׇ�&{2'����ҡ���p\\�#y�R��p+�\���â'KF����B��>+� lx����l2�ٶ0��2�b���K�L]��愸��G�p�6W�{͋�h�Z�X{�z�G�JV�p���44I��p�2Z���4��P�~���|F V�~�xї��b�@��������ԫ���!'B~��x������9��W��L�Ep�בS ��Rx�]i��0��+�&�iq]$�=�Z���,�� ��i�x��rB-��tۤ`9�7�'�^7����ظ�M�K�C��(x�&�%8g�tQ0s���V1T�V�D����$��*�0t�D�'�k�q�d	z���*��O9i����ɒ���li�C�ʬ䠛���-�S�69ș]u|����������m����>d��]����㬁�v�H�@+��jY�<�庳����������u�VhB缭��^�:I9h��h��s���i%i�,���8����;�֘$�쩵���h\i~T���ݩ��p�#}��թ���X�ڮ��\2�4k8=Gyf�c-ͳV�N'� ��SVӑk`�mm�����I;A��b�BcH�p��k��
�!2ɍ�ݦ���k�GƩ8�����=���M�\�hW����Hצ�";��ύ�œM�Z�����6�Q�Ƞ�y�lI��y+�0IwK�k�6A��:+���x�k�m��!������a1ਤ}N���#�aP�9eQ�Wg6�P���u��+%[���^֎r�B���	Z>^pc�Ri��%.�1���]�$��!P���F+<));׍�FD���}�7X�]i�%�,H{��d��z�S����c���*W,s������)І���G����߱�_g��E:R�d����S�!/FD��e�������$.�c��#�����}�s�7k��ਐ]��Wr�/�h6�-�p��y~���8�Q�����j����ut��p$J�0�Z#G�=>�����}KN���g���m�˞�{O���1!�J�F�7�Ds�l�3ʨ�$c1�z9��Yw�Am[��^����r
jǌW�J$�q��A�tހ��tj�!V��������F^�:�q��������Z��)��R��#��Nz��iI�@�6�x�������^�UW��S�Wj��f*����5��!s�h�Eg���hT���ӋK�g+��w�������̅��yJ��^]s��ʆ����l�q��ifj�;�&a�w!��^sM���!�l{R�k���R�lu���s�~�;�?��\/wgn���L:(��?�C��S�����k�p/)�J��V�#�mRt'�y���.S"_���P����=0��Aʱ�<��ʤ���j�t�|>���Z�p�v�u���=�\s"	�ڶ����`����ozj���_��{g�����)R�/LfO�~#v�,s��H/��2&�^4UL�9c�~�n����R~��p�3��p�^��A�⽐eܲʊ�a�r"��g$�:��m	aO~��cc�i��h,u�Y��y\���=#���_F���3����vb�DPN�������S�e���v�A �����
NW�ӧ4Y�9��-
7�b%Z+z���\���~�8�p���U�����r�DL����˲x�N�� �26��i���ŧ,���>���x�)ޯb��:+��Co��_0�y���K����Yţ�J��
i����Q�=�W�����V��O��<���?��6-c����\�,:��ş�}=�9��t��K��Ś%�l�ꕧ�#�:�0��BB�)C�=�ުI�1ok'��l�o�zg���$� ���)���.�m�����BΟ[N�� F��M��c�w�9 >��ڀQ(t�w����UZJr�i��o�)-m$H��bh��:�բˉFÎ�^[����5 �q�ڙT�nx�u+�6������EY��h2L��ݺs�"t��ʛ�3ڷ6S_�)\"�w�*��ĉ�u>��{���[���қ�Id����<p�|Dܔ���g�+<�qmi�]ӧ<]����39�ѭW�c� I�
X�yFt�?����w\�5��Ļn�=�Q��4��?b�� ��S�>��!���>Bi�=k����c�״b����e�w�3�,a����b�qe�`\�t�:8.T@��J$�⸀�J%�O�刞�cL�G�p�ї��
��ܒ4z��CN���5joI^��h�X1\5�K���*h_�B��K��6�����P��/�I��XX�P�W2[������S_^�J�5��=\20까u���<خ�,Pi�Y]n~��9V}W����i���)x�P�LW���0��8< <�K/�U��O~�
��[W̪𧁇�;g�՟�^?��n���z��D2ܲ�(�[ԏC�rţJ���:�eS9��5��*�i�ŋQ"'mY��_�:ߗz���yL�vU�xF*$W�R�y�h�7�]4G��>e���=�f@y��{[�	w���/$2jФZg��R�UR4���+�<I܂2���\�G��
�5 �f��fI��ˋpظ�*�z�'�oO��]!^��$[|��V��n(Q��	�������a�E͈x��?
2e��~xf�塶�v��sT�������r�3׸��%kY���p��	P���S��ğ$O��krw��;G��ړc��²�z}8^�����֣���J�<j$8��e�d��!�O�cI�i�������by�*�;C��$7�L���Z���2�]]j����W��P!�]��Li�,��,��0����k�Q"kg��u�Yc����h���Ȩ�馉?k��Y��,}]n%2�g��y��1<��ށ=��jrsf��%yx���<sH�o��'�ܑ�{$7.��pd�w�K�b'���"����^��k�叀K��?��	D�)�����<�ڥt�V����*I�g�T���5
}�l�w,7N�.��^����xc�P�ӹKiY�i���T�IZ���*��F��h[&��Q�Ŝy�y{��M�/n��WN�/6
^`E�!XJJ�j~�}�.���T��݁��l,0f�̍�oi�7]�U�9�0j4?&~C��c�Ø���Fc`+fl�!�,������;�Ѐ�]��@ 9�
?�_�>d0���A�r��)�L��z�/'���V���<M��H����`��^*�����^���j���#��yE��J�}+z�� R�X<1/O��W�Ƌ���-�[~��`UzeЪʗ����I� '&�N��ZA���?��n�*���8q�dn8������ʧ8\zR"?���Rf�Zr�4C+��`�R |�d�$�����%̱��4���1�&��_�r�k�Oe-z
*W�Ip�9Y�K�]�5��+�7���*��j�g�ŭ���m��Q?��{�����#Le�ӣ�
ԙu6S��3��G���@�hC4���1��4Q�ga�}֮S�b~}��
p
ȩ3���ɐ�1>4g��Sx��6��'y��L��mdR�ߵޑ-oTg���/����c�Pv;�x[��ҹ���Ҳ��T>�IK�`mtzIC}W����D�f2m�������/�Ό��*h���i��>���f���a3�}(�+bk{���9ͪ�*���@�e���r��p.��Q��x!��R�UG6�>�gȌ��K�%9��k���bEI�yY���4�9�'���Y?����s��x���L
�F[��%����T"Un(a�Tg��~�A�{Su��2�U��=�P�q�F]�j��i*����w�����cI�֪�ƶO	�Ue��v[��ĭ���Ju�Fi��4�٬��fg)��xr�sCg�'����'�����xz��ޯO��Z�<{
8��}�ǹm���E��g���o�t2,R��oxd?�R�!�L�n�փ�(����_(�T��(�6�n�m�����
P������0����p׫��T�g��	��@sN�]��/w"&�'�������3[�'������7�YN�կ0��?�9�����;B/E�07���4?�������0�b%=�]�a�pnz(�B����|��y#f,=Yx,�c�{1�/��lJ?��]�J�3�K��V�-� i�G�!��d,D4�?�r沊�2����1ZN�3�O��92ɭ^�В����q��`��/(/>��T��B�Ǻ��}-K�����\���`6�&C�K�H�Sy�u:����ӑG��4����D�ӎ����9��Qv��3B�	:v�2�������7r��FE�룩q�7x�Wy���~�9��$�s�H�H-�i��MI\�t�����beӄ��PAn<w���ty�}�A�V������v4')�~�l��K���}�2�}ڿ��ïؼ)��/�q���
����XM2!����EeS��&���Wr�ThԚ���׀�jP�j3+b˺�W� 	H����/e����ck��χ<��}�N��ıp�pŴ����Ì^�A��a�K�	.�.���m�y��܉�<픓虏�$b�	t���6�p6�1�:�oprZ�j�J5���Vu2����ܡ����ks<�՟��g��g(n�},xK;n^&���6�Yj�-_�&��}6�^���ޞB+>+��]���,�E�80S��_?�p�.���i��9(&Q����Y�~��?�ڢK����FiQ���{�����Ao�6BM��p��A�
�d�4s�v��W1�<J��>t�6����������pO��}�@�GO�����g��C⋾�l-d�qƯ��5�����z�-ˑ+ŗvU�'i���$�L��R2��j�3W�r��^�&޲\G=p:��U|*��������Y�	D�+�D�����#Bt�-P"?�����g�~A|�⠑O�Y�LKǶ�mq�+	 	S6��#̪H^UZ&Ѥ�o�,_�������ƋJBm%���f�. 9g�sH�u�?�������`Ip�W"'q4��ݬD࠯F������3��<c�78<�=�"�~��y��4�x!���fD��>�}���\T�l�趦��t<�e��-�`�ӱ-���I���&��iN���)�@���;Yz�>���}ެצ���tug�����Y���Z�Ȭ���=�g�u����j8��'4]�<������-v{��$�u5��-��%t5��7�[L
M&��w �X�O{>(�W�cf�����63aV��G�+�.6������a�d"m�ˁK1m檾xܞ�;o&1Q,�z56F��7��n�����4���}/�-��|��m~��-���n���n�q�gFHQ{�+�g%������+H�G�y��>�ؽV�j�$S�~I-��Uӹ�P����\�F~�����e�QTI�$�Ř�G[��JK�[=0�i�c��[��?��Tɏ���^�%
���@z�O���]ݥ�/�e!g�8�mȠ�X����)�zaP�Gɱ�g���8��uŪ�[�H[���U�d2��c&=c�h�W�prfP�}����װ	�0���6��~x|$����֯O�]��H'�1��>����`<|��	��q��g�CUۮ#�U��W������y��ᴩ�Co#�o�(,v�U�����l	۵��c{�Vp�nΑ�i�k�_#�p8�$�y;�ؒ�J��^�x;;�J��6b[σZ�ۮHW����I���Z��,�eT�a�����zh�%�o������O��]����:���_�y�d�.��U17�%�!bHg�$���F�+���h_�m~0��ب��/�����b��*
t��g"G�!��vM�t�EDY��8C���ߙO��e���,ﾓ&@��4΂U�F-Rg�u�R%4=-�"���0W5�*�� �n����ԩsss�M� ��x<�x����8Ki�y��u�i
<��������p��w�����Ճ�
vƢ��ZA#��"� �Ѐ1j�Oѽ9W�&��U��l�U:ȵ)\F	�]�푁ʮ��Zi]b�f��&B���\BE��K�O_�l ]-�P��iø��Z� ~ޫf����Q |����{O�r����6W������[���>�E�f���4����9N����f�������4`6���)|���4m�5f}�T��ue���0ηy���
s�/P�"�(�5�'@��l̞��^u��Yz��>H2k�$�rx 0��ޤ)E�H�l��Q* ��f��П�~D�É��U���zp?���Q��y4%�Nr,�6��������x�i�K�[Ļ]Q�DX�&�h"enyU��L;�^[���f��R�@me������)4M��?�����KP���Mr�B�=p;���s����h�A�S���[���i�J�X!LWVW����L$����ݧ�D)"L}�z"��l<Ce]�u�E�wù�l�7����Aj��*>����hb>3my������5L��E`&[3=��g��<7�5r�U�+٢�?�[�p{��+=��)<�G�|!�XU��WY�X���*>��_��)��a]F����gzS���/��~�,����\[e�;��x�_��q)��sW�E��I�-6-�]�4�F�����`z�2�~.*��@�}bׄ&TEC��&��:=B!*��tO��6�8��߰���Q��-��6�K�?$��,1&گx%3;#�?��ê�a�KlD�#r����=�[Iɚ���=�,�T��

���r֏KU��/.d2�����f����QYu���J��/�O
	zj�z�$2za��K�NTΒ�d%L�E���s�i'U>z<z$��͹����Q�c���9���Q�s ��鳱lmFN��[G.R\��x�Z�����Ĩ��%��ǋ&�b�׿���'�)��;�>)���	P��#J�r�e��#�r��x?"���_�Y�(�$�3����jE�[��e��l`Y$c	���G��2��`J��=PBrq�Z؂�2�6����0/�#��r	v�_��@@y��9�� ezUh�0��_CY�sf�.�u�D	�E�|�/o���_'n�#4~x���.��gZu��]W)����B��(]H����{�m�n��mO�{�����K�C�Uw��/z�H*�s�sX�՘�����VYx�r�'��i�0���2Lli�1�VZI�a2uWu(��P!�	c�3����$��S"��̇�>�����Y��)̟{�Ie�9o��=⵪���G8�j}6�FQP"�%A%r9aV�mJ�b`�5�F�nf�5p��-���G��J�ړ�R�k�"�i\θ>\5���AQ��g�gP��|f���$��y<J�a����4�A��s�kWv�H_�T������^�tj�%����F%W��=���'� �f��`D�%7�g��w���1O푢�pu	�W�x��]"�~�����\K�pb���.���>0�|Z��Wr���P��~���d��z��j��!s]n��DP���K9�x��&��N�w��O�����\Ό��$���R�v���g��&�'[��y�.�y��ѶV
�=��@�M�U�-��|m"�q�d�� ��	]��n��e�/�W+�/d.;�I��bS �O[~D��U�!E�=H 7������/yv<��	�S�k�Q�7�Q��wv��SBt�e:91�sm����݉��0�"��ݝ�{7�<NȘk�dL��g&�\��丅�� �2_<9a���Ǳ;�a�e�'�P9ͬ�A�$��¡��"4Zf��\ :[�r	�qm���	��4+��K��2�f���lkl�Y��^!䤽B|��|e��b��牦�0�᜾ɓcζ�.�)ѯ���U�5��7�@�`0T�)/-�ަrz����O�{��r2خ�S����g����}sDU��r��d0ӟ]ª�\~2�9tTlŉʃ3'墼�FN����y��2vUo=��Ir�Su>�r}x��J�	��J���"�h"+�����hvG[pP?� ��ͽL����R�@�4ؘ mD��
��xf%�5$�<�M�7��	�� �pbf�c������ �ov���G20XPsZ�������)���)�U���U����o8��г�P.)xA�N8@AȤ�_�#���*��u�'(13/�9�J�W"������L�
�y�\�����<a�2�Bi�� .Td��r"�L��)԰�_ǒ񹂌�=�{"2>/M�k�\>����_ɸ����î�����t�^����s�r£y�_��#���j��:~&��$M�h��NmZc5���F����2/^���-���ᾬ`+���0�
>��q��Z���/�xE�*m�A�(VؠCx|TB�Za'�A�(�*=j��_~M :������T�Va7�I%���i8�����	�,a��\	ȂC��Ǜ�N�dB �U�T�:_��zٟ9��y��K'ʚm$�%�ɮ�*��EQ�4��QB���\�J��k^�M^N\�cj��Z��%*�б�Lf==�,%��ABt�SZ���͑8OD�R;����0T-lc��V��%����_����+5C�e@h�%���ʚp}�>�8��j�Q'N��j/�����$J+iL+q��1໑�;Cx6�@x~f���3�͉7Ĵ��#s�勥<�K��tow�����H���=���z�d*2�"�����]�C�#�͝G��o��=�����[��$��;�t1�:��X���� ��"�Ã��.�c���HA� S�M�8�*"�ِk4��G��[�WXF��.�A9���܁Z�O;,<����
�)��X����O&x���y H
������W�&�b�g`r�bQ �i��#_�AL���<t����CN���z�m4�_�,��e+���K�}c���c�6���خ��%~����܈��N�Um�� ���Y܁$���E��G���.�G��H���6a�����YN�����s�fG�4{�/&�Ī9�b������T���_�
������0n�(�8�����H�����,sک�]��S8l婇�{�D>��+7A���S��o�I!�Cg���N�\���_�s�pR�.����״���t$PrdK�ȇ�L��h�������fч=fuS�B8�!7��Z9�!dB�T�Bx��b��W���"�@^�E7��f�WO�$_���K�K�w�/�<�a��O�j�vph��^�_0��*���j�^D��m	uk�ǟ=�`�g /h�|���#�BM��s_��L&z�x��t�y>��B���Vډ �}J�V{kb��A��)��Mp�� �R_{��=�� �|.@�ZTs�"����^�.uƽ>!�����^k�V��fm�U����5��1lϰ�ڎP��t#���a�W�Y9�wx�C݅sP^���kA���c9.��uݝ|�e�CL�I�$��o�8L�����;E�wԊ����]p���fpD2[���gk�6%�&�j	 J����#�p�x9��M��?Zi�nv���Ux���7�Fr�����hJ%rJ����\|/0K�˦I����9�K��@��M��;+%NbH�Z�U�%Im�f�������b>��N2Z��\M�{��E���T�[�:�c���)Qfr�#����/��{w&Q�gj�����\��gQV�v��u�f?hE���|JD��N�Q�	s��ejiYr��M��2SF��h�^~�y��������H޸;�[�;�����<�N�i1�i��m�v8/�9�?�M=���6��w�f �ک�vDۚ��g��X��z�Q����L�����)Dnt6���b�ؿ�Ń�ο���͢�_�6�����U��>p=*��qr��ϴ99���۟��l���O&�ۯD/F�����V�I��tܨ=�<?\�-��������1\���F<*�I��K��r�G��Dܻh@�;a��H����6�@6�6K|��?n|�ylu!���%,��~z����z���n������}�=0Ls> �B�K�
�?������Ԏ=T:���_���ˡ{��=�fB&��;�]\�H
 A������s�̧��z��Q�۪���ßԷ$?�V#V�5�p�����Ш{��j;Ex1]����)$���W��8���ֽ_��up���x��AX]�Ͷu�^�������E㳃#�R�㳕@7F(��m){o"��Bg�?���i}�%-��F0H���l�;x������H�ZHR5�� �kioH�2cr�Zݸ��&4�q�۴�Mn��Fh|�.�q/#�����d���׼�U��}q,�Z��JFbb�_#MX�H�n>j氷�ǖ������X�/���=���lwJp�:W.�<���6籌
)4�_N��0��W�Z8<�x�|�%�<Z���b@��ݿ�OiKs؄N��R��o�L|84�s�NF�\���>��"E<��#�ыp�sh��p��xW`D̗�y�w�5o���\5�gėʌj�ћ��Q��˲�,q�C�NV�EvN�O�h��:_�;��Z	�~��;�����s0om����(>��cu�j�V�2Ar'��.��c��C�+����ӥ_Q�4�@�p��yFj�`
\ZN�{�2�א�K�	z)�^��o�~C?���8��f�N�̏���T.e�O.[9�cx��|D*�����MN=�$q�б	�pk�gӿ{�PC��H�Hr ��mY_*�e�%�,�� ��I�j:%^�&�}����x(o.�l�6"��
���s�ۛ2�Q�9�Ϫy����,��?%�fD���Hs�O��(ԏ�ĪEq��<U��縖�l�~�QoJH7VR#��GS����ո�U��"u'&���
��-PIC�:`k��9��L=z��
j4Ow��2��N�V�}�����H��䰠�	�X<�p��Xa�z"e��+�Y߂uw��C;V|���Y���[h���]0�����t�2"��ߥ��M"�N��H)�-z	�uw�U��C���dV���#w[{"�{S�O�
e^�!��UX�.p�)͎���6�M-�/&����0Srk}��,j$�Rr�b	t���8g���`��;8uP�|��� �̦~����3�����l��ԟx�̢W83_����b<�y�qs�E�7ST��p!\����b%{�w
^�������7Ӥ��.E�l.Q1y���a��.Nk�i/qoCQ;���ᯡ�7q}wbC`�Uk9�@�L�V�rڏ]BH���+� �R�u�SC�
�7'�!�L��$�vdg FdW���|��:W^�dw�?�TǁO�mv�;�a�~BB=����ͤ̿6T��!ׄ�9����� �ۏ����d����="�� �J#����?�!	�N�ȝ�_5>ceM��-A~r��#W9��5�-���<��w`h|(���j��Z6�F�/>���������|2�Kt����n�8��P�)8%ތqb�	B�B���9�9�;H��Ne"G�8{����7�?���w��=����/EDzjS;n�n�_�;e���e�x�_C�c��9��'p1x!���#BXv����������ᖽ�����2QZ	���AQ	��ۘ�.���1p5�\� ���B�m������&�|�ri�'i6�����d�'{��8;>T�/�sI�A�\��{�:'�A���u��s𐉯a���]Md̎n�}��Ίoi�}��0�HEC5�I��5|��r�u��5��@��T�;��x|Pt��z��h�m6�F�n������~/hM^ ���)�ea�̋�� e��6�+�ק��	���	�g�����ɲ�g@2oL�/k�f�`�SW�٬���w��-P�I�>ݽ[s>B�N*����9������+��P� -Ew���O�_o����m\eB�g��ٵ{EcޟF|%0"�y�!���p�ڪP�ߤ����<�#�1O3q�ޤy�t�I�4�Oi��C択����H����N�+xɇ{F*QM���ĐBf��䍨r������&���>Q�RdT`���`_zD4�ϗ̎l���w�wSwƫ��:ͼ����f�j4B[_e� �䇖��6]t{�Dӵ���3���m!�+
��B��g��C�,���>�KY��T%r��>�'�KN�F/q�d:+'��񋎭�������D����:��V��x�/k�y��6�X�����dI���(<eVZ+�Ox�'��|��ik�M��6���j���ȍ�2:���>�\?	�fN�!`$����#mfQ,�A��� i	|��=��4�T�a#E�H��@�=p���Ub	��6�՜�J����T\:���j9����%}�'GR���T�&~џ��L�B��~�r��	�^6Q�4��`�cl�eQ���UeҤ/�D��� �t�q�~O`��WOS�Np$�ao3u�yD�kjW�M�������[�5�<A1g��<�$P ��a�cՏm�'-;֟ʄ�E�/�����H6�D֣x�Gy�y"Ey���\���*�.�ۂd��>��ac%�tmF	1�q���M�qK��E������L�H\Z�V��jR�M���l�ʈ�N�X~�?w��w3v/��K��ơ]g���-��<JD#�4�8�� ���,(s�vw~*,Ѱ����K��#���V-[腭uodgp���E�=)���XEb�3y��_v�
h0'�j��x���0���?Am���c1�4�-���;�ש��eġ����a�|FM��&�7D��%���M��>���B����ss�?K���'dt�+Vͤ=��~%򡙍 76@J���KH�s-��/��� @�����C���?�Y~l�H�!1`�9�ۚǹw��|pb���์(r]?���l�(C�`T���o��H������LYƕU^��/R_S��safL���3�
�{_ŖFvjE���qf�.��D�ȃ�,���]�&�3Md�#�%�4or�*S)�uRa�lUn�'d�=�2'�	j�.��v���t$��?�c?$��X&V65;�O�բ2��&Q7�����G���0�<Е�§D��D*�*���L|F�Y�?���B[�t3�.�e������ҽ--���+G�����{���KĎ)�I�����$6>�si4�d��em�ૐ��6|�2Ϊ��M�f.I�
�D�����Q���_��i�P>���Z�r����A��ݴ���>淼�%�;�8))�JXh����I؟a��*}��ʉ����F>
9�k�	����#�gt�S��T�B|J�+�+��lU"k�Ѕ���i�t<R�m1*d\2��Y�d4ܱ�_TI�e�,H��'�2�k/�0~P���X�}\^�n��%���O2�d����&��S�E��Z�����|����ny���'|M��ʥ���>���#r�	-�ѯ���m]��A�F�/���D���d�����[mk��>�X�l����s/�6���wJ���#04�ն���,z�8\*:��O�7Ľ|�
�!6��a# "��{|��`��h^�ߺ�~[`�6���k��:	ɪ�2�@�Ͻ�Y��3x�9�>�b�����I������8��}�˧�oO������l�D7��v&��Ҁ�� ����(VN��㰴&�}kY��W"\m��la؅����_�:�X�z�~v�-0�5F>~<�O]��Q8ȘE���)0<��r�{�4,T}+�ܠ-����=g#��\�fӜQHr��#�X޲�Zh��YC^.K�S_�K�j`Ġ��m,m�[C�AV�����+����F�l�as\=N�s��c�\��MǔqO�qߑT��r������|���]��	-A*m{&}� ��=��������O8�}h�Na���v���:�~	����Ӛc�`Y��C��g/�s�'`g�?���p��>_C�wB��~	��lG����}y>Ic}�L�a�}�����N��BbY��`��ja��2>��"q��~T�//�O[� S�����U���������	x=_����_�4��6���?G�N�nj�-��\m��%������X��	���w��6[����\#-}{[AKp9�/�X�W�e.'�e.ƗոǗ�����%����ҏK�C���#cʾ�X��@�<c�>O}�=����#�hq�b���c�ҴJ༎vBhc������2�lzm`}���M�
�>�:��bY~<��CL�=�]Ӎ��FO��ęvrk��:@�})Wj�t��w�ф��gH�u���"3
�
������4������8�Ƀxx�E�4��E���m`�B}���c�����t�ֆj��Qp���9����h� c� ���ӥ<���+X�!8��/�4�L�W�će�CD��OΟ��q@a�l�jQ?G'mg1�&��Kuo2o�;���aF���C��;�~x2`K���4,��LZ��4#稟�t��vc	�Ԫ%%��z�$^Ɋ^8�=�fO�'��9�:K�/\~S]�$�Q��� yv�*>{L�q�D��-h�I�-j'_�|+\�$�|j��^��ӽN�)���셉�Ա�v��5+�=$6٣"Df�j6b�Q�����4����"�c��(�2�=�0�|TbSk����J�,d��}�K��@k>-R,�1�~��g��K:��!+����f���Z����ZO4p�&����t��,���C�C��]�3_i�_I#*�IXy�}ĵK���(�}g��:��D:��\%�
]D��(����X%�$]���oU�7`?7�Hv���]B�܊���X%r��I�Fx#�F!o�"�q[t��d���C*<\�79�� /ԈZ�Z����j1����}q9Tb�2�K���[�Jp�ME�q��v_�n������X�؃��UHo��hY�0,�k(l^��M5��֙���]�����z����i�1-Jk��;=nw}�oEX�5&}v1�����|JO?�ɂ�Ժ����� �� �	����И��d��0AKamx�HJ@�4"�rݦȶ�������դ�{hC";9~=�[~e�Hh����ܡ,q�����U:0Nu����]f�mZV$�KKd��L@yU�w"C\�{�k�4��X���h�hl�&�-�)աD��G��x�Vu���8%R�m�402q:�]<f�dV�Ew�W�p�]�jK,�dϴZs?������	�R�
�/\iQ��b��d@P�j�M���~p��u�-�W@�c���q�����-5PÇ��K�$�*�н	f����[�9�YH�=,�h���[@ϡ�}F�ܩć�y�缂�����Bs�Y�ԡ�l|x���0C��uyQڗv&F	�����K�<>ËO�F�p���r*|gLV}#��㬚�{'���t�Dқ�p�	q�%����Z!��yGڸ��%F���q�N�B;Y��Q7�y	8��㈌�jf��^f���\�c�4�:�<ͬ��t��-��S�M�;����o��*5��Y<�׽ߘo��ʘ`QX-b��rFHQ��N	���K�4J��)��k<f�f�=�W�X;.�-/��k��/�T2M��APbL���E�@�pZ}8�x�4e<*�x}\m�u5����T"aQ�Yg�`21�Xٖ��φ��Jt*��YJ�2#�?��B8���� ي�[�v�ۑh�����4+Q]P�F�[���m ��Ǜ~eA� �<3^+��,J��j���n��D�Nt[�Bo�5�Rs���Zjg[���f ~��v�x�|$Jd_!���cs�f��Q�F&ōMK�j��n�=�Sb3��2���K��=)��ɂ�n *e=�D�FC� ȉ�h�_l�Q1� #%Z.p��$D��J����uŀ7}�s�6~D����Q�FӠ�7��E�F.��ny��&�Q��U��40�D�~�Yʸ�<v���C-�5f;��Vi��Z�>��}P�+p�D� ��_n�.~=�EԨ�v�M	�g��n� 9J��_a����J�&���pJF��E�w��#�`���}Ge�ޑ�j���b��x)'�VK����y]@�ɺJ��MgՄ0�|0�ݷ���1��ba��S�'+wJ���7��RF� x:�B?CMC֢�x2ٙ<I����(O|"*Қ��t�U)�X��"�KD[;=6S�
�n~$lI<|�����8�ÅW�86�ar�o=U��Ne{K��ͲH��:yH��%���4����]����kCc�2w0�)�n��1k(V6q;D�ص�C}�����*��<�S����ݿa�r�cz��d�M���4������K�o�E�K,�$�!%[ә������NB����;'6"��5��dݶ,��e�۞ӛ�����y=�Q�mq�����H���MlI<Fk$��Ў��00��J�:�R��+����hE���A���}�\1#W��f�*
^��B�����!�)�/�(��<�a���K>�����A]b�$�.�̼E�Lܾg>��S��[R�<�T�bG�0~�f�ܻ�I�a��������	�{\��^K�~LVJ���EJ��)s���m�Qb.�����6�]~�:ŮM��^$�WDh�D�v��b$X|CY{�l�R�2"�-���e !��8���(�R�)BIp��Ǧ���iSm�d�K4+O�nW���gȒ �����=1��h��C�#���	��\�z���
vEwG$O��Y?h���v�E~)v �����,i���{3 ��%�-�R��\�j�u6�Ʈ�h�jl��ri�w!�u6����;���[���a��_H~nt�;��~⥣\`#�A?�f�]b�Ȓ�8�~ޗ���`˴�tUOW���fI��M+��\����"��M �U���}��F�=�I�=�2�@�S`��'
S�}$�Ƨӝ�T�W���_z �7d(�}��׷�V��ڔB��@���<s�����'s�[��>9]���3���4+����a6�%�[׻��1���nx�+����
�˩�R��&W��/ev�2�f Z��ֲ4���7!���n뤷Gқ
ov�]��i5U/B&�AL���R�V�j�z��ޔ�[�z}���-3շ8�*�J}�	&&f��&�l�F�S?��������Z�ģ�լ�Ɣj�W���=`;$Nټ��h)}�D�!HM����/A�pC�A^�� 1簾���^,��P�ɳ�o��"�O������ˁw����"��'_E���4v�6ŧ^cRw�"?n�Y̮*䘿/ޱ�,d@���tr85jL����[U�;��{}b'P U��cq�>*7p=vw��[0�N�u�o�x�K���X�ˌ*��B�u�$��?��.���g��?�.?�L�A͵�@b���X�]��-�*-������$=���1�ˣ����ԃ���X:��'��(R�]�Or��ꄬ�K�V��3�=p�~��Ͳ��������~ľ��r݇�����Y�	Ѷ�e��a~9��&�i�~�4x:qoK�AQwPg$�8�oC��Kү~T�4��,�6���Dw7_����)Q�h�%/�_�\�7���~Ξ]9�]�̞.��m��!,Ox2�]X����)f*m˯a��S����P���Ŭg�Ǵ��-��G9c�xH�lⶔQ/UME��Sq��΢p�v��Z�,jT9��I�/,C�����ʜ����i�>u�c�IZ�u�:��9�?b�M���8@&��4<��cig|�д����5'�8:���{�sHHW+p��@V=u�����d��AՆ���B5��6���/Բ:KρM*/ܓ�D��U�`�{H�>$_���`���dv7%a��i��H�ICD�)�NZQZ����r�j

�^cE����d�Q�!��������lZ&�2��FmL��ӛ��Vf�����5����f�U�NOI�#2��L�h�v�]��p���v\�A�K���9���&��BmbWq��< ��U}�=w�F��L9
}kޫ~����\��7��Z��D�N#m�s	i]�&;���A�(��zK���W�~�?'�s��f���0"�68|�pB�ה�`6����<�@�4[E���|2B�9���D'�
��T�nW��������\u;�Zb^J�U8�5�u<�%}j��M�z]�:9sG����˗�:B�瘔ȁ,��,����Z�j��X%��u�}�J+���������w
u|w`�L�},�y7��jr���3��(O�P��e~�
���?�4$�cZ�N���J�sG�� ����y` 5h�R���вsMb�J�0"��="wp/|�v�ÅKFh�8:[�_0L8��w�(#*|J,c�l���3f��-A��ӛhV��j�M�=8��V��7��ȥ�K���f�{�}�D1��/�=�j?1�S�����fZ
%z�E�b��NZ�)کD��yYPU��d�V�KT(�rԺ8,�:�)cMn듛I�b=qm�<GD؊����KJ4��k�d��z����~4v�^���"�zX=�����AnK�)�Z��l�d��	l/�M6���`��3!(��(O?Zd� ̿��k���^��u�2m�7x�����&���ѭ�����o�~>-Gf�j��w"}Z�K˿fbn�,Dy-� 1�2��]ZM����p;��5���·�Y�ݩ����a1��T�;0i���?zeTS���"�tD�Z��z����'�y?:�ʺQlr��pC,��G�B!b�!9��Ec>|r^1�e�?Q�'[�y�C-&iQ����?��������ce�}�lu<�%0z<�?�~V� :9��-�萴R�ճ�Z����j�vq5�q$ۜQ�&�l����T���@��-��C���^1���Q�L=7�2L�Ɣ�\��	�#(kQ��^��e��,�9�8��Z�=8�%��,��&H��ŗkEx ��(K|_����gd�V�S��E�2�U,�k�˗�Ep�|�V�_7�6��j���v���;}c~��R��H	��/Cb����H��;ѳ�񣀄��A��_����թ�L��2�Ȣ�-r\y�Q:(�F�K�9��w}�:�w��
�����{�2c5"�y%\�'xV�l�8k�Op٤�Z��y����Z�0��%l%��Z�'V�9��m��Ҫ̗��Y�5�X)��wkv��:B���Q2�dxS62���A;)�-��d����ԧD���8��Q�X�@����h�z�_����8~C�=�C{Y$)�����kjQ�w* �~�B��8�ٗ�I�k�����$ޕ�f��{�	�W�M߯�;��G�h^��$cǢ~�>�)	=�p���U]i��f�%��;|�D~���U�s��Gij�6^�L �>��0"��Tq�|�36�li� 6r9u~�Z�P�N�17��f�(���{�����51τ�����
g(a��%��ʀ=E�˰�o[�o�?P����<�d�׷i�V����5��#*�e^�K�/ԟ�K��Ga`�&5��}d�������).tFk�eG���d�گ5#�/,@+�.�&�M�ּ�q�(���N/��}�p_�g�b�,wu�B��ǰ˗�OY���0�㕥�ح�����V3�~�wVV��fxmŽ�H��M/���a���:y����7^`�q�c��.�b_�������4PHjP|�'`W�V�j�G�S�u��Z�-�6���!A ��<�z����H�y�isr��.�K�H����|�Rn�S"��)�G��O�B�O��X�.��;�z�-�8��`� a�NM�e�h:�����+O�"ע������9�N$�/,�Q��K��٭D�21��
�f��S��Ë�ѯ*g�[��=�6l��{f�Ӂ�C^�6�Hs���(R�q��(�\%��5$//"���dj�F@��k�Ѳ'�Qn��_��G4�-�vl�	�/|X�M�� *��8�䟴Q�A��1~ί�?cW�L��\&T��q�~{_�/w���o�Wd<Hug�D�ۭȆ�x�o�T�Z��4Ğ|$��V2dK��o3��� ���zr+'��Ud"8��*r��H������K]����DR���:b&}Du_j�f@���V)�1H_x�Y���}���=|�[�a
;-	���A��nc���eq����8�>�ـ��of��*=|mƁ��'��{�bg{������Uگl�s��׈��=~����7�kq����*�Z�_�5Z�<{�x��k!=�'��f.�U"nb�t[�AR#��x�k��PPb���S2��_PR���3D�ACN�g�YCr�9WO� �g�Km�fs/�=m1g�	H�������x��N����X֔z��2��R����O�e�6�yT,m�8d���{�~��!��
�~�ik���J$�;>+k	X�߲����� ��5�j�O�K+���2�	��#����I���`���~eE�I�D�0Q�d#TV ]��Q&q�s1j�|�T_iӟ^�-I����[�8Nth�5׎P'�C�T���Sa��AL��4��J�W�f�hs�H�tD��?6m�M�����>n�-��jV���y���W|cJկ�4���z���^m�����oE��i�\���֣�H�X=��DZ��2P>qAJv���V��p��ȁ�W��R�ؤSf��ā��snRu�R����R�Մ�l�F����g���5ݧfŬ�AI��G�֨%��-�Y�%4������7Åߊ\�+ZQ��E��pP{��n��|���fՖ�y>�rb��I%�)�V�������y�v*�C	I9ǂ��+ؑ��p}�!1[%�֛�Yr9�K�p�ǽ6�IJ���?P��\�*�t��C�X��(�y]KcA�4݋|����J��Fwӏ��p�ۏ�Ӊ�	8hkd7�M�M�f,ԅB��i�3K,F�U梷�N=��ݍ�I�P���J�w���`=�犛"&�U�/�_y�d��>TV�z�Y�����Qo�¼��F2O����p��D̍��B��+ڔ��!��ں7;Ђ|�� �$4#��lo��R�2�8�N�6��%c�;�A�kH��=�h{��b�Cm����}ǡ翞��+GT�fS���#��x� @������r��1A�Q5��{N�E��fU"[kĴ�U���W�[����Ɵ��Kc�a��Bp��JGӥ'&�T�ħ�OϪ��p��~��E�b�=J�S?c�f"zJ�%�r��;��!��.}̴��ğ��j��ء>�"Ub��I�Fׂ��r�Y[fUʅ����Z�A�P�Dw���N����V�[�#�W�b��TC�W?����8���j�^#�����vL���暷����Z��N��}���������$�g��;������N~Y����r���`���߼�R�Z█>�LZ7u{@N?Ă΄�hT�4����D@���6mz�IT���>�Z:�+Y��o-�-|Ȑ&C��f��w���S��z�H�����t�ӌ� OU��D��u-+G�T^(E��3���n �~�������M8��|�YKֹ��ğ�ڤl�UO�V��Qk(Q�W�S���طI!��"���u�Rѩz���7��WV��A�[�s�^�֐���T�|�k�A��l����QK��E$�'P�M$����^K�lRVw�4���x����E���8|j�{E����ô���*%���&�%|"��� p춟p7/�M#cp��j��X�VY������ʚ17a�m�8^��F��$��9��j�d82�w�r���U\*+O���V�GՉ8��wnZ��X�x���'��j�g��;�8ZLSzGY���n�C6YL���ӝ��3���?�N�X���KXʭ!hwx�D8>��9��Z����>�J��JLE�8Iʑ�)QlŽ�T��&~��l������=���N�b��e��cך�Ww�]�abz���G���ʩd�ߦ�{0O��!E����$@�&W�J�@��@uR�<�e��@��5�B�Ik}��E#�9�p�!O{����3
���5k����p�[�����Da�� *<�.��Vmht��1�5���&I待���3Q��S��P��Cm�Y�ɃQ�^u���ٖ��4�y'QoJ�3�7T���w�Yn�p��E������5wT�k^8�|�9�a��6�����SkO�ؖU_�q0i��<��*������Cj1A�>nV{��l�1g��{�~ꆨ�_�Ɋ5�K�u<�����[G}����A³���1}�;�;ז�P�U�r�E�������9^9M,�>��Bt7謲�g}�~��^�`�W�G���:FR�`>�\��j��`s�����԰��Ɠ}��t����	����ǉ��k��L�qc$�ݤ?��cs$ ���
Q�����N��C�+#� �p%�NJ�V3־��x�17j-�<a؅���̿�c�f/b�T�U#�&�1W���/N��F��m�me�����hS��I�,m��-����=�NDT��X�����9-��� ���l_�m�OuV�1�+��K�����i�{茉�oZ8DU��#,���|R���u�ơ�=�t�D�rx�U_�H	��Ncg�5̙ݭ�Ԏ4Aw0-�ͧ��j�w���3]��^BP����rZ%%⿜��߱f��_
诬�x�6*zaۗv�mx�{ɧ�f��{���z���%�$`�m�^R�ͥ`S�^�y�=� ��C�	�b?Y�c��\�T�@:"���f�\�D���.W�Zk2�\�D�C�<�u%R@-�o��Y�?ub��H���T ����m��.�I2RU���������Ç��;=���ڡ0F����cK���w�v�s@�����$�n���k�hՎ��f��_Ҫ��-�0{����*0I�{�)b�����^�V��Y���d�ڃ�dxп.W��r<ܛlĒWO�+����u����,�����j��PV����Q�H�T;b&&�z��,���;ဥ�Øe��^(�b7spknu��M�+��LY�R��)��L����e�����)�G���A|��Yn́���K/�w�Y%��;a��C]� z����I�C%jl�PǦ�]�i#9�MTM
��s�I-:�l&�����YaN��
:!{�ׯ�~} �J�y8c�$L��M��ֻ	��i��3���	���da#E��	y��m��B>�	air9�W�L�d�fH����/MVv�%����M���{�<_	+�i����z�������v���$�hE�|�֜���s�((�^Z��b�z���P�Sk�M\Z����[�B{0�m+9OQ����S$�f�7��S+�-�X�,�v���5�&�~*)r��lZ�J���3���D��7�?��UI���3���I�����+��++�!���?�m���V��W��gU�ҁ�5��q楒X@퍓�$4�E��[8���V�=b�I�{�T/�S���+��5��-���� ��۸��"4�� �����rp�l��)�\����K`��Y��7�e*��~��5x�6%r	��O�A�v	ڈX�ϟ�_�ʪ��{}���]���3q��G&)����d����g�[�?^�/z��@]Z(�>�X�Ud�S�	�GG�brt�O��aj���ޓ��ᱴ�!�̽OH��-�(�lu��F_y�X�����o�E k'�� ���X;��ԩO)<��;Ƭ҆����e�	�v`�~���ӿq�B�/I��ԌV��$�k������ߦ]͢�	���H�t>|)�S�e��\��D&��66�Ͷ�h[=q�E�Z�!�|��eW�����ȋca�pw�=�sD=b�Zu)ko�Ȅ@K|e����	��[�����g x	���J0�TLuc����l�|��x!t5i�=�@U֍�³w��z�D�v)G���A;�!c;`�j�֯��X��ִ��$�G��a��]�� ��7h��h��H+x���KQd�~d"	�r��sfi�DȢ@b�M��R�ז��w�(����Q�*R7	�ا�Wj�����uj��&ub�:=��Q�gh�6VHq����^��#ln'����R�������	ާأ�K�~��ia��
q0W&�b]�Sji��Њj�v^���÷+��E?���"֓0M������[��f�=�^8��P�� 66�Xh���bD�B�/�㗠z��#Wor�M��6����`C8I`��LT��$��ٱᛣ���<�MB�O�d��^NP��н�94t��Eb���pg�ك�O=�n!�A04Z�9e� R7��%��JT\�"G VV	X�s$��/��?զ�Jd�d8���M��[��)}ⴈ�¥���H���/���C�kkLj=��C��3f�:�*��R�>�����g���Ɂ��Ԋ"%��/S)s����6����l��l���������\����cPɾ�Ri�'��P�V� ��b���@+��rU��Rsx��Ĭ��-���S�k����\�ޖp�wƬDX�	�n�;����P3�w�v�d�خ<ݮZ�Q���w(�tJ�{MM')k�JS�~�j���R�~�k�v��2`�B}��(�2���=P�϶���{��]�~�B����{|�M��I�:�%�D�v��bz��G��4��6�k��y�g�M��V�	Ps2$�Ư��3I���P����ޟ8�I? S��Ӕ��E�+߈��|s�-Tu�0��ܗ���8�s��U��'!.�PMQܺR�s��_��TU�9/�`E�扁�Av<�3O&ң���?ź�������2y��B�p��Ԙ	{�g;w0~���6̓��?b桹�C����o���'Q�!RK+`v�ĘxI�E5����Z�%�u����`K�^�Q�D��*��*��bS���9���e��5g$b��U�M!hQ*�1g!{@&}������넸���\�XS3� P�!�'z9��8Fg�y�z4� d����f)�
\N�0F�,�#�%ܛ
��l��ی�b�j��9�Va=�^	~�v1��%���MH��n#S'�Ƽ9�tAD$�$���;"y�e�گ\���Pp�hS�,Nf�Dϝ sޛ�V���%{S��Y�ـ�DŹW@X}+����i�cC�����J�H�� ����%`O�3�w��b�C�L7W�Ux��݆4��X`���y��Xn�� ?42#�h+4d�p��#��5/uKB�4�m@R%HI���	�)�3�\ِ��\ [Ą�e�%c��d�.vj �.0T�r�	�I$��'��}~�PD�%-�e��JR;B��L�;�qȹ�?�685���:�����Ꙏ���W]���?\��
��g��?�=������k�oe��WX�"�hՖX�}eN_*�<������S;rXҮJ${%�W�E��b��g$�s`� �0��cWZg�#;�'�Aw�h����P#��a(1������>=k�g�3D"?Wix�Ƙ�?���dռU��)����^�ُ�H��`�o	_ܫ��|�߶ز�o�F��ɄgwJ���}����|�����k'�`�%p��c���V�-/��t��<��;+9K�����3���(�I��5# _ݺ������2p�������]���AƩŜr�)�s�jws"���ĝ9�p���M��A`h�#_�2�&���>����q�HL�!��F���eN��{`�(�D���V��P���HTuj���O����_��_��L�+�$,��O�����1���\� ;�>U_ײ���ŝ��T��ߏ��5&�9Ƙ�,A~�۠dw�I�.Âo8��x�L˞���/c�4g�����,��e�fM|�ʹ�$�˳����ݽ���͆�ޗ�Z�!V!)gs�8BN�Q�~x�ϻBY��|a�E����9�-��6#B�I�<�Y�<�����zS.Ԋؒ�;�k0����T<4I�6��m�Lʹ*{���]E�g"�֦"h�">%>��|xJ �T�}d�C�\�̥��}��7�(�u�^f%mzl�=t�h�<2 D:����z,�W�>ή�����(��+��%ڭ�����#+��t)�.�gs
`znR�.���3�,h���~=ù��1�g#q	ڢ��"6�i�/-5<��7n����nsb�<����}l���	i���1��bϪ#�?�>�J���}(D�N�Ds"��q�o��np�A_:3�א/�4����Ǐ�ǘ��V��ݰ�)Ѻ��I��x�B�18Dr��^Y7����Si&��n &A2D�����E8ô�M�N�u&��J�zW�75!�������8AW!j�3D�t^+�_���p|$�=��y�-�Ī8~t�� mo�a�mE��M$�Pq�x�7���<W��Q%�"����	Ѝĵ6��X���{�Ȅ�'��㵤O��Ԫ:�T�b�0���)� �0�'jA ��?����%T`����g&��~�Q�S�!W�pV���ڟT!�ƛ~�"�IM�7�KF�)��H[���hf��ZD��~���ԽcƝS�Nh<52�!���gRc��H�	=�,	�ui�B��'J�����s��]�����S����m! ~���U����3�S`x�%N�߼���r>���9�T����@�+�Ǫ������ɘ#WO� �&8e�v7�e���gN�����w#��������C��C����g �\��J�Y��
<�����J��K���`[?f�w��X���-]4���42��t�E�a��7�WF�L�%��gD����u�����L������C�b^�����`؅`F��G�Po�6���W�)��v����jV�-/�a-�>����E��:Ѳ��\�i8�&�YQ�'5�B�\y�ɘ�fJ9�na!!�n��P�8��l�KNU�|k��#�蠵T���ൔ����]��*ek*g%�픇��:�p����`���E^�n�MF����&ܗ��Nvsa���0-��W�&�nu���~�l��\����p�gQ"�;��C�>��1����/�Ɣ����	��챲Qi��֥C��C���,e�I��Yy4��^ZmR��q�LM���*�c��넃�b���FR�p?��-c	���ȷcE�um�����0��XF^_ha���+�i��{'sI��ic5�����+2��:���Z�Lg�;� ��ai< �o�5O��˕>��WE����9S�x���cV&gk˜7�|�/��4���O�~L��y�Ty���kU�¿Z���QC���&��2J�!� �pGe�Ć�+�k�U��������p�q�Y_�hw8���a5V	|��I������)��k��G����U݋3å��Q��i���o '�תQ�YH�!��ϗ��q�	H*gc�<�B:M�#����%�p�����-�s򢻛O����T�
���W�i��|��3��E/<��ޖ���;	�7l��B���d=�-�d:+G����=��W�]�I#W	{Hg�G�����_�vj@zk�1��{�@#Y�[/[eCS!�t?�}6��=;Nl7�^H���V���L��Z�K��(��pn�N����������q����8������z�-Ӗ��zb�	��!���<�:����_��=x]
��%ĥ��%.�u�Zm�MY����*�_�^�:k�g:<��pV���n�̟��@�҉��XSD�	̡v�I˒��H�$ֿ�!�ٽp%���%�r����/�[6ӑqV"��Jt��b�;+F���[��Zd��,��YE�H5��q�^�	Ȝ��R�~*�%Ηo��Г@%�&���m$��k��K�|��l��� ��Er'~(K�8ŊY԰J�[����-e���-�u�TwO+�x{ �禷��k�\%��L�q@�q�&���z�=���ץ_uR_�a>"���Fx���=������0u�5��낛�8�A���$s�� �	��׬��s�u�n��w�B��)�0����EdT'1'fD^�.<"���t�P�
�a�Ĉ��^c�n��{�8)n��[��I����-]�"���©�7���P��i2��}���aJ�L��@�8����r�az�i�{�e�޳��2�/$=�Ƒ���m6��zE��ko�=h������?�4,�R$�f:�{�m����R(����P"�.e�����ڃ�&h2�|N���NTѶ�����z�V)蕡����s�����5������V"���^��%��S�$�_��n���s���S?�k]%6ቭ������Kx�	�lB�T���\�����EhW���^��Y_��@�l��ٳ�-p���\����%� O6+B�K�ic8�'��WD["�g882�4��a��1��D\q�����mx��������.��%�
���A4���;{.j?O\"ɩ��ƓJ��#��O��v�eݽ@It����"��[��z�)����y�L����a\2xx+�^��1��m����R�{�k]#bݾ�������lu�+����(4h�-������x=�B�m;�B-]!�F6	�m�(d�[�RY��4���3++�0�,���$���5�pI�1ɴC��~�����H����ٗ�7Q�qg� )&`��U�nԢ�m��R5m�)Xh�"E��,��ՔC
&�������x_(�G�i�)�E��[@�f� ���W��yޙ4����o������;��<���<�9����B٥�f[ʀ2u�L{���5��v�ז���v�<rC�4��V]QEU9W�#�0�p��|5��?�0Y�����B :Շ����y��ہi-W=՟�6���Q��� &X�|��PH����z���G�V�I��A7K�ٸX�`��5���\��ڵ���;������K��ԛP�=s�35n�~Ċ���t�j �pM�k��R`�]&�&�Ӛ�A��O��-S���dW?��5/'Z�"�����;��+�l ��ll��Ƨ/�y�2,�AYNA�i	~[\��*��Q�v��Q��<��-�X�� ���W���)3й�J��'��ojÁH�Ԯ�h�k%j�D���� oZ���gE�x��wrM�*�k��[{]^��փ�����L 
�|��H�0�%h��].ߍޱ�#�G���k/���%�<�K&�$� 6���O��yp�C�[:d`M�h�W,D��+�]:�+��������c	���1�V\`��Jo��@���fn��W�.�RA	κb'�4���t�=W�c�<0I>P�d#z�\�bh_:�``c.��Z��9L�f^EJ�[w��� Μ���q���`#��J��٭!����^��h,�M�2J��N�����owEL�v^r��dk�>-z��Ի��N�p��Հ�I�V]�r���p�����F�c�Q��B�������;R?�̢��C�x����3�(Y��so��ʖD��K�`����Kl�*�Z��+z���A�O�i٭��V�/�X�0!��$,�A������S�	�=��Ty<e�C=%�iUJaš���)u�+NN/�.Lֈ1Y����7K5���X�������s�~��~d2�0�̫Y���T+�n�'�0���bc�Ĩ.�;�*���y{��Q�{���zT�
z��M��#b�o�FYUJ��pb��?oU�zD_���m���U[u�������jNWH}�Ph�3C@G�}� �W0p� ��o@�� ��h��KZ`�UB;̎��L#�!JZ{q�M�.���pw�@z����@�(vT}�s����*���j3�X}M����	��B×t�5�K,Rh[+��7��~ݯ����DAm:�U��Ϳmywh����t�+�^�� �5툂ߋ�ߡeE;�;���V��j���D׉���Ri+)x��5sa" �3wg��� +"��J��*���m�L�ʺ�\*�6��S���bV���[�o�w[jhvg��p��d�k�V���N:��\�f��í�Dzg�w�g(ţ,��s꓌���\��պ��=�-z��2D:�*��;\�` G)qW�W*=w	�� �ȭ������uZ�/[�߃~����+������xj���\9����%� r=υۈ�~�=���rK=P�'�Ul!�(��
N)�'���V����uy;4�@S������3��RE�a�N���Mjs�����q���+����tlS6��_m�ھi;�^���i������!��o{�w�^�a������yo�[B!�}+��s�ؔG
���&�1��RO��8\����� 4��!������[�G-<��.��Y#��eeg Z��LQƋ(�׺
���s�3s�`��|�>�iaFFIt��9-�h��yEߖhå��/ZH�uм[ȹ�nw������i�;#�����'^��-���J���]����` �v}��[�:��ƹ�ё��.�9: -�s�ocxH������j���������ԘoI���j�y�vq�	/1�������'F���U+��0d��\�^����ΐ@�h!D�0c��2�P�9E�~�W�9U����Mt�s;�����5Ϥ��i�w�!/_j,sL8�S3sx�C-:I�,ˬ�+������(r���j߂V;��e�����x��xi ��A���VTДc�~�RF�R�q6�q%!5�aK�{�ׁ�/3#RV�O���-�m�EE�f�d
-�u�ǌ)(���AT�q���/�zK�0xS��a�'���]����ﵠ�CQ�O��0�0� ӦWF@����ɊU�h�io�j��R��kV�>��([h6�EC;�x�\6�|�|�I����1hU�g����+,���r��>�֡�!&�u�Q fÊxEouU!ݐ��tSHm�Q߭��)�{<u�]V�=x�X���ˁ��O�@�Jz��訒���M��!��=r�r1 t[g�K|�Hk�+�v	�'��:�I	��f������*'��|�f(ꏍ��s$|�1�S�P���#5#�Eɣ��&^½�a�b�s5�!� 6ͤ
��9W���2�.���f��?�D-G�u����Yf�n2`���v#��D�:� 5
)�%'� ��rg@�)����#:)�ڟ��1^��DP��6ru�"qM�, q���������!������Z�?פYA�"�p��{�IJ���+���R˳6�}y|����/�C�����T�#�7U}~|��c���aK��I�Ʋ�be���3����+ٳ����α�e���m4Q�P�����z�FS(��{��>R�^:�@|b�^��ܤZ�_M�*>����5�(�.��u��gbz�.�$��Q��[,����}�'"ȳd^#I�M����c�>qM��r!�ϡ6���)`R�b�-�(���(�����%�>��5�QX�i#*���k�&�°�S-;+�ƒ�)������Y�s�b�G���<�'�Ӝ}���J��)�Mc��z~�J+����I�h=`��q������f�[�Vї1"B�[{��0��q�;B\�N��wJ���j�u��ү�Ц�;�Q�!�@�k5��?�$��&t/4�G����o�B��Ki�x:3�9H7U�KX���nPv��8K�-N��s�AO���U�GZ����/LT2��zAFs�i����T��q)��ٮ�ƒ��[<����s��-�!$(���B����D�"�d���A��2m�����J<=�i.Z>�^���h�u�>�Vu=~�Ԉ C5�d&:N�S��F��w�����W�J�m��䫧����h}r�>��{�cX�.X�nf��%�4%����H����r��k�U�ƙ��e�SǴ��jO��{��5ﵯ5�v&��ڕ)���Zx��k�F�w?&4� a���������=�=}��i0�~	��P�j��>{O�-�?4�f�G��B{��y�C�M�f�=c���a��հ�1��K�ո�~�����~bA������П�[)H~��<�񒷀Hʣ����f�'<�{+E}�ޯ��/����#�YZ�������J6����&����:�����q�Q��A||�9\�9ǉ�n��(7{�(�ܛuC5��#������PLIS29Lakn��=�QY�؍A��(O?�����xVfň"�R�z{I�H������t'��8ΡJn�+F&��^��,�"�R!�gc.��Ї�PQ�.�@k@���+ni�XGӵ��k<S�>���Fu���kZ�˧�$'c��z`g/T��b⸿R��	��ǉ�[58���r��Y��Y�@��.�61��qP,��{6|�5�bu˛t����v ˿��3�-k0���a?��\�
�L�<#Y��0��S	z��椧4����7���A�������������yv���DWƜG�ʮ�oJZ����T[�*t��K Z���8��,/ai[L��$���	&��g	��$�d�#�ϱ��F� H߶A�C)CfE��f|"�*��4����n#�� ���?��(|u{�&55��P/�N����)�Ϛ�oD��:0Ȭ�M��x�$b��1nR��1��b�x�gW�������Uf�sӞ)@���d��HL��p
G�,o�L��p���=�c��]�h疜����}�������9���3(�N\�H�itS �,�Ty� ��ʂX�g��
�|������Hy�U�M^5���PP~����%b�{�G��L ���m1��4�-0�%��0#M|�Vb����u
�~��bb�;���j`�Z<" ��'�Q�"�r�r�{Tl�g������YV�d=���N��E�@��:vG!�ر3NW��bѓ��V�M�j'�<.+z*{"���u�e�	��3	-)مl}��䒘�.?�M�{��y0��wq����O~J�҂9��L�Ps Ŕ-2��4�d�#$��-��p����+=��٦��1st��Y��Z9-Y�%�q�����4�_��Y\n9GZX�����*�:�Q�)������Έ^s?X+��C����x񳤼�����a��XR��
�����I��|��޶��Rdy���Z���v ���,we'��>���D� '��B�I�=/i�����;�A�X�Œ k^��  zb�Od��I�ꢨj�K�բN�� nGW�w��ߔR*����k��$z!FW��w�"�����<u�z�zB0��1�W���G�JMb��w��������N�,�k��j$�ߙR����[�Ө�� �|�d[�	���I����lH���"��C��k������}�|�i,Mi5y6@߰��ԃU�QY�'��l+�� �B��>�%>^���9��3�W�I��rË��m��4���i>W�f ��z����b��y8k������z����6=�dWj�b�A�!��AT�����9I�/;��Q�IRFN�ݍm�r�c�U�@�3���Wz�	��<�� �O��3� gզX����?��3�����=MQ1�>���ho�[�r҅G�����^x��S�L>	ݻ�Ӗΐ~<���c����O8h��˃��xv@׏mv��(�t����B_�#�귅U��[4��}*|�o����*�G`O�rѢ��
������P��m�[x{�H����VV���d5�A���/�}��K0�����0~�TG(z`��^����|��]��@����G�UG��ly���dKL�7[��ᬁ�LLu���3K��C�
�E�l�I���a)����jS4���Vd&C�j}j��vz6���^�.B�y��(���o�w�t�I|���ܙ�]��
;�B���7���������s5a+<n>ɇ�����8ZI��ʑ]�L@�bWH~Ц>uA��{�9�O�]��sb�0r�f�_
�nf�0���#�׎�*�5��M�Qi�%�v�����}�ʣ��c��������4���1�����];3N�<��>M���~���\G}��8�0v5y-�au�{hO�v@o��q�U�E��&�p&˹v����w��x5=(�Vb��E�.��,��f�_|��%�JQ ������A�b��	=�cN�� K�5R��4�$^�z}��������|���V�ń�4���!���<:7 �\#s�*�{�Z	�໷h��T���t��O�ަ"=u�:��i�4�FDomǑJN�w	0�g���u4�m☖�RS
�R5��H	��=){K��-j(�f���n�B iz�n��
�A�O)��l���⪫l���d�D���n����8�G����ћ� �������>A|�|��Q����e�^��6��w.V-��������.�,�Lg����~��ű�SU�v�Ѐ( ����Do(��G.�zL��6#�?�$���8_*�x�>?_h���`�0���ܣ�ܑadS/f�2�2���?;J�0�#3̰!�%��Y�7(k��X�7�`�j�InB8F�՗*#
;s����y���#��FII�~�����Y�@W�*`����攃�W,KK�b��p$�O��
�|Q!J�`4!F����Gb�����`l�^�����J,-	k�5�'����ċt�u��b }� \��<�Y��4u�ǩ�'�36�0�i��d�����\���m���)�u��W!���n^O���K��W��f�v�����N6HTwT���+���w�h5,��t�݄1�e��;�ξ�؛�/f�gUrV��W����v����@���e��G����X��������v���1�3J�\A��:�+���jREi�D���ʛ���%Ca �Lԣ
?�� 8Z5����&.��/ѰU}a���)Ka̩�/�l<EZ�W��}l�tZ(��f8T8ȩ��T��]����z>�X>+_�򨞯��^"��Br)�9�e�l��셪�����جAż��*y���c��ٱ��d��:���q&	��r�����<@~�~BI"q�Y�S0�߇Oq�x�+�>�ae_�D*��4�7������r�����ּH6�)���ՄD0#q�Au�ɽ�G�^يN��-�������\e畤E�KNk*=�@S̀���NrָP�����5��q��G�X�<l�O���2!�6���p��)�gI�x��.U9��d�`�����*7{�t�ܖ>M��m��OSo���b��[�o��i�s3�ߚeG�1+���s�7�3=9�{��Gݢ�ʝ.�=z}�g��1h~��j�s��j���~ݯ©���y�]����ɏ�c����Lt⟥���#\�{Q~�@�şB�MT^i������;�>B�zW5nZ�E�% �W�x����dQ��-���p��lZ���p�-@��7nM����R�y#�`�m'(a��� (z_��c��n1�@����s?�+)g�e#�/�c#���J�^=�c7��UB�<�Q�[�c/��q�����yĸ��GgЃ9�"�/O�Qo�DB%��W��z䒿L+�R�Xh}7�H��z H�n&H(q?r_�[p_��6���
�/�_��G�5R;���8'�EEms(--�&q�������Z�T-�:y�����>.%������]��M��������(Ġ�;;-���p�7%͝%���m��[�ٱ�q�h�q���3�l����a�P�x���:mô�&W��V�{e���,g&�u,=��ֆ������3>�ǵ��f��q��4#{A��+O�a.��=�-�}<�{F��}�������"�A\��T'�q^G�u�w�Uzv��A�%�X�t��i�����h��y�3ĭJ;�'q^�F�C����8����$٠Ը��_�!��l�%�s_�z�藐a�bHez6�v��#ya��3n,�ӏB[�&��a%����xd�o�M�Ut�w�+�%M�����{]���dc��~�J��Ag6�ȩ����xq��qD��3~R��IGHQ�{*�k���Ȣϋ2�-�<�R-n�,��=r*窸VEy����6Yy��	w��Z�S^�W��ܢ_�������+�w�&/]Y>���ab��-���KUm�m9�dv5��V��C��ַ�+O��lӯ�Е]��W^���P*�X V�x�l������>?q�a���(�pP&��}І4J��%���o4����`���Љ��L�u.�0X��� ��N��l٪�'=��:[aO_+fhZ��na�<�[�_Gn���U���������2�i�Q8%¿����tŴB�s�CS�;��|mNK^]�O��F��m_�ڴ��Ӂ�W9���=�F�U�߫����u�ӯ�f!����/��:�*H�J��~�t�חO�z��[�ͤJME���IQڦ(=��-Ne�~�	r��ׁH����d4��ۙ+�|���6�J�3m�+� �`�M^A�P�[r�+���M��İf�CQf`qRU|Ju�i�;ЛY��d#6�f�pv/�V�Ӻà^;�p̟~���}��FYr �Aj�w�Nw���֝}���T�R��"��g�]��̸����L꺷ϟ�to�|�aA��_g܌�R� �\j�%-ķ4�iA�D(f`e��٣N��Q_\G�$I�#]�Z��^8];8`1`�� f�j��
���!��ρ�]@.��"S�⇗�o�d�I���4B5.�����Rg���Tvl-/J)�y�����݂�B�zX���������~��%ZI�ϵ�u���$�]�V��߂גK��?&�%�E�f�����vѻ�2��C�����|��!�Ũ�ȷ�#������	���j�:��=^cey I�t���8j��Cj�����$�-�<j'�i�P<_[0� ��z��)�=�S�n�Ǝ��~O�a����z}Hp�)gK��s�������+Va��HDx�<[N)D #=��m�S����O�M����dw2�=�G��<m����-�IoF�Ǟ����5�9<��W�Ο'��s��$^���MSx1^C]�2o��CJ�~h�z
�Un��{`Y	�|���,yA���9�>���K?߯++��>�+��k�%�?}��X<��)�9,���|�|ZP&>��)�|�}U3A�M�4R0�M aخK���1:�O���1�B�6�����&!o`f������9���5�S�2.��нF��	����^QYҾ�o�j�qIfumS/��*+���E��ڈ��Z��)[��v�W�㤒�� ���[ИC�T<Ӥ�� *Ε۳3����΄J�����zV&�7��q��p+�n�S~U�ZI�0�`�x������8B-��!H������.0���u��o�_����V��n�9�+�U�^���杢�M�"�5?!c�4n�T�աg�������0.� ���}X�y�I�q:�e:|��g�Tϟ ��#U(H ���v��Jw�yv$tNw O��cy��R��>6�;���pGHwr�cb#��g�r�����ͷ��7��wx�#.��b\!�ԫ�|3Q؁[�Gt �n�����V�_�����whk9xע�l���p��#��Ļ�I�G��@��;��'���wY���x'U��Z�B3N|@[g$��v�z��Lv��^���ʀ}�Gt���ϝۀŰt�,a6Z+J����)_�u�6k�s�����mϗ�J�i��,�p(�'Q6���@7
��RwT�f���6�T�x`��9��J� Hء�����eC���⚻q�!�.ތ�7zxI2�o ��$�J�JZ�y���o��o��r>�Q�2�D��1Q`Rǽ��$G�G��L���C�;E�7�b���L�\K� ��v>$�JU�)<��q  �(i���U-�
�n�1�W��P����@AGvU�_5F��j��xJ�C&}3���Um~O��?���4+�9���H�߱{3)������4سHI��>	�ى0��tΰ�
�aI�YZ�mٌ�!��4�� N�����^��5� G�[&��G���p��I���OK��)A����
Z�*���Y�4�.��aQ�ݯwM0q�O����N �}�^.�6(G�Lj�������s?jB�sT#����7�p��<�GS�c����6��\�}���tG	�#+DH�����o�j�m����V� �K�m:PB�98�Jn��r�[� <'��?j�s��eK3a��Js��1D���J��E�8ѫͼSPn��r�m̵i���63� kN��td�挈�q�^��_h����L���p�gG�r���#ȕ���PJO�W��6O�h�YhO��y�I�J�f�z���;p��Y�D�{�<M�����R�Q��]��
��9��V|�a_^�9�jW��H�ն���(�~�9'Ly�p֛�[%j��YK�-�ac�s�ڎP�����A��3��J2�4�	�E�8f���P��F�2�^q���c`||R[�����*p�kq;������ǉGČ�z�*��Ur�HOm{��t_+uH9�}×�o���)]/��n��O5��➗��AX�	���p8����/#$��B�����K��_-��(uF�`^�eцKU?y[ip�*c��CE�o��
�n�����B=�Bpa�ooiS(�5I���ͅi�^3�Bb��/�����qa�@~',��
&�W�?H*!Y|�e�{��݄T0O�8(O�w�;��< �4*��*Z~�9�V!��@Fx��9�_��-�X9p�q�ذ`�)�&G	�)u�V�n�[��9���,��%n{�c�2���/�g�8A�`�3��ޠ.�p���H+\�A���gM�k�)�;J��D�
�H9sy���P�>#�"�uz��cڹ2�U�&�N�	�R��U���T*�vc�!,4��2�Z�x���
�˼��i�6R\X��1�3��p9zȪ���C��[�p?L}s-�N38n���i��P��p6�P|�+�������HkS�l�#����|�F��ua��u�_��w�{��U��������B�1�ڦ6�"��;>��;�uҚ�f�&��r-̕������~)�Pj��*�U"8=e���b��<u:�;̤�,����Ti��׷5C(�DS��r�NA]�6�`��q��C�68�Pt��	���^��������'�a}�:C��D�prt`#��8F9�Z@����������Nr�-��������!�<'f4�TRm���7�ڨ�%���ryw4,�u��N\�	@uW���]�aw�?G��*�^;�+vVz8��׶����ʣ�P������xE_#�7S~��vv������7�_�QP���[/��h����ޟ�.��0�S��	�=��u1S���;�=��k|�v7J�x
ޟ7�6���k����[9�I���/hle��l���?��Ӄn�b�e77s��C��kn[�+�㨱���娒��z]l�i=�Fx˷�d�+R|���2J5Qc5 �I	��(\����~�)u��q!�.��O��DO�J���d��D�~�I浦<����7�I$�e���=2�v�,�������:�	�Li�*�������Jڔ�P�~q��.����ca[r�|�����JDmҳ�����_��j��V�pu�nU3�uQaF��?�q/�}�TcX�q/eL�`�*u�Z�@q���N�:���5���~�]ݥ�6�e���4���M�+"s^�`��r�o(Ϻ3�A#K�uC)R�D�z�k���}���&~���� !7k�g��rᑯç"�o�x_���oa�H���v�i
�l���8~�������/��'����:����N�xCSc�E���X]ކ
𱗉k(�`�?����2	OeX��N�o|���y�a$R�X�,׷[&����8��$�iqA�S��ݯ'��1��βL���W�sNrr��f�LK��hl�71�o!���I����el�I��b+�%��<��%���f)ʦҏ&�0U0RCZ�����|���r�9�8��,ˎm9	r0�ai����z�������X<���J5B�:��Z��%4�H'uV:��[?�{����:Lw�i �:/j��#��ӝ��[���=�7c$��ꦮPV�*�f��&Õi3��7i���Tݘ��[��E��K��n�c_�E���&97�*��H��v.����Ƚ��r�!��!��E�Iҝz�
�X�R_B͌9�#uY�z�Nn���hP}ǉ�hX����t���r�[���]����P\�Q����!�Z�S����W>	����|���~�K��l�tyYd@`�X���-�Й�ӛ)Ӧ�-��>�k�����e��N���� IN����;sx�# ~>M1A2�ٲ��w� %�1p���C�����>��cF��Q�sL��4�玠+;CYl��I0����C��IX�C��	�>�^�$,߉��q�}3k�<LpZ��o�ȯ���.�LU�0��x3�qJ�xV��٤ΐ�8w��Q����\�G��@:U�!��ۓA��Gvu��D#�,�����,p���bdu�l!�������$f'KF �����y� H�^v��㥒�(+�����^���#)؋5O�z��O(�&�[ ���η��ԣw��$���H�-0i�I�J`��<�~�粻������t)��y�?�3>�rJ�E�2�P����R�e����m^�����d�:֍���Jɔ�pa��]Ř�U��hf��F!~�\�ұ��1cs��.3�|P��	�q�%[Z����7(e��|�~I�Y�sL� pC�pq�I������k:BR�m<(�Vü\�PK��E2V- z�u�[ﱵ���!p?,��ي�ʙ�״K�CE�ߠii�=z}�	���s��2my��TAOb�+Q����ꥈ���t$ρ�#w�֠�?sN��z����LR��v([{�;̈́Ơ"�U]a� �7�K�s6%a3��^gAv�äs��1�Q<B���I,;	c���D��(�$�%�tPN��/��0]�̞.����M���$���4Wyhw�������г��Ӎ�����f�	�P���y��{o&fb[��@�����t��C;���^����K���Pj��g(���̞ѡ=��m%��v�w����
�U����Ϡ+����p42�����o,���?ts��T��"O3�T/�E�����	�[rF��w��-�&w�#N�E�4ؗ�%b6�qw����f)�DS�M�G`i�R`a���+�g��R$�_���T
 �E�I�0��!A�Z�SL�DoC':�)�JNk\��o�89L���������o�7:������4+�m�M]$�3[Y�E-�z ���o��&-�f*;�;Y[�Ζ?ɹ���/���+�|D�7A^�@���P�R7�C�.�-IF_��� q�M�&��.�ϥ��WYܯ��Ex�t/���Ms�p�N��y�< .�]�Q(��n G�|@��� t���3Y]л�-e�V~��n�\�ֲbh��/�#��zr�
򗲅� 6��Y>�V/�-��t���r�e�c��@�Yu�y�lZR�i�2;I�㾐���í,��l��tj�x~x���ic��H���:BZrE�� ���ژN���d�*&�����ڸ�&�o�����i�%�������\�JPl�*�D<�<ز�|Mj�� /G~�v�'�M���Â�6	n��80)?�Յ���=S˟wX����G��g�������+�%~���O�[���=����	W����SV�*��z�c$�>�b� =��eN��4Jj)>1��9>Uk�-�?M�=R��h�Pkݷ	7���ؘ�/`�O^�=��>$�w�%�q7`W����Ԋ~�za��6Cq�GX!�(�3E�o4r����G�pW3s�DL��ԹJ�I�	_�FS�6�nE�@�;�*~�N�9���=�S\�F��W��p-^2n��Ђ�I@p�ȶ�vmՔ:���>��|?�!!�D�sH���x����ݴ��	����W�}f��6~�-pk�eR<���+ � }e[xs����M%i�vC?Dʟ������^jQp�z�4����Ci+3��|�����
������M�'���m|=�"�J�5����X��?��d]�
����QM�ԇd��;���ASJ��7�ܲ[�lա���j�'����n\U�B���;� �]}���>�S�����ߔi쫩�6��~N�*��0�a�b���5)���ս��ntK�쌅U�G,��kv�w�t���ʄ �Ӗ��
�訒v&,G~�L�mJ�ZА�o.L����C��lы����8���k9v^�<�َ;�m򌕧ǈ����3��q�pX�gSc��7h�lh���ciR|�:��J���J�۰Ǚ�2c��(FRL<�S����2�8f��є�o�ifC�Wg`W�G^��m��lr�J��rVb�L���=��#e�ū_���L�L_���aH�Z#�b��&%[���cE_#=j��0q������ߋS���8�L��@O7�E�`�7��X�YӍ�F��ݯ���K�<&�tN ��)��qp�
����?����u~#*���rVV���S�����ht���l����"Ǡ�igl���$	�j�O�>�AuX<( �]������%H�$�o���p+��?�!?W>�y
��I.	�Z<7��J����d+Ǎ��/U��rc�>eop�C0Dv�d��X�����4/��~΁��j����~7�G�� ���V#��0T&��\�w�Z=��ʩЏ����&���6Cg�J���sᑨ��1�cV! ���\�ueˆ<е|�+�dW^^����:e�tUG�Μ��םE�|��Uj�Y�j�\k$��5���|%4��ɥƷG�����	k|�{[v�qU�p�Zv��_h{{��ߑ	/���T�f#�rGk�\�<�(/��d��=uz�Z��f��墕2���z=���w; O��Z8�� �/L�΁�� O�� Q�ve�H��pQ��d���"�b���;�0TM�y
��4��o69aK� >rYJR(��.;�.�!y�2�{1�y�A� y���O;|&�����e����<x�:%���r���:@;�KRb�[%E�~�[K`1�� t���^C�DkW6�x�g�_1�,ό��I���<��R�N��*�߽��=rb�ɱ�#'�Y�.Nx@*5���%�����T������bU����|3��b(й^��[�iۏ����4V���?Ƒ;k Rw��苧���s1�Z���.#D���yq�0Lb�1\G��B��Q���AW�2��#
�b��R�5�itT5�۝�	X�+��b�-�?�<䷘+�w�3L��E_�j;U���!Fx��?TR�e��q���/h���]�I�׮�!Mv�2�Չ�,��Rv�0�e+�3�Z-����cS���Zg��)ù�1>!^�����"�ڮ<�=��d��ڛ���#*�lUVb�+���ޑp7&;�.�XbI;���k��sQ��ظK�5� �c�G��T���	���q=������2��J��'x��T���6;��_�?�(�ogkx -P��]����j��%#x�m�,ƢD�DWJ�N�Y��$�4����q�Tv0��~N��WH+�m�}�ǹ���٠UǾ`3!���sTT-A.]Q�q<�����,��y�Sov���.i�/G�b�BE����&՞`!Y��gP#����$^igjD�鉖�Yk�^⺕�����i2�\�C�A`mԞ��s@@=&�8+Vf[I)0� l�����pz�L�s-�s��%�$�
���-Ϸ�����Gɖ�,�0�l�1�l�ea�V��c�+#�`�6t��<*�c�kmY�n�s��cH^b�#�򻆖��9?f�n�e��n
ˡ���x�z�l�"��6�ٶ0�����]�YX#۶�Q�?x�����4^8�[]�,"Vv�pɧ�< ύ����g	�K�����24�4�ϴ.�2��3ba�f�)��̘MK�eG�����NҌ��QQ09
�C����1�6��мJU&zI��oZ8�e��}��?��nNO�^7'�Zl#w݋䅩y[�j��3�;*��o���0����Γ�e��8`�n?t6�eK���V�3��<<�k��=�/���;=�-6LL�'�o���G��+0���Y�Y���
,�=VV`�'�ۈ��KZ[�~�|�-��珒)���5�H@#;�\�ڼ�[�3�x��y�#J
)���{���~Kpi%tǆ����)�3�d%u��W��1�7���A�Z4
�3;��(�y-	[ﻖ��e�p�3|{ZrmZ?�4oy����oal� �f�(2�$�\����"�i�q��DP��>���X�_r����h�����W��#�(�}�Tn˶j��+[��Pbg��]��3�k]��+�B�Ax�HU��a���[���G��j��o�������\6��Kn�8A���� �9Y&ٕȲ̲+�e�JfYVٕʲl�c��h���L�^�����(z�p����-�478�T��||����uѹ���8��E� 8,[4\����>�>��~3YzA���@��T�˽���Ԕ}���X�r#��F�	��~2"�t@�	`�e*B�� @~�X��?ƗB�X�@�X�#W�5E�r�F 2	^ڨ�	��x���
��$_�n��(�������fK�^r��}1̔����0��+��JTsa��P��,։޿�$��M��B[$�l�m���+� �;����8/n�S��|�`���-���V�q��[يj�{���:F����i��n�2c�5OǊE���;��eZ��ҒYZj3�x�=�G�cyRj
���4�8��,Ѥ�5K\�)�M��ya2x�g��!P���T�Q36D�5���F6$Ƥ�ؓD�+<�!���ß�v�<w��hL����v4WK�*�a���;�N`� bVV�9�n�����O���<�Z8F�]���c�ؗcw�H6�E\l.��Z����~S�c��[��,R⏋���	|�c��4��U�}1-����纹p�̖S��B��l:%���S��{�[n����t��
y�򝸿�jU�V�߳0ܮ�L!$|�ԝ&�6��W,7ߓݴw�iu5^q��<pJ�.l�3A|b���t�ۆ��e�3���3���=����\��s�ڿ���+%��<j�v|����/n�W�7����o%*�L�F6nX10�~>L ��Ѵp(��H�Ǘ�;t��$L�O�JN"z��n	��*ܥ>,���Y�̽����s+^�sS�9~��K�o��Z��	��,��Ж���7~�G%�9�Z�RW��F�TŽ�D�]7��*��v'�G�o�I?�k��5(g��J;ͬa������f�$$�X|��6p2�C�3�Y�/��. ��gX�qW�Aګ!�;B���`��n�
"Ы6R؉>̋��;�����xn��\�>b��q�U; ��M��L3�0x�)qsy/��K�(�2�%��f�E��g>�)��m��m�M�ݻd���!ݾ)�6�����%�N�繤dS�8���'�-��{�@�2��ly��녔�?��t� )|'Y��ڴ�@���d��e#خ%@�%����i��1�̖���MǻOm!�������jA��W��8}����8�kI�u�C1��O�p�X�	t�ը�D���Ɂ�Pb�p9�F,e ��1pbr
+q�~��C�S�I@H��C��o�!5(���08� �~�ZH�������s���9���(�g�A2��\��l�P�,�L��ب���~'�<�����^~S�aTK����Ū|�Lj�z`_�G���.�����V� q%3h,կp_�>�����j��
T+�Ү���T|b/t�.�->j�k�6	kr7f�{��W����,�*�\Z���U�rd�@��܆V��ػ�������b�+�֑�$�rR ��TKC�:���(w 
��w�3�S�%����s7dc%���89k����v���Y���-g���<�s����&��M�ل*�+ctV�0�޳�규��mѵ��O����%<.�2e�7�������+�~0���C_������q�
ȍ�I�Hq��V��Ei��<DQ�N@��N��A9�3�2�Wr���pI�iuT����i�߂���E&;�� �����]fy�t���k�Ay�g!5����aU��gOӎ����X�@M+=���R�p� �F�~�9���* q��������ԧ:�pzz�×��\���%(��Qx8�����$Ry*W�����}�rM�'Y�nɒr0��;X�*O�eV�`P~&�e��L��2c٣��=�?��Gj@�A� ��-�I��_��������[���G�R��>�7F���&���ͷj�O�o��u9Kh�_���Z�$�-�8H�X��r#������N����(�s-����+^3�<���Iv�e8��s-�cf��`t��=j��%ʅJl��dڟ"�
��5B��*b����=CMb�$�0��E3מ�tB���iRiQV�L
#���Z�?;
n����F���8�(��6n&��3)�s�I1ɏ�p�Wh��)S��@�	�2�8?j��r"	1u)�K��u�<������!��LOs��Q�y��rW���^�B��Xr����i�4�B�Un]HԜ��M���SQ}}WH˪d�5�ڥ7����Twe_������������K��.]O�í��ʿ��ό�����u�ja�e�?��W��9E���͗�Y�M���]�+�5��-�i����&�M�Z�ev�u��n�2��g"*�O�6�
)݊ʖ|v%�Q�X����D�؝�%I���A7?�H�!|����U�?��$�'�)���m�^( �CH��a�c�Q�q�-vsQ��w�Kش�u��H�E�fF��߶5�<����Ζ��
�~�d�IvӜ�����-����Fd#jy�)��,���a��|���0�A��5�k̍�ˑ@sl-�E�ܽ��M����ґ@S��˾��ښDx[�վz���+@rIvT5T�cg�[����n�a�"�Jt45�B&�lk,[bôM8z��ƪ���tKc����7H���ڱ��:x��Q��`K�A5ʖ7x��A�3�|��y�#�<�Zx�:	�p�O�k8ڍo��o�{��|>��ܙ�rz�'��x �фQ��X#�`
�\N�K��J��#�kvɏԡ+�IR��~"Pm�h���'�X@��c���<���6�\�<��r���r-�$+˵�1h���ȓbYn�<)���ɓ�,�.O�g�����p�*����Pni�X�]�)׻�9�Gi�[��f�-S
����\&��s�n�I��(��X���O���v���-Q���~���f��uF`��H��T"�m�Q𞔃��M��pҷ��w�c��3E��Q���F���}���f�t�?fH�ޒ����D3�O�D�?��� =��RՕ{�BeR(����?���;�Q�'�2pR|����0\1͌��i�m�f�3l,�&gİ�9#��Ţ��'g�Y�]Έa[�H`i	�t`(�txo��"���*Y�QL�U��'�>���;��4c%�K��A��5Z��Z�:�� U#��¹�8��b8|�&l�����D���6Ѐ���Y���><�/��1ȏ��jw&��%�����\�q>��ІD�͆�c=�0�� ��G�&���/V�D�l��S��;!�)
Y\���.�^�M�e�1�� H�WƝ'�j?2:��[�L�>5��&8a(y�O���8K�q��b],��`�^H	��sT���Sc"wn3\E�?�$Fhk6�}��ߣ���Պ޴�ud�(UiDIvDL�x��eӳ�9t2�Pb��j��Vb���P9+�;��i%�^֊_M��@��4�<�[��E#:��0����})J��8�g����S�[�'�B���>��m�t�.[K����Q�S9����3���7�n��(�*X����T3W\�3�7�$�bk.��у�+˕M�e �N���X��nц�� ����td�#�}V:���M�z���:���X:�ü&td�#;��Q<9d�#�v�ZBgL�z��M�Tj��gr�K��.9�]r����RN�K��.击T��})�(�5}@RkK�n�q�s��i|P��������h"�M��v��Y�G{*Q{*�=U�G���S�ٙ �kX@�M	?�����Z�h�zq��΁Te<��� ��{�k��.���f�}���H�����[H�d����-	 �"}/��F��
h��©���3����~���Q�mt�x��Έk���yGTx[Jݑݞ\�ȫM������Of����e<a�m���)&���x������\�O��	C���F�Ph�&����PC\:���jb{Xq��"�ӹ.�k5�:�u�5rcX��\MQ���א��Q3�mR�U~��H@/�%�� /����A|U��<F�������s4�çn%��w�̽S�����I#u�~?������߸�@���������'�W��
�XZ�D��P+��N�5��i^��X���/��Ѩ�M����U2Z�F�V����D����<.��L�ҥ�wF���99��2c�1�+ۄ	�ȬզBK�j��m�#�ɶ�y�d��y�d��y�dc-�*:����ʎ�#�+&2A�Ũ�)% $���A��T���:�"}��:�R:��$�D�(g'�_:�j��K���"O��Ĕ�4T~mH��x�LDT')*mF�{����,@�u�b�ABR�54l�R;Q1:B ��^��=���G^jC]�.���Xٵ6�`� y:VF�Uq��ak�N!�Խ���2�5���:?��O�n_���1�[�#�/�I���ϸVZ*x�"��)#��6�f���I^�`�m!�V����yf �=貟d��꣥���sZ�HG0T93R�"��Hg�_�ڢ
L��h>��)�D�!�U���\�n�I���|� ܉C�4�y�I�o5�#<5f( ���r��,��k �~����"0���TD�zGSQ_�xxE�����`F���P^%E�4|�Яѡ�Ӣ"pt���<�z����y���Ո���k^��/���(�5<����\5�/0#�&��z7r�ޖ�PTozߡ���|��ZLC}���ܯ�u����;�,U���mb)n9+B߹���Q�-�jԷV���
m]�����qù��i�.��w��c����D�y�o�R�"t-��}z{���JA>�(q/�z�=��r; �1���m����3���J� X�QP�R�R�bhՠ
���\��h�*��ҽ�/m�K��$6��|~IQn>IsYr��,��Ks�a=F�(>�h��Q��g�1�3\���n�tq���2V;�Kj~L0s_w�Ƈ��{��>i?q�(��'�U��e�_��=�v�B�}s�Y�h������[���5��ռ4���@�A}��Rc�tYWH;�Ƃ��p@�޻q��)1(����sqW�bAN�5���Mʄ��C����֖(&8I!��_r�	1�!��*(�?E�ƹ�#��Sr�	]+ ��`J�����$���u���Tw_��<=�:��0����ڥ,� �Tj��&��6�H/�.�>5p��kp���c�,�g�o���o��s��n,����F������S�2Q�5j�ƪ�=M'�Ͽ��QU\����_�E�7�jitJ��K�ZcJ���v���cEd�GO�BkoZQx{꼐V_���.���[`{mK�a[8�24��e�g�7����Y�@����p��+��+�t���|u��>| �3B��Qe�Ѯ�O�!�q�����g�2pyG��I��"yƓ]C����|'u�&zGqu�jN���lڰ)Y�C�ە7�8�p�aM`V��6M����ZxFڏY,D�i>3�xʠWv�$S"��:~�2��08�xIp�9�FW��8J1��J{�[��oa����;��#F��4tgc�����e��+�ew�iK8��oA���p9���k�}���̏��T��~�=�ڒH��C�j�վV����D�8΢�7d~x}��U��ݟ����e�f�3n��b_��??��~�a�G���9oDyh��C0��~��Z%��`�PuO�ٕ��;�C�T0Gg6��C��|��[�N�@K�	~��Y�oQu��h���}n�l�P�߀���3[�.��8Ϟ���6ioRnD���N֊�Q�e�Nu��A���YrF��+��vP�\/��a��t?��@>�t�c�Ze�����Q�����*������2�	"q��;Ҙ���aD�y@���)�ZӮDo"�9�T!�X�ڮ�Ƌ�ٚ����
T%��` X퉘{�1�8n/|�����KHi.��u�VA��$=�l�8�2���T��&��̧���F��o-S�Zԣ�S�������C�$>�О�;�yz��U	m���+��N�����E�T�~����_;��I`��1؎ڕZg����q�)I���)���h�V��BJ�)`�� �� �+�W��X<i&�M;�f�<������˽F���w��'����I�>:���n��a�9������R?��]T�g_���Q�I�M�l���Oc���y;QvbuI9?�"?�x�n�V�v@Xh~>��XK�f/�6���S�R�N����x&�@�h-��U��z��;#��n��Ó��\5�۹Tz&֮������V��\���v&�x�ZW��?��,���?;|����Q��W-����Y7��+u���tP��Sh�?��������D�D}���G�ϣ~µR�B�]�Q�n��/��[��3��aI��R��{ \�VK�ĵU���z�	��|'�\����w��u��(��b�$_�[i(Me�78�9�$!�*����ڻ�7U��I� �S1J�
"l�Jk+�6�Q
[�E��T&�V(PL2zv2��ml��sn��^h���(��"Rn�M�|��w���{���y�'�򻾿�~�3(��FG�=��_r���K�7UW���Nʖ��_�{���Q�����o��N����Z�.6�l)0��\�M"+�L���9%��&������)�����	�%��9Д'ss��Ú~ʵ���0rZ."Q��g)��\�k�	?��>���$��vZ�c�6H�͘mpO2J��+���R#�h����5�bۺ��-^�$d4:���Vu�$�"sL���י(=��ؐhS�����i;b���ꮈ����ɇ��=���̋��v�����@@TJ6���eG�9�A�0�Zc 5C���[�x�з�a�����ǀ4��-���
��<��'�Z�j�i���P�W�Sh� ����X��m�����ن����k�� Ih��J�K��P���c(]H�� 4���` Mu����I�;�(9� �ԔL!Va�ʟ�FV 񔎿1���f�Sr$�T��F��WVٲ�C�|l�+"�|vDC	u�Z����W���j��[!~�i(�G��>�����t��8R�)���$,F��DHpL��<Q�l�ٺl�Z_��;�n�:�䧵;�=������]ᛛz�H8M�S+��ʤ���O�f�n�5�Y����i�5��Oz����h.֌�Gkz��|рg�~g|j�GB;c��o!S=��*�� E�桽������U��S� ��7��Ԫ.~ ,�b�~:/"�����`�'ݩw��Wҝ*���~���(�
��`Rd�z�&��ڸ�͘�����𣨿��iB��T,'��Ma΃��c6@A�0sk��)�
�ɭ�7���j`�#H�]��:�|�Bd��#m�no�cW��E��,�����)Q���kɲ��[nK_f%uO�|����^��������%?f�C�� nV�E_|5
��M�בc��s��O��kc���$s��v����w�ih�\ &P�\��c�h<��B\�h%Q�F�&�t�(�G�����R�0�8�4��J¬i�:;�}˝��ʡ����&YE��̅��i�� .	���akۓ0����+�f�+�����o�y��`�Iޡ��H�1���+p�I7z��$��Qݽ"w�+d�3]L�R��o�5vc~6RddpB?�?@򥪌Ǎ�;�ocF`�٫��a}�S��g�@�I�������U���H�m�X��l��x�ْ�At������ԧ�1/�x��WW�A�ރɫ�5���o@�ߦ�띏�g�l�3�X6����Wxc-iE�2Ñ�|=1�á_CR��lJ�A�g���'/M�hu4lFI�e|{s���!�]�03.���̹M�t��[-pe3�ߑ;��Q�t���%}�E�[�nF�y��d�Z�wU�K[.�8*uش.��B6I��y>u�*���,�RW�M�X�{�.�_c%��e��H��V����V��K]�.�?��I
�׶����Y;����ӻ"����u�#�X��(�]���*�WoT���h`���Ml#A}�s�M�ȍ�ag���6�dT}�29sd(�L���XZ�����o��F����R(g��_&g�$�5F*��=��MsiU�Me�Ox8��ʰ���s�1$:�q|��o��7;��H��E��,}��ѹ6�\{w2��缮��%�9N���1��w,`(��>���D�9�H�;O�UD�J<n��سu��wq̗�4N26X��4���gx�g^�h��h���n@s�?���pFj��ۿ��joǆrE�_��<���k��������&�`�}��ϭ�C��^@�38����4���8��H�x2N�@���K�-Lk!�kOޟy<��xp�.3�^�z��r����E�x1�IO���Ŏ���%EYbD�ߥܝ���E�C�=�})X>~��	\�>|Γ��ޱRVj�a��s��r��M?i��.� ���(�SB���4z�HK6�Y%�0~S��*�K�T�$���H�+$Q�i���r~�m.M߀Q�U�<��;��=�\.Z�/I�W.5����|@�F'1Bv�E�L�F[p�o+VM� ������g`-GEf���_��|SF��!���a�KEX�[(k�\�Ȇ�3t�a6&[�J)�����R���+�X��*7����K$:�͂������[]9�5���F������ߢ��;��SLX�l�3�(����譩l���U6�a�0��Á��V��	����r�|��c+.�0 }ESr���-(";۞e��|�[�*��m<�Z���܀�
L�L��Q���|��]�P�a�o	V$?=��;q�E(�\����m�W�E�*�-�Q̷9YR�
���$�	`���) n6W�5:nSQ:��!iJ&����Y��i�`k��L��y�i�Z�y�CYa"Ѓ��V�8�ڴ� �c��0��Ԫ���/��y_C�G��2N�#��X�gq9�fNh=g9�BC(AnR��&��`!�������i���
xgnS!ͭ�V=ut���yVG�1���o�S�;�G�"�w;r%�ҚN.��k­+�H]��b.�R�'���/��0�[�G�Y*m,����.=��E��̗̏�����P:���@?,A�b�AZC:��i8X�ݷ�&��B[V��Җ��t R1��\l��d,ła���D�H�`��Gղ�	�n#�b1��f
��E Y I��XWI��?@aB��z
M>uq�Qz����;��ܑ�u����z�c���fi(ٷݘ;f�3�<fz��� z�r���裣\&��8�-��A����nyy�\�=�]�J2���$PhƖ �:��y&������M���͔{�-�La��ĩD��,��w������$P1Ut0S$�E1+	�	F2�L�}Mx:�&����b�)�� ���nw$��ejF��@�(���޻��H7�6�"^�1��p>J�O���(r($�͍�����~�+���&/	QR��v�%�D�t_��� sۇ�w���`�Z3'���>|�Oc�t��㦓���Q�'�=O��Be<V���C/� �_�䰴ј����|R@�NI�<|�N���JO=��%�#�P1����0[(���C�B%�t��V�:ҥu[Q����}�o�H��ItX�i��C���R�ɀC�C*����J	9���cyS�&�B�
��,x��0�*#|W�֜!Қ=I��"�Е�)y)P�V2�U��PN�7Q�P*�A�}�,��?�)@�]�t��܇�p1���� >�s��He6�^�l���k�{ҨBh���T���.~���|��3���{��$5RF# x2�(���i��\�:徔�)��oi�?d�-����Dd:��{�4L�z[����[��h��r�i(�D�f�)'��ßG1������r���p����Y��ּ��y9��^Ng{���� �b)e���t������@�3&�M��EE_A����UΖ�'���Q�֜i�E+�M�`Vd	g�%��v�2�!	�,��4c�r��?G��emB$jOɪ����RD�0:���; a×k� Ŷ9�W �S���|7��o(]zK�Û��y���1���h������hU�ғH��(���j�tr��O��e�	��Q�腺��N�d�^c�M� 4T��3H���n�� ��A`/�u}�1Ww)���F����D$�����D�� 2�Lsʐ'�����j[�kmz8��Z&�7y>����`\W�0�?p*�R���t�hx9�}��OB(�_��Nm>E������s��Y�@���D�$|i�#�2�F�F��]Q\O�U�Y�LɀcVH���8��'n� N�Oظ�F˟��"���Y*r|+�0�CO^�0u��:�lMZ�Qxj�Dȉt �:�-Õ(b����E�����z��9_JkЙ�4o�du�]eJ��\�dP���,�{T�/��(g<'C�/.��3(�C����Nʬk��.x��e�H��]j�V�q�j0�qH�p�9��J�.��=���t�sD���ȵg;G�@Q,=џ$cAμ��F���;Y��7�5c�dd���f��6A����ڟ���:2l�1��I���4�&H-��\�\f��C)�>��)��(A7h�䲓,��L����0�\�Y��5�Y�_}���K�Y��3XZc>)�(��V�@�}{�D ���{a�K���<,�eV��N�,�2~�i'-�j�ϵ�fA�Lm�/��j}	u"��M|�=�t�	F�Q�c0����(TZ@���#
Ѫ1aCI*@y�zm-p�yi��q��Q�M}�����sSu��G*�;P��3�=d�X��8T:(K&G��'�\B�X��;�CW�z��B{n'%g�jK#��	��q��Qpy�T��!�׆w0�{����9�"E�]ߏ��Ї��ݶ��v(I��MJ��Id�D��$W�t�w@�Jy{�צ��,�d$���5� �/:o~P��r��ԛ�\�H��Gt���6��(o{&(쎬O9Ct�QxY����i�9�-{쒪.���$M���r�ƙؓ(�)/�DD�������X������0Qq��$�s�xr��h/�d.����Ji��&�&���<H��X��Ov�;b��_g&��1jM�2i�������;y/2$�8|'G�U�G��vU,68ɠ�E�Z+��bS��I�Q�0��kt�h4H����Z��C/mi���z5�V��ŊV���5�Mo���ՙ��}�M�>�����!X?uM���u:����I!�_�����l������)��M�5;�(\}��U(C̢3'�u$.1I[�V���0�HZ�6�g	���(�L���~o+2Z�9���M�դ-��|Aj%�M49����dj㖯@k�"���Ol�
�ԔR�`gN�v��{)8(ɠǑV���R��c�.d�T���e]�Q���t�#A�_�eF!�`DE"\8�9�JO|�$�k�Ky1�{B(����Q�9S�y��ia�@AwI 0�e�,�R��
(P\fD��V�]`��ȍ`��bd�A����3�%�V���q�4���S�d���L�Ҧ�� Cܬ�v&Q1���w�������!I�b-P���a�[�0���(	����5:G�X��lz	�r��-�p�@-7w�2X�X~o� ��T�*�H.QNX��y��%�P��T�C}�SXd��{��dr��S~�+Ā�տq%ޡ0�o�Я��>��,�@s��,&zB�%�����0����������:n��#����m�gt��� .iHDV�U?�����<�_!��sH�Y��ڗ�
�D�a� &�[mTJ�~A���y��9�\,7�&��@|(�~4�l{�܁��X������8�KX�t�Cf"	u,�*⺐2ʠ��Ų���VO�x�H��*��Y°����xZ{"w���.t��c�AN�v%w��E�L�z=� ��ۻ"q2���������&�h��y��[OA����N*Um�C/\�@AqL�w0����/El}����P�/�KU]9���j.�l�T���	���V����A��a)�є��������hС�{��P�s`�����yn©�XD�I?#Q�n�W�% �'�'���ŅDގ�JN�ȁ�~�bݰ��:��� �e>4���p���)F5R`G_tU��w`���oL�y؄�n�N��Cw�Q��F+^�`��h����*Q�?�Xg=�����Ug�CY�!>e@Ɯih���EP>�����RsTi��X�ʶ0���;?l�D@��@��W1���vg�`��oB<$
��<z�)�H������ͭ3�*P�vDH��T�ە|L^���*S��QOk����d�=~�}���4�A��r�������,����-�dz���Y�����^달.Q^�C}�Էc�����6_M5wE{���re�;���.)0vmX��� �Dg��������2X�ft4˿	Ӑ�&�]\��%��$�O����|_%Vw&x��y��&A�E� �b��!q��4��1����bk�Ǟ�'_f�^>�.��D�V��n�Gt,Osi�¤d�c�Z�s}��V�ι�J	(��$_����`38�y輊9]�d�T��'���=�w6_�1��D}�\'V3�IbS���`���M��Qv�{O��c�_�X�s�Hh"�u�T]0!����^=�	KR��ԇ'F�;��iZv9��ju�mb4�P�T,)15ϖ��H�5��`Y�L=��r�yb�q>u��R4��c�@�,��z�`E��L�h[��IS��j:���+�~�h��u�vTY�����Y���-g�Du:���d��;;-Gf���n���l�_��`?�@j���e!�*F�B�`���*~]l�$\{�א-uw##�Lc�?�2v�Z���ޕ�]�ӵ�7�>�{ss�&K{��-���Ds`�Xj���c�{�OH�
�
J��X|Aq�ȇˑ�S��5��D�W���f1D���԰ō��0�ʋ��ʤ9f+���ֹL��.�׬r��ң��b "6!����K�XfWD�Q]��?a�\�f��\2Iu��9I���Q��h"�ec�"�\y�,��o���Q�1Q��X������;��J��NE�?��EW#��-�M�|o3��A^�*�������A:1�-�Q���L�Q=��	{	�z���"qJ���,ξ	mF!AQ�*Ӕ�7M��>&)���狼�@�1�I&�.(�C��\=3|0�@�%t:���B�^-�o���lXq(w��NF*(��[�C�r�Z�(�����)����'��%�/���Ч}��9���xEfuY��WnT����|T�:o��󝼟]]�E���y�\h&�pn���	8!���٠��4��v�8��i�+W ����(�1�� 3r[��c��V��m�k�v�X*`EW��ҧ���g�q���9[~�>�c��/�C���}���6)O�'9�,m�4�(�o�C ¾�UB5��M��A^}߹H�B�s��;��`^�V4�
�SF �Ӏ?�^�0�$��v�3���W�M�f6�����v��B���ļ�##	��3Bf
V��/ȠE*���r�:�ŉ�2,�-��qܛ, �Q;����=v&J�	�g,�rb�;�>���.u�A����0�u4�,_���wu��A���T�@�ơ\�{���Mj����]���#���v4*/O�l:�Ͽ�ɒ�g��̉x;p\vWʨ.�C���1$�@.�A��A����� ~b�р�F'A`�J�vT3	����$�����E��W�l~`w�h~^��,�� �ጰu�b� �qK�J���Eޮk����]���nS�YB�����x��G�.R���:輡+��_t�C����]��O'/�Τ�3	�M������:jZm�c~��I�,��qC�g>#����z�>� -�z色��;�^��P6��n�"xu\�lq����X�<t��eLƤ5O1���c���	ӈ�'�{��������"�7{`�%xP�9E�n�BRj�Q�j�,X��S�+:V�?j"��~�u]�Fdk�8����	�ڌ�6}E_l�/�\MXԾ)���q�}��a�&��v �m�7�	�yᲣLC\+ԧz�pvm�y"x��Vw���Ŧ.�=�}���%z��z>�^3�S4(Ix#��'�;GK;t��"�@�YEU�"gQ�拹	� {[	4���➳bY1/m|;QA_�K���g/�_��@̧�)���0EnT�e���	��m�WFꚸP�H ��[^�8����.l+�Q�U�ר9塿�%f�}#��4
�½*<
�Q�u-��_K��6��f"�iɆ��ßЮ��16�dBf+�D0s��柰)�����
���e�V"���*��'[H-��r�&�M�f�X9�KZ�����)rd
�$��;-4����0SivHZ+7�u�����Zs���0:�2%bDHBm�88g����F~Fp�gv�����fDS+�̘G�|7`�o,��gQ�rT��'(k�2��:�)��\Y��idoAO]��pyҩۘޔ��M�J�|XW4�b���g�fYn�;Y���!�+ce��X,=\��4UQ#I1�.��ڪԽ?gk�`�Q�)`�r�6�!>��E�/�u2H���� 
f6�yF�M�F�M�'�\-w�,1�S��$��cg��M+��DY�<����� �p�;q}g0��R�sυ����x�n�C��Σ�^T��,�fN���Zq�k�%X��h�m�����J~��q�H��X>�Q-�x��mB�j����i�1t+���26#�_�<y7,�By{�4� !�Ts��Vr�7�L�.�x�>lJ����
�֖�ۤ��7p,tuF�Hm���s�X5��@�����b!��V1�;��������^Ek����! 8�`�"�m�-R��'}���D;ƈҹ�)�o�2Ea>N���D��C�UV�"S�0�B6m�K��l1��m�nAdp����khܙ��h�XG:z�5:OL`��Hmlt\�5MJ�Ge���Oq�V^Ʋ_?�\�.�%�V~L��O�g�- �&X�����3k��`��
'�"&{1�ǌw8��
+̚b��\T~����Շ���0|*ЧQ���aެ����K��0^��EG��'���ע����p�y<���*�3HK�ef���/OB����E�y}IҒ��&O[�%)[�@��$?M����"�&2��P��]d������7ٺ�&�7��j^Q���Ds$�QC#�v�@3�Q<rS�z/������:�2$Ƨ��G/y����O~�s������3���~����遨�Q��K����c���߻h:��f�ǧ1K�T{�:)��$tH����,��u�^4�Ǫ��=�~�N���~T�9L��a�����0�t^/���I�z29�z�A�C��J�*�L����R�~�%����A&�ꓩ�G6Zy��JM�K��J
ȳp�kv:-

 9�@�i�i���@vN�ۂ��#�]KP,�n�3���Ǿ���°�&�G�|�@/�1�aZ~����ʧg8���m0l�^*��~���5e�ͪy�Z���!�W�b�)����_ѥ7��/�>*��d�·KA8hP}"��Y�rض|��54X�2�>$̟gS�_�̲x���j��%��3��e�W�n?[���t&��3������(8?�� `��j��u��ErY]%���&��a,|̡^���!����]:���u����ѨZ0Vzu���MS�w��~�=2C�WB�A&r�(���jb���@���R���,vy0vy$v��.�\� n6�(�=��'%��n�0SG�� *�1��T0�n�<�MA2��b��5S�rA��=���S��P�\�l���g��јs�{\>Q��ɨ)F��G�o��\:2�q���SI2^�z����|��̂�량w���3B��w^䏥L�Bнa�2�����f�z�i�<%GO*V��N�zL�Y�4-�6�=:�p��5��t��s\�p�r�������dΡb+��nNxR	M}�:#Ъ���KW�ɔ��9V�Dϑ�g�ldVW
Fz�hT���[��Ӊ�F�>�o�\��<
3�8��OpK'����I�V�"��e���<#�ژ�'X�m���p����<��|u	h
��꙲�87�̣Eg[ڝ��tt}YTw49PW�E���}c�q�����##Z��7E���'t�>�j,�RB�]�GZ,���q13o�����@W�~죔ӵ�a%I��V�\�t=�9�g܍��$gC[���{1f�4�U*���s�D�����a��a9w��ϥio�N��H/�P2>Z+����L�h&��Ep���~W���օZC���3���G��F��g����a�Z�ǹR�Î�g���A%��~�baEOe����pO������R���:�26�F���j�&��TH�M2c� �%�L8^������d�c����o�[�1����dq�p�j�h���P�2՘�T��A��sN��(	
�����=)���u8�9�;�=귰D�3��
�'=�f �����j�V��'3G����|I�q���������)�u̝z�*n��7=��]�y��X��nk�t����2]'et�Z��|R͇�F*c=��؄8�|h5k�R-7�E�-�t����g8�m �|�f׵�N �����kH��pE(p̓moB
B�m9���o� "�A�p(�&|��9*�W2�y�/Յ��@;9v�e���>��� 7���	�j��6�q� ���P�F{����I�N���l����a�U�y���X2C��8��@}���䖒�h� �O���7����Oh���OUÖ��n9V �~��"w�v�D�PZ����F0�:�lD�C���̕�&pDۮ��(�JfkȂB�y��D�Q�׫��a;~�꩝��|pL��j��F=���	���#r�����X��G�/��	���dX>�Π��#r�o����g��P�:��1V������!�"�k�:
�%?�x6�M�7$�%�� ՜D�;�ݻM�܇|��:4��X�/M^sh`����1uY�=)7���U܉�vĕ%N�	��Fr�MRplbto�����J3�ݻ�q�0�T���S���L�SX��`M�p*9 �IO`xq̓���6�(�$��@�ǜ;�J�����0t�M51�᪻�����ãnsԌ?�0�W�` ���؎�2�㉪���9�<f�8�q���b����5�`>d+.�K����-�7�"L��t������D��v,��{�嬵|.q��S�2)���8H�0w�@ąR<"^�#ⅽ ?&��8y��`J�sz�Ź�]MHk��������,2�^g?��;�0Ǩ�Vo����~��*kI��u� ]�r�t�����j�t	�g�h��S���<�֩y�HȜ:�?�N�O_��ч��8�p�ܧ����;!?90�],3��8�q��J���l�U&�؍�l�6x�{0s���	����,�m�S�w!���Y�%`G�2%�qw-���2��,˷�	k2�fr^��v�Z�`�5��x��tD7���0��俬��]LO��
����oI�����U]e��F�W/�U\��� e����II�����ˆK^:L��:�#�b��w��-��w#w6�ϡ����8�h���/�K�ڋFß��R`<{&r#v��]���7��[8\
�_���͙�~ٛ��<M��!�d�~� 5��ﰆ�-�Uf�+M�S�ƒ+�g^!��23c�[<Vd��L�զʣP�u��~�Xz����W��`�It��3��R�Ή��������$
���c�ɦ��@P}w�����k�`�$��Ы Gc(P��z�h�㯘z�)�1TW�0-�4��^	0>Ԛs�s-����A�L]v�Z��(J�#�TNj�
��-Į��v�Pk�Â�bx*��sF�L�RxB�q�:��Ou
���}o�7���n:,n��6��a���d�Rx��;Fߎ��$K��y/C��`t�i�������yv���q�J��L{���"Nڥg��Ա����N�b{o�Y����	�������[������ҥO�H��i�p�Sv���Z�����8�A��m��g�ԫ�hM�<� ۢD!Sm���Yr���b��L�	�t0��=�{g��U��5�8G[\�����$���ȍd1�6҃~�CC���O�������4��c�.n��.���D�Î�'Yܡ}��|�!�L6��|~���~����89�1��4H4�Z���e���w�ȶ�uu�]� B<���׬�a�0���ۼc�P�BI]�e�5�z�ݟy���%���|�3�'QfpT7����;�oq�s�Ke�,��@A�ī��S}�$gD�vd�0ս�%Wx�Qo|�������`��RT�ON^%:�+�oh���H#P��1�(c0�#�b�xungD{� ��i�HkW�9���f-'�G'��Od*a�O1�5���?���7So(z�Q��E\1�D헄e���[�SS�x$RS0R�����	���CN)ڻ'#,*?����ih ���i�N
x�{�`V�$D-O]��j��[��t
�w�C2	Z��,�p*	��l��+s@D�;5t�TE�'ک��[�a�ִ�>!Zj偖c���h�@}���pu�Yɿ�@t��� +�2ɏ	S�*o������9���L��l��o]�"��Q��'��i�2:����Jn�(��q�K��P_�c�7���&����D=�r*S�B�v�{AA<I^���X5笼[ޏ�e�ͽ��j���%9��C��ls���~iS���9��y2�Y��18��D`��u�g�Ȓ��P|/pNRaZ��mt��Vzk�xo#&�8ǍT2Ӌ��a.�}��V���ŝ
�s9V�k�����ڌ9Zx���f�g �oI
f΀g/VK����=�_�z3h�?��.+�-ͭ��.�<��SjJ����x#:%��/O��r��w.�9>��ޭ?�j����4M�uY��V�S�h�4v�ʠF?Z��)_D��n���4M��� _�d�=N.nϿ�,�ݴ3R�_L�ZU����_t��0>r�}���ݝ5\��r����o&��J�.�P	e����^��l�������B5s���k�Н]�C�z��Nze�~͆�E�*Z�
�QS�m��+W̟�D�H8,w�??f$�n�~��A�z�@f"�2-�,��q��m�		��_�ʂ���:�H�����(}��V���"v�";4� �]]0��h��n؀��	��q��C1CS{NvFDa�x^	��� ֱ���Aл߮40e�׳7)�YN/PpRdj
[�QeP'~���N��q�[����*���~�!�<�R�
��}K�¦�Ϟ6�[O�{��A����"���3Aޤ`O�Ͱ�c~��l�ª@D�'���T(����pT��{|��/���\�+��h���P-�*��� �l1�q�S���}2�*ΰE�?Do�P�^��RE:â�Ѯk�S{n�r@�#�(J���������2�2��и��zl��½����ġ�	��ic����MS2svKAJ�R���6`���5̵Me�T��WC�����j�8��T�.��;�@�'{�w�t���P
�T��]���z�Y2����4�O�Ř���ED��0:�����1�����R�E�9��
?tգ7���5���9'��\�Q;��ƈb��)1��^��h�v�\{e�%��|8�X�:�Tw�"�=�[�b����$tHsP8
�}���f�f
y�fN������t�i�;c�ŏ^��� Ҫ>F�ys�pR�29�~p�v��v�'�ֻ�/0㟢�҉c��~R='8)=û��9-��"�֘�l�4:�+7�(��#T1��^d�����繤��R;q"v��1o?]A�9���z�?v�Y٬��H�Ğ��鷅:?(n���l����3�%�ޕ�Q�>�Guo���oW��Rd-����ME.
�C}��.=�G�[�5F�,E�SA���J]g�U��6+ ź����9�9��Rz�T�?d2�Ř)��D$I�G�I�
�����pԮ\�`�Hး,u��N�!;K��M�8C�O�����B�O+\%BV�C5�u��#�gYl�c��1'�uj����>���D�Y0��e̫d(h:v={s~"0�`�7"�{z(�o���}��7t��#ͦ�`+��O�(�x�Qq��.���m���6��b�0�i� b���Z;,�P��6��YAMˆ�����Q�|�J� ���REp*�,��׹�V$2��L�/r���B� u�b���Ɯ�X�$�6񣮠iV�����|�D8(����C7t��˲���o8T�Yz1V�N�F�KO����@�he��^j��iX<��J��ák
)f�?q"�X(�cz��5�a��� Kw����m�����KL[`��[f0lFg0��}��#�^�� ?����.hV��Q������.Z�{�/��å�Ёz|'� ���=tl��-�0�����7wuu�+5?6
�r2!�J4h4Á�i�8G�+�`�Vw_����,{��e�f��u���|�/�؃8å8�:X���n�����B��nJ�z�O�d*|�2�m�<��6�}a�4�A�k�)��`5�XW���ұ�P��J�e�[O��@����S[]	B�~o7�2g�QBw52��Jὦ>�����Xs�vnNژt�'H����^]�l�2A�8ف�_����of��,�Ys�C+�5��"�⌢�g���c�!/z��)X�<��������6�vK�]#<�: l�������c w�+;z�������O;>��Ë����CSχ���\~ا�Á�p��_�C]|�cI�����5��d\!�-{$�N�݇�g��hoM�x�iͅ�H��.~)wG1�Cu47�4�~C,�\I�L�A�6T��`H�Z�F�ي��V�;�g��$|���:��Q�O=�'(���hF�^>��c����߽�����
{���k#mq'�p-���-)9ao�� iK��BN���Wo�-��ߋ�a���3N�'�}�?� ��X�l�'@�{k#��7uE�uѷE i|��v
�΃��}KQ��i&�)�JA�-r�2Ӆt^}T�aX-~����rr{��K����ށ� �����`�Ƒ��	��q6a�_�A%��Yߔ����M�&�'h��{n��7��Hr&�[j�J������9�m�Yv�������K�Le^���w��wҖr�+��4��j ���*�IvF"�,�:��/h�#���#ig�b�-��D�5#I��I��,I<kf�P'm8�>B�(�?�����j�d��y[7��
�J��F蟒��.�_�k��V�6�@oᑛ���0�l]��� ȊC��*�_�ǈ�� ��L�������Q��IyYr�<	]Z�V]1�Jm�R��@��P۾3���]"A�O!��S�������T���$<���I���9Kq[ѵ��5��{1;�n�G�j&K�OQJ3Q��\�jO�͢<�[�P`y�P�c�{�+���H��y���Os5r�H��"����q���NNϷG�ه��BF��)����'��2�����Ak�UȮ�N�@֨�`Hw%��^���S�"�ܥ=��^uh�*,�����w�6vG`w 	v6�[!����U1=�ޥ��fg�Q��_���b��E�,0�:�J~������|���O�:fU=$ϨΗ{A)�!Jy��w�2>^�;J����wzx>t��qwQ*)C�}h����C$(.�D��p�M�C~{qA�(��P'�:&��O��t��N�S��t汋�V�v���2cV�e����l/T����P�{ͷ�œ��<��x���}<��w��Һ%�۱��6L�?���7��?���o����"����s�wt��܋q�O#��Ln�]6\Sۚ ��e6��}��ceʤy��"�F�x'�y|�q&�o�"��jX>�~@�.��'��@�K,LQ&UIGrf[W|�`��Iu)���ÆP\+�Q]��F d�aRR�a���0����zr�E�5���}{Q�Z9���q��
�$���eU|xO�-�G�H����/G��y0��C��z>��՛���˦���%KA� ��n�-G�$E�T�S�WJ�T����E����>�F��
M�py3D�eV@�sA�tb�M�k!������8SQ�9!˃$��
�*V��*uɝxC?�8I��Ԯ#0��F_(��x_�֝���p ���xr�$�-��y�����5N��-
�,tRD$湨|��e{1ɅwĲ�F#��&�&��xղ�H�~x�m/$�T#�2A��f�P������W���A�L~א=�^��wQ/�)�Jk"��w9p׻_�'��g^8/��f�a]���I�)�P��c�W*f�� �W�R���x� �S-�<̀���Ve��� #Yȑ0�g�2eT�(������:W�����D�F,�,2o�����r�H��HJ�BW�<\n��aQ�h�2#]ڈ�Y�]��Hߓ��U|K���\�YQ�b�(V�?>��r~gHW���"��''�8�ևF��1�7�Ň�9^��}�kE-�����m��o{[sdFi�a�=�Tf�`�r�K�@u���mR�<d&+)���r���`�é�������P
ҏ�Ç]ݠ#��^���o�G��Av�:��M����S$�?R�
]Q8��| � ��MdE.2S%p�$V�7Fp�{ ��ׄ	,(�>ߕ�$MmB���"b#���f� ����^���e��AZZ�� �T�P"+Υ sZ�5�Bw����V�7�|�����g�W���6��	��t�^�mUo�����h?�]G�xm����LaRLJ'����'��I܈��,��
zJ�ߙ�w?�?�!�!�i+��%����*���'��"ӾNK�#�tt�.͝��I>�>/�k�1��ڣ=�̢B�3�J����cI��X�Ш�^� �0���^���_���"+7�� ��s6�� ށ�6��q��ћ�L�Kê�BcA��Ч��jb���%Rbԗ苿������8��Q1Ḹq��_�M�bM���;�hUh,`;ڠMD�ڡ��;چ�E����q�ѥ�9��nT쳲[�h�~	�"�?>UH{�*If�YK���A�X���y/
��C1�x�ҰȪ�thH@�M�޵�F!n�U��÷^{�5�'u�PЯ���÷q��HBv�:�R|���^����+-h_Z��4���I�$ָ�%̽�Z�!�ƕOl|X�~�ň�o�����}ZZa"c���Jt"?��d�d���*�n�W�Q��lt-����?J��,Ҧ��|�@��_�&y��1���� ��cV��G)�P���t�Fe9�'���E��4�f�T_�A
�~Ùm��z7SP̴9��.����f���N}h��Ș�#��Rζ��BX����F���;��ѝ+�xP(2�z�\���O����O�"�\����{�3�=�50�|����Kk�	���H&��ޑ�l|y-�i�5�w��X�K���̦Z��o{�lΗ�@Lٽ��>�!�H�&�R�B�g���MR�c�HkI��@濾}_ ��b��V���:�i�1ݼ�Wʓ%�[�(�"�"- �vw:���2���W�h�U���u�������.���>��:"9�^v;��<It�]V����T��o�q�/xKHC�_=�g� -;/�-0I��yb�8������@�����Ok�
dU=r�����R��U7���u ���Qʽ:�s��Y)UMy�	n�sg��+�/O^(�&����L���x��ޛ?�Z�*z�W��뿠�JG������C�U|�PB��m�^��K)^�f/[�R��D�p��F��k�q��L�����r<6	z?6t��~��cCj���N��Ç�z�w�<�y�wc����/�aRχ�ć��0��õ��p�+�h4���lE��/�� #^��D��� R�����]�(m�SL��a����`�䊾��9uG��i���c����x���;�׶��̺�]d��'����%x�7��1�#?����{���fLm�p?V�sq��d���M]d�.&݀1u��k������ެ���s���y�d���A�y��2��hB�@d���f��⢑���T�|I�{�#� c���JwapA�3'� I~�W�j�'��r�Z�� �jOH��r��?��$<�����X�_n{9v��/���|��y�x�w�-�#��t����F	���"pƃQΘ�O��������dW�l5\��$�����=�Xm��N��5�ݬ���3U����ppD�tˤተȹ��rE��[�LyQ�K�(�P��g�5�`�"%��=�:U�|��!� �JT�݆��;��A	H�(��;r��Z(	�;�����P����8�3�JēOg�l�/:e��ۢ�Zڹ'	�v�ɐU��>h��wq����7�D��\;O�fӀ�l�����h�g���/�=@��� \�b�"��|���dj�
�����OG6���6�eE���۳��������-�k���`�[PS�	���iX�y����k�z�`"/[�I$\nP
,����:�P��`c&R����^/xPO���>	���ؼƢs���/M��J;-]��9������SO�?v�Es qj�Q.�"�Gq�?�en|��@�o���"�Y��i$�Vր4"����#>��%̝]�(���8L|�z���X=)d!��
�`�}檛�ӕi&�QcN����I*xNZ ��eq��k-�ɻ��o�=�#����������;0=��&���y 7|UO��>+�n5�b��?��6v�{���e��+��6����^t9k{3�����W<�.���u21U`r��]�umUwYؽ7���'�$P�\������ef�V��WhU?�'oG�G���J��D�7�jJ3z�v���:zb��Lt�_aŪ;�)*�S�-�\��c*���n�': `f�0J��zeq@������T���F3T{-t,m*ʬ����녽5=����ݽ��P9�����XKw�Ě=�u��Cb��]�hl_��H���}�~7��Ż.���ޙ��nM�h�a�;�]���2>��S���zn��>X����Z��*R�wFdWY���Hf�@�?�\ߊq������:�	C�a�ơDغ�B5*���ʀ���Aإ��R��zɪq���%�M�����ad�¨��>G�m��y�g���N��`�+q���,��]�é]��Y�aF@�h�Ϯ���x�-��x��.���qY}�Է?�:�ʴ���M��֒UOd89U[�!�e�c8��!Z�33Ɖ���L+UnDO{��-2~3�C!V���K1�4Ή^N� ��e�{��!TT�Y>���8�����P�������>�{g�r�BY�iFl�q7=����F�|ۅaQ'p-܋�x6�ů�{҅[�:Ώ��ղ�dW�(0���t#T=�T�l�t��R�"���UM[
uw�b[%���0����e�DQ.��oI�]�X��w�\��'��(�"��`�~�5�"n�|K!��a�;JIN{(�~�40m�ߒ�r�������bWba�x�O��V���A����vf�Mq>����:�������r�'�5��A�b�;ՌB�
S�ӍԻ+ʄzV���W8����cӳ̍�^�]���ĩ��lK�=z&�s�UZ3�<�З*<@��:�&���-�v���:��B$����1(sX6�+2��fuB�`�]�R)��!0E���<FG7�<��xB
�9��$򃾻��S|�tx�'kg#���S����O��̿��Qu7�Ӟ��]a)�Yf�v�ê���\��9�C��#�����+O�hI�yS��~/*�tؐ8���	;������Q��i�ۤ��U+�w��Hd�[b\�\Y�8v��+�Z�~)W]e�߹����ҫ�ރ�^t7�P���Dl�6�<�m{ț�Aͭ��~��P6Nת�ۜڎ}ȗ �K"-yz���P�=�Ѡ�}��P-�h&�@)P#�oY��z.A�nV�]��A.Oޖ��B<;���W�N�J�Q���B��/�->������X	ڗ�5p�0u��W�y.�7t1�n�!�o�O)�������Ьv�hw7@R��n�i��IDd<����TR��@:����!A`��M�JK��>ѹ����4���}�kv5��} ��/�uq�&�&�km��3,A5%IF��,f�hkB� ��-.�k%Y����a�I$2kW�a�G�0q\���D�GD
<gdE��qR���7�8�R�^[�$Ǥ����^�[�6���������׻O��i���{q!�S�YV%y���`"ZS
�1�th �}5��9�ϋ%�3�����Uu�cC�=Z���O��4Y�uOygDn�6���	��V-M�틮hG���}�-�k�Lr��O�4��S�Wu-�սG9>T:��P;G�ן�Ȍ��w��;��C÷�J~���k���^c��
��wa���u6H��H���{{����m�o7;!b\�dsx�G{{��U �U?����'��^�lmr�M{@��F�E����]�j_��K��v_�'���U�ëpxgl&{��/p�=�0'n4L����E���)�Ɖ�g��ݣ�`c4�N,�}�S��~��p�44��0,���W�K��w��j�4f'�_hI�1{��(��D$��iyz�l�£�lxFz��ow76m�������7G�6���{Y���M��g�Y}qh�oE]�N�Y4Q4Ų������@�v��j���~�3�[#nƇ�gz�F܊?�=�(��7^�n� �R�#�R�d�FS�D�� ��[�I�p����k%�r�I��U1��	��S1<���+��P,׫5����E�6uS8a�\�_����+ns��yb��B�P?z�3��J׀�a��oU�jI�0%�yHgN�6�&~��hP4�F6o(%�H�6�A���O�.�c�'=��9J���x������+I۝���Vuwꅈ������+�w& ��y���������ƳA�}�]m�~��[��<�4c�ݚ'R8_��Ю�=	�m��( ʓ͘)�����A��p����ܶhɊiʕ��/�S�J�	c"�h���Pɓs�|K͏���S����V��@W��Mƕ�pxy�l��e����j�]�?����&�Y�D�_�m�`���,��w��Ҫ�� bT��V.2E����.�<[x�sp��I��I|�,S ��ӍYG����;d[�r��z{�|�\�I�A7s���"ܕ7�R���Na��<Ai��A���3����>0)Y.�f���ՑH�ۿ�׼#��+��|����`�$E�3-�堂�豉Z'6ճɿ ����ZUu}''�hUo�#�~\��['g�hU��:b�`�_����Фa|Z�:��Ye��[s��`��uc�G�zl��\����E�iSUxC��J[޹�b������&�J�6_y!Jz�띴�{������W�p���֡�|�\y���΁B�� g�й�p�Z��4C4��D���������13��7&Yb�Xct�\�xA�ɽ���hr|X��p$��x4��p�ݵ� ����O&C#��;%/7���e]�}1�0��U���v�Ŭ̠31e��]�J���O�ݜL>As�&[���@�6�%,����%br��i~�7�6G$�|�c��+}����u���)��G�]�q���;���'�D`�p�q���O�{���Z\ԭMS��h��>�Dk[8,�-(��S{V@TM>ݥ���[h4<
-���׳�e��\4�I�n���M��4je�*n�3[��U��i,��
(!�y�V`������ss���F%& �]&:Ca�����#v�v*�;��C�8���Zv�����|."�Q��F�ѝ�ײ;.���"@����䤍�{`vy5Q�n��|y)�z�Ĝ�����lz��&�]`�[_m�T�B��j
�� ��ְ(�V�įʠs�*ϋU��9�fW����Qn�=��Q>��7Y��#�=�4=�rIj��\`Cz7;~H+��%6鋶P�|��cؖ#{7��ӳe����.�v&tE3]�h~Wx\L6�܆�h��������u&z;��P����m���#�����������o��� ��� ��q�՛|G-�¯����|�ͰX����a�������joQW���o����aת+'(> �����?�z&^�^�~~3�7�Ql�z^�<Pq� z�I`�-.� p������\<s��J�	�j `ۜ�� �,ά6i��E�^��6*b�1u���۬�6k�b����qvxs���V����uJIڒ(h�^I���bW����7�O��:�W�Em�.����.�:,�Y���N@*&,74��q[��t�����6v��lS+(�t�[���κ������|��=�#"�����& �\Mt>�z5�SP%�����;�Б���]LJ.�c�A�Wb@~�U��3~6Fg;vDɅ%F+~{V��?���=�8O�s7���6�x�6����_�A�KKN�lb���Ďv1JP8�c��F���χ9�r��P~k���T�E��$�R�%��kyC?��շ�L�OX�~��;��#uSw�n�Kw��f���\;u>#��*�H�);�"�%x������4�kB�Vŷ�q�V8�Jo�
�S��ڛc;���N��ufW�����k$c ��Aؕ�̼���s_�2U3:{:�W�ڄi������=Y��c�XOSΡug~\Oj/=�83���i�w0)��Bߍ�~��]b�0�x ��ŋ�^�+��D� �ΨW�üy�W�K����>�2��;{|x)Vq�)1�ӾP^��3 �ڵ(������ԡ���Xɶ�z�K�bI���1J����y������D��`'Pt�G�*JTP��u���J�̯�p�8bi����XA挩{��}S��3� �afق~��֧����	�|\;V�H)Hn;6��r�y��;i���A��m�3NF)���G��Os���:�8N�z�gr�����D1}ȣ�UD���cI��)#!H�s��g��y�)J�V�i2���z�ٰ�x~_�����P���)��c������\�l���+g�Ѩ�#�O��G���t�w���g}�n+������o#��QCo2S��M�[�P�獠C�m��m��K���6]>9���`�s���<�K�{S{�y�`�X�����3�i��jz��]]<���1�񃫲��؍1��{6um{��~�ж�N��(\y�8�3�FA�addt��.ѽ�8m���I�p��M���6��ѥ�D?�};yG�i�W�E�ن�������S>�[�R�>��3q�R��O��?Ԉ�0��$��ڵ��ل�DC�tL�8�$P�6T�ŷ�l|�=Tg_'���h��ͫpa�AnF�� ����#�Z��n�Z�,s�R#>̓30tj� �#t��s�t����#�8�*�9��<�j���嘾��"7��/�)��:�R1��y�(0���2�1�����ӵp�������Cӱ(@}�v���o2��.*�ֈ��n5�u?m[�}����.n����Ȝ���w���Xd晃FFp��͸.�&�e'\��¸~e� ͯ�'ql�w�L(���1/�ʑx7������;��8�L���X�����ЦU�1��W�F]�P�/��o=q�(� Xl��_?����v����ېδ �c���<?��� ڐW9E��^�<]gT�iű�h"��b��
i���I������+�#��G穴����"�(;����6�M�gp� xD�Z��l+X�����\hT(RiATT�Z�Vd>��V($���8q�8ݦsns����� ~Aa|
��C�B���_�}�p{�������s����}}{�Q��ß���+��_8w@BO���x��r���������n�K<J�z��X '>f6�P�މ�.��@2=.
��M#_	�_.�.�GΣ��������W�x���j�F��n�:]��w���Pd��p�m"�3N	?��qO~K/��V�9)*�n�l	�h�۴�YZ��N��9	π��0�
`�]
`F�K���A��3qR��<����x�H�I�W�2������ vBi�?�1X�O�� �'b#�m��q�x�6g�ԥ���6R:��6g�&��@�!ZvkG��a��.zq�|q��]�)Qu�q�������<�9��c�<�|M�$dQιQ⠫��ǹ��D�k.�K�)q3+ys�M����˜��VjS_�YS�����q�ksN��t@:hS�P���٘h�������l�D����f�$:�5���Y��0~�n�Nہ�Ȉf�"�J�j���y������O��u%����?�MN<|�1p�ɜR�s����ꒁ�œ�h/߀]ɇ���n3�����C�����t��y����{I���=B�Tݫ,᪎e�2e�|D{�jq�xVkh�����=�H��6͖�,�翀��ϩ�2Y\���}��VN�M�t5/�%�Ko[	����>�U�Yg٧�;�V���l��)hUp��Ba��b���ܮ�ڜ�(�}N�06�~j�+��ں)��>�! t�цH" $�Ј��4vR��M�mN.|��'3��N�Qt��>>����L
gU�e#��w�o_�f9�ر;2��eW�!�	�x�:$���F��?q��拃����a`���C���T�.qBvα����9,�AS�"I<�/>�,��Vd+�n;(�[Dq��~�W<�<�5��*�\z����K��N����ٚ��@'��]���ي�љ�߼Q6�����D�jF팾�sV"/�oh����-T��?��x���F8���+����}6�qA��+�E��L�,Gr}_�e_���Π{MsV��1�Wy��0�9`޷t��=q?�����#�o�j 0�R��w*��8�E�/���z�.-��/y7$� ��R��
�Y�O-����K��T:qi���&NxD��X#���٨��ZI,�G{-�G������F�ks�Օ�����!k�xSI�E�nSh=�������[�i|�����w*�g������@3SW��I�{@H�Iy���Htqg�.v�K�6f��d?	w��f�C�S��>����"�̴���;[d_�6��\x��M��ԥ��6&�7z_�(�"�߄���]#G�l>M�VW�)������6�*޲⮵�6���&$�ph�?�P3V�[`r�=Ԗ�>��3�34?�p�����@r|bu{�d=���Z6:$�� ����Kt%<�6})��
pz�{�P|=R~V_�p��o�'�Mm���T�ֿ�x��VG�i��>`L��*�G��N��Tk�f���:��U�%��k^��q�п�۽���mq�"{��e9�'�v��5�C�=�<�F���w��NɂH}���2j��4�9�h��P������t��'�����J=�(@T�����k�y���{��,��}� ���e���'���s�	-XwN�c2o�=��X��<\�ۓ�>��t�N��gOW\�ړ0���� mO������N%�g d>�Dn�/�a6a]�}�|����n�2���W��zQ�u�x����7��λE�cҎcjC�?3)9aq������?KAT�j�X�&�g	F7#�aL�8��67������1tSU3jy���?���(�]��|������Ľ������,��kw'�O
�I��y���$�S�~N��L
!�������Ըo�� �r�v��F�wI��]Y2*�HG�F;D��w%T5����P����7���^�w޴��q#����m�Y���}��䋬7�xt��sV������8�3���:a�a�����agB��h+���	��%;M&���C������S�R���ڨł�pݛKYZ���qPh�v�v�/�#��@��w�9�I��A�V�>�x�����b��"nP���g��������t��Ƭ������v�=gU���tH��+9D�,��4�yu%�@���?�������U�铁��iDk�(��<������н�$M���8Τ8ݸ=nzq�������2��|C^Zo�{�ߗxZo��i�����mRa��}��c��m�Tg˟���x���m��������F���y��Q��`dC�:͇x8.�2} �B��Y8�����La�ei�@����ˤ:E�#;cŹ<S-bBn�����Z��V�
_��d~v4�Ez��v3?����Z���>zݝm�f櫍"%H.7+��ۯ���cпe���J���-�.���Fx�fYq�@ Z/Z�G��T���������������	��^]�l��ߏ��o@��V1�{���7�l0H�]���l5��6�-%M^�TX8:���_��m���"Z��7��"L���ש"!�G�����������2m� X�lPV	�a)�u���ͧ�X�MJ䍋-�EiJ�"�U��K�~š�g��x�e�u��j��c�0�����<�?-`���I}���Hob�QQS��C�����U�JZ���K��R>M�-	B�Xt��c���X	��O+qicݕ���6։�=ʼ)���|j��i�#�>�R��	5Q��V����� j��ȮR��l�5���Z����W�߉p��P}�nߊУ���7����}y{G��!Ɩ�-y��d���z����a�̕�<�7"����(<�q
�=�*��k�C��IW"��M����/I���dsF�zy��y�{t���'��[z��g�t%D?P=�_@��l�ǚ+�DX������ӿ��+�(,U����z�݂-E�lŃ�ng�Sjv�Ie�4�t��84�y077�櫷�4�m��R%���!_mQ0��;�+0�e���R��aÉ�ύ�1H1m���M�w_I˔��;��ƻ[�L����+ڑ�l����ȫ`���Bº���t�ضR��h{�8�͌�<$&S���C~F�6�mp���%��§~���Mo��-������5��y��t�.Z���CM���q�l�d>3�R�"�m>#�)����جH��%|iko�)��V��<�LX�������G��cr>V�ru[K/�BhQ�Ȩ��~W�A���-��߸�Jn����26l�8<��5X�Pf�J�U%*[̻�@�+G�_�Ǖ���o�^��G�Ū�~u�ʋ����\Ͳr���ϣ�������Ja�R����V;�͡r�4�(���x\���&��44��^�ϯ�"��Oio��
��S��3�#6%l����T"z��n2܀^N/����G��sAs7
ͨ%Y�Gp�≖�nc+�ü~8N�����$��ntKm�w�=[�F����pqJ��vrx��/m�O�Mˎ�<ą��R���}�9O�En*:!�����R�[���ڏ҈2IE�3[��Ȅ��%ͧ�Ckƨ��wJ��0��M�ڜ������Y9�U�'
��X���#>$���Y��%��K>4�kH.�S�h��#\0�8�r��?bd֭N���ee>�f�w���Z/��#��8�-�j�v�G)�A�x�>�O���{�O�fMp�
�~	]�Ac�g�m�mN���ƗǊ/?��<h��E�$F �1YȘ�?���;!+K�;6�&�q3�o��ō^�a%[	Ӆ����ֹ�9� JKs��f#A�?�t^#��3��:���X�+n��+��>�b����������`4*j�M(f��ޡ��nHJ��.���T�F+7��֨�:Ցv���(���i��r�ԑ��/��D��Fw��!��T�c�'���)�VG�Nđ���g��t��rD�N��G���J���?�G����K�E�}y��Nhuv8�;�����ӥ{PyTX́t�Y�!IM��}�'�̑��z�0�k �"���B5USwn���� v3�ޥg�n[�C�N����a<��V.^C��A�ԝ�K���a�ױv����.f�JrkcS+��"���z�i������@J_>��>LK��s�[�3�����O��&��T���|l*iY_C�5�ͩ7-����P;}r��|Ӈ��A!^u�|�7�0�r�ʒr;K1�HU�م�8��o��z��@�� DD8VM@�X�la�O�g"�5B��	�mv�IN���^���No3/q�`4Zǐ��U�j ˿C�)Aƾ���\;+zG��8C�]Zi@֐��S�ޡvu���d��!fG���W�-��9�.��(;���\��f��W�fa>�C�*��u���t`T��3M�Y�`�K�t$����w��t��v����<�E���Ld�I��cv"Y9�����%fw�i(V���)7+�:D��?���V�"y���,�B��b��*��_
y�:5'����bF1��
�kvKػ(�\���k\�y��C��@���%�!bOq������>��i��C����I(6���$�1>�L*�hJ�V[b��.jb"�����qf]'x7�o��%)��;���M�r�B�������	R����p�s�Z�R����Ӣ���!����բ2i��N v:���(�s��������^�����|A?����}x�c~)o]"�V	Omd"�Swh�;���/�gc�"�Xz��s�5�vw�s��(�Dz����1��5'�_��=�4�����)f��\Т�L�6[���W1�
gSz���n�J�b��Y�<�g�݄"�F����n?��Ao���F��w�`����FS�>�^�j|$��� �z���TZyy���7C����&6F�nb��F�9I��N�n"��s�"�;�ٱ@�B���񵸔|��^��@ZA��~O�>���Y��0�J$;O2� ��eʒ���}��2I	G��Ɩ#B4��k��	~���5�|PWky��<kY��inڕ����k��Y�2�V_�����#�i�P�C��"C4���6 �Tga�#���^@BQ�7�V�����x�N=N�~vD[��_'��>Vt��SU�GXi�q�1)8���t[k�]��G���;#d8���ޒ��iJm�Įj��[zVUX�<�_�I��y���%� _�Y�p���X�RmKL&+cDt&s�O������`��GA1$a2V"�I� "�\L���J��Y��	|��q>���B��9�b%�"j�O+��6�%Ha�u�K�E��6���C|-�pc�>AΝR�S���}�7$,#�%�}Ҧ�\���n��]E�3�Xoի]��ޑ<0�vč�"m^� �s_R�*�C�!���v�Exv�]L�ZѷsE+\���\����:�x��J�++��e�yr���ҕ֨	<
*=�5Cf�
>|�S�h�RS]=��s���*�\�y�	�ڠ�/9���v*!��T��6lt:cyj.oҨ��W4��NS��e�I��3=�ƮF�Z��k�Y���lBR�VU۫��j�@s���J���ۜT��V���W��վ�be���!��cj5��J�A�OhW>YZ�y�܆~���8���R�ae�Z�C	ϴp�9^��~j<�lʧ�F�![��|���7�M*��/[͂�MG�2����ڜ�]U��KB՞�4��C4�4K��h)���C�@�ԫ,�{W��2Ĕi>��>f�V�K�$�Bko3ma�s��-���V���4�����9U"ϧV�z��[��	ܺ�J_+�4ӵ�Nԝ�/O
8�>'�t�\1�1S��8%w��}Ur�������$+Y帢o�)���_��F|�*!W�����ŏtyh�~<����I���J�#Iw��;u�PY���3�7M-f�/�L��u�L�Du�Q���Q[��Z7��Wߡ���H-�"�F��	�)�C���H�aT�@V0m�4w
����x�_�9�&��L���T 8a7�oܹ��䉕��ѕB���$:滬�5��F�}���5�?��_�F�2hSkqkjd�D�1N���.�q�A�:w.U��s�v�dy>l�V+8�9E����5����2-[EJ�2O�6l"��E0�{�"��C����{�t�/~ef�~q�Hp���#�I��%�J��=�iS�@F��9�Bo��9�ş��im�ENn�sj��QZ+}�Ҷ�5VP��!��*ss�΋f���	A���l{��7�7n��C5�1jܛ�"��N�TϜ�r�����yl��R�UHxܓ�U��ރ�X�Ȇ�O@$�zd[�y^ǳQ"��9u�ZR"�il���L�J%2]�@eo3R�����V�d�K#��+!���
6��F��j��c������E����:�k:j�60Z�/ޡ�VqGs�z��~�xb�:��/��Ů�����[����	~��hO�ZC�j�~5���'�F<	�jef���� ~���&�����-Y)��E��q{�LT�ʲ*���!p��h �����r[d��:�����\;8��N�@w�
���%����:�_)F��tX��.�K[f�Hx�j>oP�>���E�1���|Sz�5��n��Vr��1|g�xo�q��Kw�����\F���_q`Z|�[fU���U�������й}���Y����0�|]/B�]� �7���g�k�#H��-�!%N�(�j����X*]u�/�!9)2�����J���&ЃF����ރd9�Ц��$⭸_ ���'R�ez�բv�a�ٹY���j�m#�5��k� ��}xQ�45
,U-��4��YUw���p<�g8Z����%�l����
f��e@s�Xd?�g��{��`>=�Y�����d>���|X[���C���F4�ci�#�MsV�
t�/��S����cm�/��?��{�X�b�C�$�
�q����I�E��6���m���v�1b>�*���$��-G�%Bd��C8s-p��ҕ5��Ʌ19Zr���ׁ�'R���!�Ix�8Qrj��uQ�2?�X�V{����+VK�L7gy���w�
`��/�$T��wpIl��76um��8��cI8��;g����Κ��i�ju�TG8�s��Zd[�;<���Ȋͱ�mW�Ȥڡ��k[~k�3;o�υNy����/�����~����F���1�jS"�:i�8��k?*���&��.Ԟr`Y���N����8B�g7�w���*hO�(��C�Izv��W��E񐞴��1F�~BHO��	P��,��m��;�&-�~�.R/�G��j)8t���k�:�ډ1.�yVZ��$�I�s	�����`OP�R[B��h�ܚ�=V��y[]jͻg����j�����|���Bm�~�?�mk�0�q� ��!���xx<Z
%\����U�0��gBtԲ�zH���6"�VeLS4@�*��0ތ�	V��kD��S	<$� �&�D�g�<L�:͡�#�$5�d<q���]��b�s����;�-ۙ_��^u9��:Uܮ���pV�gf�?�ƕr&޲�k~ƙ�9'�BVѐ��:~���O�b�ɨ+ٷI+�a��_M���&��4�J�:���E���'e�O���(m���%}�����x�$�?���X�xS\�n��>�D���ӱ4�=v��fo}��vjMډ�*(�B����·5��4�M��g�*���6��u]n���1��lw��D����o3u�(�ě��Y�=j�k5��F�������ND��_d�R��.������45����Ѧ�bi40%� ��}�BHO5��K��eAS�U����E޽ϸ�s��Ci�����
|�-hJ���+�`�3nE6�Sr?�ݡ��W�Cwx�f�*�H���N69$�*��a��S(-�:���ן��26
�O�&���C;Y[�
I۩@�!ig��5NlÒ�����S����#�6)�j*�=�-�!��$�9�E�F��f����kCqk��b+{��\���_��n��E�;ӧ9i2��?,�mב�M=�D��=I̍ ���+t��:����t�Si@�1���>?��3/p[��ih���
�dB����Cmq}�%L�w"ED��oj^�����J���>����Wipc=���qZ��ஷa���g�8G��r1��ԫ��d�G�Ca���0東&�hu�u�K}l���dG������������!�uߖ)��R^Z�쫘��^�7E��i�e0_t[���p�o�.5�FZ�yz����� mAV����V��^���_W��C/X��!��3�*��l/M��*�%;e���t��wٻ�AISw	{��ߔSC/�×-p����^�dV�t�E�Sé�Ju���D�~V���xr����򻦾4C��P��l������ȑ�1��]��j�|Zl�q�nB6{Y��M����+��*����kL�I1�p�4�ٴ3ὔ��e�y��R���3Y�_?gI�x���|�a��.���jf*}��-&fw�*�-M	��?�$�@�"����訁�h�M�%��BΩ��k�ՙ�1�t�����
M��Ø{��q�j����Y�uIS��x�7�zV��Ʌ��d��lR�/���l��-����sq���j>�<�����I�z��8	�8a'��ϚY ���u���q�u*��ρk$޴�]ӽm��ΰ�c)!���MG��R�/��%�'?�I���Vj��#.�/����9'�c�w��5��dL���3�8��a8���t�Ԧ������ �t�	ù�V�J�<�����o��
�(e�D��/1���8��%��2e�P���n�����Mf�ջ�/[�%�j�|<ʀC[OgɘO���yO��w"]�e2�u�����민�7U[0*X(x�҉m���g��`[��Hx�XXr�#�)�e��O�aY$��%����f�Y�_�t�a�c�*:�@}WU{���?a+�hw�X\���G��驍�b@v�G�8����
P��6f ��XpF�ۊ�`�j��-Ad+��*������z��@��^?3+�ԙ����N�7Nt����y�
�Ù���y�ޞ&���ׇ�2�c���@Jy�˄�'r1nL�4�<��f�7.=b�G�����#P��i��MSw
ڑ�v� ��x|�˳�^���ABe�e��W��xJq��C�?I�9��Ds�tШ�d�/_S��i�<���O�=�(J0fo�Zihǥ!m�q@<����~#'� �~)C]d�T:�Y��	vv��\-�����-}�|��CB�k�������^���Y�ҭ�//��Vv?i���3�Orռ���H%�/����W��~&��k��ɻA�I��w11E:���m�v�E+�c�����]ؓ���1�<~�L@�ăjgy����Vs��/�����������ٍ9�}z�83(������9p.AU1{�l�����Š7t&�g;�a���
����^�x�X����;���	��
�@��%N�)�x��O�N�E}Ά/m��g���^&�����W�q��v�W�� YV�^�RQ_l_!�,�z�\�5VڡS�FC����[��җ����6v .M��+��F��4��=Ź�f�ɯ�S"u
㗷��
�� cVy(��o
��!-X��X���#Z�H3��癷vs�BZO�8U�C�}�5��f�<��*8<�6,�N�r� :9M��;Y�����*�
D�n�*�7��o��'rH&X��0��S¯�&:ު�GN�%�e�kJ4��EʒB�,q�t�u�Ӽ^�������=�cS]�y��	�;+n�1�NԆ:	khv:�>�󅗸�Ԋk#7I�_����P���)�W���|@DOj��:,W��2�\�K6D�Oo��[�g���6q�I�M���NW��#7���#G�yǄ*����(|�r�g(�.ثD?���&�Um��bn{��ӂ�y̮��8�J�+�OY��`�����6֨�jWpy�5�Q�+��!-=�Q¬�-�bf��NĦd*K�¶���gB��'V(j{���m\d�V�����B�@VN;@+�B��B�����wㅩ�
M���=BT�w#��VYj��e�je�1 Z�Q�n�_�^	����I��`[�hU��\+��[g-�g�"y��g[E�Yfz�n�2�,O?I�J��y�z�"��k�<��D�P"?�&lC�sO����tul�JD��nJ��4�PjWK\��{c"I=/��)��a�$Č�1�&�X�;�͑��ix����R�h���z�Å���w�m�7���
�iW���A��f��1f\�%�������ʏD��>�
*�;-�e]�.V�`�^g+&��S�:$UN��<��+A����C�mn�/��D:�����uB��
F���U�Y��J.���ג�5ƈDӥ���S/'��P��V�V��"�q�j#�4�"�`�U�� �uek%�u.�H˓k|�;��QI�?@�H�I�iP�a1�'��D1�A��4䳛(��+O=����h<��e�@�kF2y)�x��F�U���6Ti%nu��/T���\�ƌݴ4��a�C��4T^���k���db\��,���6��H�0S���v}��˸7YO����z���rW�9��Z�R��\)�`���8�����/��t�y�����w& ����J���ښ4�f��*�X�w��P����a�k��V�iY]���Ʋ�$�L㢲�g����b��tcb��-��.4x �ݥ=�������G�vxܦ�%$ӳ�`4�v~y�0�SY�(˵�,���[�U�~}�R�]U��X�?�\�5ۜ�5'�3�<��(�dy�[�Q<@�%�.̐�:�%w\���D���_����YԶ�\_�S	nEy�V�E��X��=^;���J�+^�q�ڙ�O_���)IA�V
 ʊ��
�� �}��*zN@+���]�/����x�N]���������Tfh�K	��K����Ҁ��3"��w���y���v��!K=�?3^�\� _�TG'�b�is�R��؜d�f��9h}��Vv�����ز�_b��Igs�vM��f3-b�ył]����ȓ��1B�j����ಜ��AO�[�k��MTa���X�_�q���V�����=��97���%��OBً�a�V)/ţw�� C�g�^xl���\�6�*5�ͮ�/�5~���X�-j$&�?7k��8�%�T�1��Γ\����V.��u4��K���5����ͤ'ʒZ�䢶T��D("�S!7S_p�=<�m���0ϙ�����CKp&�^dS"���-/���R膺��Jx���L�2�Os%<��,Ft>�<��S��+5}<�q�G����A�1�ݦ�eS׵���/��Zwa��y�Z��Y=��)F����Q�� �χ���$�s]P��Xr��
�����ū��	#G�t�n�R �Pd	@����}�({�`j)��GO����Vo!��mL�+�L�*u�����2	�KB��>���x�'r�I�	t��.3".<y�.��~G]kR�짽�W�����Qۣ�J}"��?{�` r�ȫAe�Zh�Q�)K|���+g����	��f��Z�I�̼�)}���T.������5"�-����6/-WY�Pp���Vz&C�P7��P�
@`Q�7�j<��3 �\%x����T	���f)�[�Æ1��K2O�=g)�d�
�iBMY�n�6�C�gjO:���P�wOQ�Ca8Z��8}��0�����J;j��z7(�G��E����'��ָ�߆tk�8:��9=�R��6GmQ~��K��v�:<[{�9�����K��)~��v����F�O�v��R�e�`#ie��Va�c��K�hRnaʒ�%kٕHEO���nr���I8D�t��K���g��f��x���:��R����ѫ�~��_��|LL������F3�ز?�3��#q)P�+a;��ڴ�&j}.]�V�����O�ҁ	�	�'���l���H��iv�r��Kħ����#�ڢ�ϟ&��|mj��6�*�6_w�a�V$���D��7D�h�g�x	(j%�	_y�ʜ���l_�	��
sXYZ��`��F�e"�k� ]Ψ觝̛���C���N�^3�.�aH?��)<:��6u��iC(�������k���ej����հ�ib���]u��W�����p��Pvr��"��Y�z��"-�D��O�:�y����`���
�h�%��1u��=������X4�-^+����+���o��/�`���\��!���h B��X�%��2���2��b�P����S4�	���e����nd�n�m�C=��-�c�A#Ԑ��mY��3H`��P��0'�eo�I�{]����OHٲ�~&���_c��mF�_�5��i�_����[�O�k:F��`��n��1DP%��[igPb���	��̯�"������+�mگ&�-�4ת�3�,��	s� ��i��Vm%v���1�QWwz���=�A�C�$����Z�q?}����UO~���mqeU��D�5W�േQ7�*��j�ȓ�n�i���z���,R����&�-خ̝$X�	��a}��F�5j�E͢A���ʕq�Cg����I�T�-��Y^�����%��,�pX������� �~��U"��xB�����U����Mx������JOl\��>�	g���`Ɩwc�\
�ugg�=I{�;�،����ԓ�`J���q���������𹺊����,�/_>��$��,�+��n|ɽba��#���#�R	�D]/4�=�N�B�fY��+�xD圃����f����Fb!�B )���EbV����YX
���t��8���x�_�1 !� R���;5e�1��I��1�7�(K��6��lh}Z݈!L����XI�G]	��³JOu-�Ԗ`	���e�k�ډ���6�Y��ڕm���klԵ���e~���%C�p&��v(�N��{�ό�VGd��>cĢYh8�Ӄ�R�j��#�!�;�L#����k���i�I`�U��!�9��7��V�=G�
���\"�b��G�(��Cp�&���|�&���tDnA���01��^�g���?�D��c��=����d�[�o�;A	WY���l�1BM��C��a+
��$_Ӣr����P��ڟ^��Xh����+P��$Q@�[����x�\��w-�7a�D�M���gzO��6�Ɩ�ڎ�B�Z��z	�I#.�oU�&�Z��#���|�,E�;T�>J�յ�2QF��).�x�I��N��u�e��S�UO�j��H�����4h�޳�u饡��jI����@2c���B����4��K������:�䐟�:�GMYz�@e��B�&�,����wu,}��i�h��#���s6�۱ �-�����$�d�`mͿ�w2^�6yhV��3��)�\�X������0kW#^�Kf(#��C�V��6#*Z��rF�d���^�H>o�Y�Ո�| CF��|*f{��Q"�ڟ�\c<}��I!\�������$m9�S�<�����@zz)0�8� Չ,��\ X�=*�#��dl�z�4+dX�=�r���m����h��S��ɶC1A�l��ЁQ���n��l1�j�Bh0'i}�=��_F�ۉ�5I��jٷ>M�ÚL;Ue�V�xa�u��=�:��/�'�,�qF�sݝֲI�]5R�N�G�T��}�)=�Y.w��-��Ud����-�W͏�0T����Z��p���H�
hK#7h�]��H|z�6��/��hɚ_Xv�#� L�i8`+h%|�
9�۩��'zr�	��@�A;����I��>�֛�f�1B:��~��&t���#��G1%���RfR�ob�/2Ti�:�I�I�[�^�I<aw�zGh?Lř�s��H}4`�O��A������,d����>oq)K*��h^�y����u��d?�E���M5�9.=��cN?L��lv���čQ4[���BP�-:(�~�f��=صsh��c�%S��y9S"m�m�Kg� �\%��*5ͷ��Xन����*��7�R5_=M�R������Y��u[�zܻ��3�I[�l��)��{2���ȇ/���� �����[��;�o�
��b'�%��nk��spr�Hj@;�[e�`�U :��]���X�@u�V����L��ᭀ���A�C�n��ҧll3�,�6¥��`o=Ϥ�j��
�2ǽa���qk�j�w���
��*��i�
Ts���<����:]y�0.�~#7X���TL���aQ���`�?c>q����ɘ�;�U8̭� �=��mH��l���=�kq@�$��V�b�0�h�&�׉8�|��~OOZ���xv�#�s��X��\.;��4�.�h�t2�<9��E[��-W��d?�=\��'�ۛ���}��p�G.�goO]I%|1����������g#�y�E�,ur���q��ԄFW�_S��	�ޤE�<��O��f�r	� ���ʖ��S+�c�?�v�4�}��@�ə�$����-�E���6�����T��ͧ2ڪ��_�W߄*y�f���sq��sw k�$ҶDCXw�oj������]4'mq�e����7.�����S��m��fD�i��?���c�N����]G���熧k�f�.�>k�5ϓAuy�����������D;W�L�N�e��4)��cV��~I*R�gtD�ڦ�S�� ����Nm��Wq��.��@�\e���c�"/��~�nC�9���Uܞ�4��S����4L�;t����J��p���y��tЎ�;�t�a�?�K�n���a���0�i4�6�I�bќd=jp�c�%G{�P>:�,�ɶ�������v�kN�p'��DX�z�������ӷvo���;m����ls�T7���i�+QQ������3��pO��IE����$x��!�3�Q�L�ÝZ6}����
,�At���������4����,���-n<��t7ÿ&y���+~?hV�mi�&�V�k��FG}���i�@B}�E�q���}�Z0�5��4�h�Zw��3�׉=��"F�g_��n���'QN~�z�.�����&�^_��&t�xA�x�p7X>�z�?߬���Y����ϖi�B���A{����c\�z�˵��;����_X��l�����㝚+M=6�6��,2�l��l3q�01�yw���	����v6y���2�Nw���p����Xh�:"��O[E"M�<w��sy�k�r�7Q�>u� ��:e.���ف��ǽ�`�;��w��U���@����x��x��K&a�,��8C|�i�[���;��c2��ݗ���3']����� uS�`P�	�8yU�t'�,�ie�eL��5�2P��/H&�<����N��,����Fo>{�!]��Svx-��0�Y�pF(a\^˄��4a��I����,�s�x�¬�j]�gIt^j����B�7��ƿ�vL=�1.w��Xk���K�����Z��<u��I���Մj8�A6�}`��P�81�	���(�g���t�>�U�Iw?I5�,�u��9��⍉}����
��$_�4�����m���]�ƳQ"������g<K 3���(�8�>��\k��r��\κL�f׆Y���F�,�졟3��Z��dރ(g��4�ZY���L����L,I�<W�7HbzL�MH.ڙ;d��A�:�֯�nzh=i�h��D�t㇩�I&~��c��N��DN7)����C�Braf#��J�M/��uyOi���#�s���S�zg��ؖ젣�R��������Q�m�oKG&��Z�DdHI��yR8����ס���pr�j�W��*�"�\e��^�U&X�6���El�-xH��S�X���i����z�J����϶_P�>Ur����Ձ�y�� ޗ�@�˟�*�4�FRKXM�G��l��˥$nSw�>��8jxX�E���<t�?=���<u[��&�r��X򍝭��T��G��w�G����N�`���oʒfS@�ل��=x@+q��y)J�b��!����5�5Vp�. ¹�B�q�ձ�V>~1[���Qn:�V�����cy��֦��7[8J�և۠ͦ�[p��!r�����H����!,�����B�NU��$,��|6�e������l�st^^�\N�!��&������~�"O�N��e�~���Y�ka�z��W��2������M�U�{���v}X�$B)�Ӎr� 7�`����xL3K���i��qj�TBr_G�H����t��n2ڍ�77ɛ�y=����I}�௡A(Җ�QΎ �ã�_�_�B�:G��f��B�Y�����7D����@-���P�����ٜ�z��-U�{x��Y�N���E�&[	�'�m�������ݍ��N�'��3��B\�<Xrq2��%}zr��7�[�I���T���	�6�L�CI�=n�֓��V2��nd��Q����ҷz�@;��|S����ÎI�nlG��j��x�!a�_MNXr���x{J){��P�&��1���)O)��/_/���\��%L�nhG��FY������܌A mD��l,�r�"�Q�ׇOP�6�i 06�Tw���Vt_������������0 �w����Yn��9>��Y0w�����F���A:(Y�v���&�x�6ܩv4|i�&f�ή����6�Dh&��=�(�ZF�i˄���4��2K�\=A��Y�p<��ج7L���
j�'��<�ښ�8��[���LT����,�p�6N*R�S��E(z�I�M�ϊ"Y���DL�n�#����c�Y��f�П�9d����i}�`��&��9K�`��辶Mv�-�	�.5M�H���|�	��<�,�CI�>0������$ ������f��é�:�k�e�=�'ڬ�����|��W������S�4Rm�]fe��[wJ(0�j��9+�u�sZ/O
���1~gh_g�Mu��=�����(�M�Eh�4Y�
%�𢴄;3a��^�h7s6�
/}�6�!��d�M�������H&�����S�	=�x���+�"�W �'4�̞I`
�A�~�{�_��,}�B�<~�z���	"Kf���[q37T�ѣG��yG ������߄,
���(ksiL�4|M'%'�`�v�����Y�]y6�����
�fmp��d2A�#�L`{F��;��ן�(p�� zHh)��'f�#`6��M�Y�_��l�x@h5��qj.;(�1}�gq#Ϝ�D���t�/���*lp�������8�� X&3�FY�p�66~�0=4zЃ6��7�cmWsiG�#�p$��M`�c��vY0�[0>�Xw�-�$����ڌ�H<0-57��㫆�e��Z��;8	�pUp��q;q��}@���{�����h�[p[��q"���Gуe���j9��o�OպC��g�u(����4�]���p5�ʄ�f��mB#�t�[	�vXj.ga6п�(�̨�I�Z�vק��qX]�?g��z�?�`�L�I܁�" ͽ��+Ob1�cz��w���&`�"�`)�J��j/y����.����}�#HI��2I岁D���$}�拱NWS���BƋ�O�V���W���*K7�G��m�&��Zc�فr�J�f��Xp�]���.�iTuɯSA��ʘ3A��Ͱ��E]����Fд?����D�af��a;��l$�0�9(�P�ܥq:��W�����]�9�S��1~դ_�T�<|X���h��h9�͜x3��C[豰%�����QBG(� �A��O���D��yO�@�x�f{�f��S�;��(M�̛Y���3�I�(�o{_%�[��<�cY����]d��3q5F�td4�ݙ�8a����b��z�+���j��䝠he��C���=�fč�)`���?��ٖ9�At�/�^���Ɲ���)��R���gk���:y4�|Z��jO�D�L�jsv����l&�fz���x�D^�EK�\��^��@�L�r�ϴ�z�d�rZ©���?E�׳����Mm�W�:�	c�Vng]D��ob�u�V!��AN�2C�����w  ��SU�#�r 5����B:$$4E����z������ۣ��x�����D˳�o�h��2o� �ˏP���WI�wB�q�Z��w��c.���g�-���{���POͫ[e�S�b�:��}ަh��&W3�#��B���}�{f��5C-v��\R�=p1��[�3q�?���ѳ�5��x>��O����|�aF����ԄuB���-���z?ܾ�۲�$݊;g;�8��1?i?C� -�4S'j:�����O��P�J���3qfq�(�~5���=�f�����ſ����6,@[H2	laY�rk!�/Ν&�9�9�Y���d�v�2�T��ۼ{�Z.b�Og�7Jx�@�6A%}w��Ke�ﻇ�������hկ���j�g���W�ː]�׍�n:���S93}���`"e&�'!$�D#��H�pu�� �=!֣�Ppd~���pP�!y�u��3#Yb���U,�=G�ˍ���~m�E�qt.Re�9��>����6(�O�H�ضK�k��4���H
�^z�51%Sԟ$����kA�XҖ�6%���3	o~Ր��I�G��R$Βe���2}߶�qa�彠��:��@wh��j맄�7M�;XjA�O0�pn� QmA}�&����b{:�����!F��u�@u��pu�Ū~�ڟ���0��-���眱b�G�����M��q�7������2K�m�!�e�:c;r8i�x�ܼ,�E�,�����-1@�p�6�wG�2K`��d�-�����8&V��	2!z�WY���/])K����4>�F}9,�����,,-u�}��@7�x]9H�
FI>���"9�'ll��[$E�qnm�-t 3�1]�n������#�e��o�p�}Z��P���j��~�zCl�T	�)������Y����ⴍ���H�F�B��)��}���W�|z�+rEo
�~�qN��j�F��R�6Ү�ҵC-uh#�j�S�RK]�H�Z���f��F��>h,85<�>V�6s��F����K�H�m�����O��h��ő=ڍ'觸����x�4q��d9R��%ڙ��"��`i�~�s`\-����Gg���ɻy�R�gI��YC���s"e@�_��L�$w��	���C�U1��lu�H�ew���ɬQ��)\�f����_ZD��7�<7�(��K��6���g9��y��0�Z�,����	j����<�{�Ǜ�y�|�ǭ�<�*�[p�ڹ�?�n��#޲W�w'��xNw Y#��P[?G���Q���d�A���FY,�V
�'< �m��.'�G�G���S��w��ە0_xw}����1�r�ˢP���{�Jy��%���)i�bh��w�2�6Z�c���8��3¨_��#�'F�yu'��Mz��S��bkh-9�[���V��$	6���f2�Lj�|f5�'J�.d\Z��B�G��X�N��k.�ɿ�ҍ/�%�
���)�$U��Co��]�p�'�`��dR��B�c�[��̀j�w��4S.��8U�Ȧ�_�H���e�7�p������y�&M�=��'M2-�G]����F�]�/��6�K�x����c���q_Pd}���8�&q��Xqc�E)M�'^`2˥����7�.�����g	.��}}��[��#y����|af￧�����G����
(0f۾��J%,��ݞM=%I:D�b��52!*᫯��?���SZx�U$�A�� �a�=Y�-x�S&���;����*B�{-�H�۱�.Ý���A,��_kx�~��Ѷ��<N�,Ʀ5b,,����TK[�>�(��21Ӡ��D�Rҿl�p����g:�W� �/���֚�~��	�<NG��4ǳ��]Z���+i�]8���|��6ޖ2�.V��d�\���|��x��_ ��&�T?%L9��������"�j%�+k8���KQ��yF׹\'�+z�{E4�2}�Q��K.d26�۲������y�1-���q<OO}.���"�[��f#s�����F5z�	sEu�?asr\<'l�":���H�G���2V�2��}P�:�����Dz�oG���t=2��$ KT�N����yz|�ܴ��u��N�3�SJ���澈:h�L��DŊJd�gC�TK��d�t�=�H(�d��f�d�rv��~,�.%�vz���dG���Jos:��G?��7Y�ѱ����S1����P�P�Ѷ�hZZ�֑M�����X�v�gC{O�5=���OOftD�:�y��R��N2Ȍ�f��Md�Ӈ<��>����6*j^t�W`?~~�����[-5ݧ�4=�6;��0N"��̰l� '1'���|���䖖���e��i@�!ζf;� ��\O��Mo%;�"Gď�GN�El��?٤lŏS�LI4�E4���sg,�|��P+K�4�?VS�O���6Ld�]$���|��������m�9m状|�z�3q}�c�G��:�
�)��r*���>7�� @�]�Ǜ�g� �<C����Z#ʼ��&�M�w���Kl����R�n���L&~c�t±p-E_�&C�:������ �(p�y���Ҵ����X��>�c��e��AΟP��\i� ��|�^�E��y�?�Y�}�֐�z�I	.K!Ȏ��\�W�(����gBf�����M��T!lE�(6�;	첮U�l�*�[ݥo`@V��~-���ײ�;��F�����^�	+ �L�}�)D&�Gri����e�uڴ���A/��Х����G��*�Y􃱔������H>����q���
���k����6`y��
���t��n�@�떕r=8h���6�)?�����eC  ��xr�SZ�;P��l�CYz�=t�Jeɯ,�=R��-pim�u��~p.'��fS����Q��h߲E]�w�W3��&*�	+��W���_3��VY̋��g;��a3"�n$�.o�Y�
�*g�@����e�n��mZwe�/�N0SN�+��X��W�.��J�F��&�4O�Ek�G�����3�HBª�:P�A����Q�>��ҵ�F2^�H+�ȗ�~^�Z+j��oI9#G	g	G�|Sv�ƺ�C5wz�T��6C�טZu�r�hIS�%�����Ї��2��=bu�Da~M;��bƠ�VB�u��p������v���u_�L��T.����9|`����^0�����+kT#��'q�O�&q��/;D�ڴD䂈��@U���ӹ��jM����Ǽs�q����֞q�/dFI���H��G}E,���E��`HS�rF����%��R��+����p��l6�y��ì�m�:����`1�����qIC>�\Ir&����sFn|���bE��0�zu��N��N��[��i����kvzeĦ9B��A�l���Lȋ�Ԛj����!SK��7�S��? TK�:/Kǲ3�	}��j�������7����c�_~�_�I^ba�,l�&��3�-*�U�["G>�*!ҥ�u�0@��$W���ĵ������R���x ݽO�M�|P�`gԃTS���Fn�o��OL����3��˂�Dd��7��#P�dn�&6�}(���k.�d�D!�����q+�Q��?8+V��o��6b�t qzW�&%��4�����#.<4i܅b�` ��N��U�`�&o���K�b6����a���;r@��� �?a����o��UI�V��VJ�&V����75�d�z9�2M O�g�$�#ɨ>��F�T��Z����e.�G�������g$Z|���4w$裮���}�2{Ay�^<#�,���%�ϰ�)֐h:���B��G�ݞָ����m��&x�sVI?��&�e�:j�I൘L�=�Ff�!8ԃ���{�AD�F�@|�g��ŵ{�H��n��+�y�+�Yǭ�l���-7�-b%"��`�!#T�����*酂�ne�`�D�w��Ն���uSm�%�\	���K���a���@��L����"�*�g����y�ܩ���}��o4�D�Q�^Ǯ(�gH�ge�=*���4�گ�k����'˿��D�o�p�]n������
h4V���o�/��K 4��V8έ����(0�WG���DѥIIΜf�Vl|�}N�k�0����VT��}��p`�jn�8��X�܆�+Y�oc���*S�t�87&��	�vv���X� �T�[(:w��H�#��7�rc�H,���������ݠ�XΦZ�������9(*[t��Ͼd<�I����1����i�D���>ΦƋf6�a�*���F��[�5я�d�S�g�=ڭ�l �Gd��������RE��z��^C����V>��B�YO�Q�6G犤J�KY�#r$P��y`��n'��k�\#�Jrx�{���h?�ڧL��,ft�F����H���(��E	���iC���=�PB�����,6uHna�[���%!Z2&�n�4�k �V�X�i��=Y�l�Q�N^�X "+ХH��G�Lh,Oz��e��>�M��>J2�-�&wr���2��lD����y"�/�AÈ.�!�){VZ���CI^t!Y�Π+�3��\ ����d�)`��EF�#ӯ�[�E�����ɑ 嶫��ǟ��1uM1T�(0�"���� <��.8�,JAh�*ˢN%�I9�����Z̳��l4l�Ñ�Gb�.�d����%��@�Gs,�sz���MΆJ�!��K�r|�b|t�����ng�u�JSg��^\�65�!���[o�����J6�,��eF/Z�g�;4�
������D�@��E/�z>�k�a���J�200$D&�2}7%�g���c����Y�q�r��T�s�Rs����ξ>���{'Y ��	��U����PR��T���"�M�T���c)F�ʮF	!����H[l}*��ڧV��DTH�$������Y�H	!!�{����l��}���O��s�Ν{�=_�����L���*��FY{��/;���y+}�;�
t��a�l(
j�
}�����Y(�1߲��X�g��� ��kj���"����[ c�B�1V�|l�PZ.m����<\5-}
�M�[S�)�r�JK['ˏ^��{ٙP��e�H�j�dS`�������j��>{?�\-]����D����T������FK��������Oo�0�p�`W۞	�s�(|�1���N�er{�i�j�%�_���r����`T��6vm�9e�7(Eʜ�c�����CVX�~���U_W��ÝN����Βwnߧm�m�f�
7�3;xU����A*�<�<�kD�(֪e�b�����"�W1�ռ�[^���wiz�aX�k�۔ĻG�p���J��Iu�ZI<�	f��a����BLc��{%P��Ę�P�~��A��{�� ��,�����ї<.��՜��0��5�[�d�I=��k_�b�{S��o�mD+t*-{fV��LT�l�u~�.���!�@��h��j��}Ԏ�	G��;̰�G�ަy=�~ݮa�_I�ac����3�z��[�+e���D&jKG���c���Ě����!�	]PO~١x��6�]+��f��D�u��=�l�7�������F@=�؊8����O5co������������٘��Xu/O���+���t<)̹S�q��hl�!�~y����n��<�èV�e#�~K���A��EfX��@RT��- P�(^}��M�#zd,��n�&ɼ�p`T��3�|C���^
G,���&-V�����imYΊH~�:'V����*~��7��M���<k� �+>�`�����s���.V���y��������u����[�tse|(y���_�d3�<tC����3^o�rD�3��ޯ��x�gF@���&Q�V_��u�my���k��yƎA7*�� /�d�̏!�rq��H�U�-�ަT�R�"N�c`΢	���#Jj�AV����ٱO�8�W�A�%���c,��dt��Vj��g�Zy��r/LL/h�lp�<�b�͌�	�W�Y�jn'C�4l��J�r&�ї�_= �����+����d7��/���̲��[C�d�aLY֘jWI�� \�GG sB��>��#���&�̘\�m�ަG�V)�rȎ/Tt&D�����v����<Ԕ� E��vD�o�φ��'b��)�__�_k�e�(c��"���+�_����Mi�;��5Y፞�t���1D�o�w���m�d�~\��z�*�����_ڭT[�G�&�/�C������Y�����&�9�<g�l�)A>Si����P�����3�l3�`둸��5(�p���eV�ez��4�#�������L�bU���{`�J�����Q��4�=�"2j<&7��s�t��	|����za�s���o�y����� ^��5nyx]&�/Y���{ ��w�Z���I�AC��߷��C[2�al3�ԁ�V�.�4��E�� ��RN{��L�e��C��#�i�נ:Bi[��6�"�+��9 $��	��r�Q"���]����:��uA�	j��G��>�`\�u��~s��ɓ�Uڐ2���Q!뻷Wć(&��i��h��FI[5���M�N�_l�m��ed�#w�t�7"�'�Uh�/AM^}t��s��K�J��йD�9;g�<t@������� ��Mc����]���Ͷs���ܚy��9Ŀ�f��p�PO��], �C�� w�k��~��	��ۓDK+n�qU�6�*�$aC�٨�,��kY;I����'h��ܧ|�7P�L��P���y�� Z�,�z�D,�'؝Fڜ�,�آ��%����j��Ni��Ͳ��v�{F� ��vs�?�/��> �=����sHl����p����y	�����5��D�9�-�����F�4B���[ۊ)�'�VJ�����{��KM.#�x�ځ�-�Sնf�yIB_� 	��Y"�m2Zu������v㽸y8�,Fk?�F�]PL�m�_�(!�""�m?�*�J��E��S65;
�g��:aw�S��(��e*����٨�1��x��f���Q�,'����}���Z��0��S��D��j����_+�{��4�6~�&)����C�4�W�������&�9C��֔���慈���X�V�ي���#�l��k|�֝|ll
��k=�i��NZ�\R����m�n	:��j��|��9J�s�+�|ؼ*��mf��M���/��f�	�9z(�k�<�L�Q�w�A%<���;���P[�&�K��:�������#��33����䅡w�Y�v�yuk����
;��~sx�Sӗr��.��%�*��t7��#q=��`R_sy^G�(���M�e�F��=�-�5�FY�Q�M�c�=l�ֲp�#���:��'�⃐�~F��"�Y�*7gՔ��.�n3����w8qܢ"��<�������[||3�������3g�ǖ��S�+�'^��7u���ɲ<_+�5�������x�j����1����`���jd���~�xv*���^�R8��a��0�b��(H�&���d&ޖ�_��
�C#`����f�7�d��l�Ǥ���W��"�e�@`�A��G}JI������;��I���F�ߗh��D��I-'��O�5�`�v*���S5�]h������[�Q�<(w���>�|��eO����p&b�%�Q��Ǹ,���kT0b�rm_N�z��-�pǜ���XVq2�.Y{rR��W�d���LVr��h^�x-dJI�4��g��=8)�
��2+rӜߝN�9=*y��J㈸mlL�?�����r����7����=~��p����9Ө��3����Q� �fR���ej+\Hp�O9��QF�U������7��J�?-�]�{���
R��?�a�5�;�M���+%������'[�˾�\��C���@��.��cQ�aX��?�f?�Xب���Ú�T��L!uSh�_�2vD*^�"�}�/*�����b%D������z�S��Z��f<VQ���X�kc�~��U �lN�q���*�͋UT����1VZH��QF�R�|2��l�#��Ϊ�.�`cq��q�4�3ړr����q셾Qz�m:+��ˡ?̫ ��km���8H�	 ��t>�v�|Ƴ3�:[�ҩG���8��H�ԣ%��e�uk��]l�� Nt��#�G��06!~_m���'g�/:-��$�� �츌��#3�����q2o�d��8�3�A-eCf�OX=�6S�5���L�Q` �ؗ����4ߘe����/u�+8M��[���"qo%T}F�Y�;�� ��.}eY[f���b�"zr����ů�\����t�� Zs��X��7X`
����;��C���(/1�v���Lr���b��RR�o��_���L[��+���m���3�kq�\1B��͠����Ƚ��L:���|cQú7���]��z�����O��W�R��y����Pk�2�����s���YA�`t��}G��?����}�����41��e?֧��r��L"�����LRXӏP!�N�p���B_�#Ŋ~ח�s�V8<��]��7�����1��-�zێ�*���Ab|�E��r�M���������L���O@�������(��a�=m?�] �öS�Õ��;��>U�wd:��E[ͦ��;�H3����=��J/�#_�����˾����8���i�(�ml�8�lmqqǌ�|���?��ۭT����T.;-r��_��G[;��G��0����[Ç�%�´����i�h��w_�F#�h��}�+��(Gʩ���}f�����կz!h�c�x+Fi��#c�ظ���s�,0kӡ�����9�+<0J�Y�:Jz�G=߼;�&G��[����l�C��|��~��+�!�X�N�%(E�C�7���lѣH�<"�j�:ƀ�FS��(��sG���Y�/Ų#��'8Rx�W�R��׌�:��Wc�������KZ�T_�"�4V$��zlF^ӢV�H���u�Fp�h����ek;H�$� %4������ҟ����}}��'l&���n-��-���.j������q$H�������;�-�C�/["�n�f?ix� ����Z����d�-JA�.V6\�4�tc�Y��bNaݤ	��լLژ�8ww_��X�5�c���3ۢ���׊y�;QK�AA̜�oc:����=p�6׸b�+4��m�<3ܣ��`ي�嶺ΥN�Y�1�(�wS�R>�%�¸16������S��y�Jcz~��s=X� ֻU��GN�*N��-�
���+�� �#���{�m��-��)���wj�Z�_4Q�@�E)�s���+ ���n�J�vs^&ɛ�*�nm�����Y'� �95�K�7�g�A�����-磱U-�c=y��9�$��M.͎��p�B�ss���\����w�r�{�cM���Cp�Wa�F�<�.$��,��C`���'��Az �w��ޱ�׋j2	]��]S�3K�&բSN�K��'��2���ʹ\��b��d�'��/�Sy�,7������tZߡ?KAL�#%u(J|����ף�0.���z ��.�u��u�t�̘l��1lh�@RIY6�h3���D!��F75u��f[�nb�ۂߋt��^>nWw��#�:ĳ���ly��d^�\���TNL�#0d��C�}헂��.�k^�ni.R���릥5��5E���:.��2��Sn�4��~��H0����h��>�H�1��Og0XP�:>��a+.��$�s��C��#*�2$J�)/e�Q��X
� #���p���Y>��z�sN���C����`<��m.���\0*hT<1i�o�˫������hw��|���Hkw� �!Z�t_RI���SA�Ic)��
�֣奣E�C��� p�Z��Y��q:
[gK?p(/��k=�T�TB���)�����?��50�K��j�6uh�߱�:W�:�(�G���D�_���4�ۅO��.D�Gv8�lF4v��������^������Zb/.�xض1f��� ������,��,}�]����R;�!�b<I��ߋ��3�HV/��׷��m��3�$�E���|m�	�w�8�i�]|*CF� ���ߍ��_bHI�&XF�ժ�����W;����jV�W��Z�=��tz��y�)!��A~Q�����Ǡ�w�À�}RtF��y9�A�8j������*���;���G>v��v��l�*f�p+�%q���Q��[�fM��O����(��5�fI*-�Wm,�+���q?EFY���|�Q��{�̴
�۠*��4��c�6ğ�������.��Y����T|2B�(P�f![q���0�+�`��k��i�qb�l̛2l6�;�˰�b�ņ���ω"W�ZI���d��ڣ��?�UP�K��X�oJhh������I�� �8�������$����1U�d��}I�����S�w+fv��ŷ�|�q�~�M;f�6��6�l3�6ˎ����_'SpK���'G�n���]�A�>U,�f�*���&�";/�b�ǅ�;�);il�L�����kj����|5\�._�l���_/�K������N�V�I%9�rt����3��/aƄ�aD�:��)4��o�4C�Ь88dJ_FOҠ峞��V�O=�~ʍ���:���(҉b���k925�[<��+�O~h=���G
�}H�P�"���㓀Y���'���}�P+�Iy_u�O��R=��
�YΧ���/�{�I�x���Y��,�'�R����о0M�v�\�/��Ąo�;}󨹴~�^묙i�+ףۈiƿ�O�F��S��O�[����]@W?Js���v�ǥ���Қ��J�R^XM��~)j�Q��RX�}���z$�E��J��)�e:�\��� M}�W��۾�Qa^Ra�
���>�0�m�C�̍#��b��M�>���ű��%(^Q�g�G��1s���P9<���Ηs���jT�}�r��2�s�e��j�Fjp��w����_@��گ�%�U"�����;�
�)X{�T���;�!Κv�z�Ȧ~8&�Z���况�rn�h�E�W"�c͞E��krM�:�����R���-�z��d����;�-�|���v=:��L{4����r���N���k������?�׸�l:���CEAP	=��U&Tp>�s1������`�������՜��.��T�\��w�׻r�~�4�K�O4��d��ϰ{�b�ȵ��������0�v?diuѷ��a%���8ϙ�K|0�^��:b��>,!��"�N���̹���'�i���#�!>叨CE&���wFg� �j|�A�o�%�7B�_���ecZ�d�t���_7QP�=�*���s�zF&�j�Z�u[�juY�'S�!�/��K�\ڔB*���}�GOV�k�Bs
9m����H�* f�z�_=Ň#�,⋬P�}��_�*����������������V��a`�.p1H���~�O�_ן���[��.�Y������W�[����i�(5r �WГ\��O��? 4�ͅNenTp^���{�Jݲ2v )�Î��,��o��CH��#K��<�_P�
ξ��A*)RJ9���	<7��*݆14�-v*ߜh3g��\&��e5��1w^�Z�������p���y�z����/��c�"v��z:8��!���&�k0*�������%��|(�X�4F�Ә�e��9-����ic4> ���cm��!� ��Ź���?5mFg[�)��op�"t�D�=V� [t�|\��F�U�`ٹFXv�����m�c1|��[s�!m-	V~��~�����'�$����}OsX��%X�?_g�֫��dJnϼ�N՘�&IU�������rj�۲!.����D�$%�j�-u�*�ݿ�K!��F8�.Pk#���:���Ҙ�%��&(i@/�����"�#M�^������,�GGAk��km�g��g�y(��ˠ΂���X]f�;0�:���΅����>�Ŏc_�B��Z��%��[^�b}����ѣ�Њ�5O�&l�Y?���b�zh����ʂ��p��ל�SD�թٲ��/)�Y���ե4����(�����7����6�'��/Q ��Fgb4|㝞��N�h�Q�9Oj�2��iOp�b@���#��Kr)���FUH�Ć^��>Ӎ����u)�o��p�o� �
6��SPmW9�]��f�
Ź7�ԟ�������N_+�op���Y�C;hJp���?q�U$Ī�u��a5�n=R+ѣy��J��z-0W�w0�sGw7�W���D�U���J�}iNu�����d0�8�"�h�z��4� iRy�򖁎�{2���S��_��(j��/UFp�7�v���;�e4B��Y�;���/����"B'o����͗����$���D{�z��Z�-�rC�t� �}5�,�g�-�k� �3�.�E]�C8[������ø��?7��;F�o��2��R?e�����s������%7B�`���$�M�V�5� NJ�Rs���./��[�J&��*��MQ0;�7V����{�q����S7�OFX?���W��F=*�E�!� �C
�IsJ�b��!wZ[�&(%V$pH������S�������,:�-1|/K�ߗЃ����/����6������!{:�A�#�4)X=�	k?�c<(i�B!C���S)�>652��ġ���� ����	�G�qD��פ${���GQ�1�{���b8?¼ЎkhS/`�qě�M�I�>bwU;�ʏ�i6�d�awR7��_/�l��%��N=bR� |��S�$[��%���wLʯp�����L��A\ ӼA�5�}V�4�gl:�d�M�N�/�ђ#?	�{9��Fo�`�]�Q�����q������
9Z��������I������P���_x<�Z�i&o����\���Dr�p*���Vld�8�0�3�m聚ѭG ���8�㟗�O<?)���2P�����s΀��d� ��Xxn�譈D��<�ƣ�����@J��&N��L�}�k�:Ƹ`'Xk����3���\�m$�ə���:�{�Z������o�YU�=G����6�zY{��~�C&�Q�X�����{ �Eۨ.h��ʵ�u D��$���4�e3pC�9��Ty��z$�;GO�'6{5VXHy���k
FF
�@��/��B���r̋su揤�k���)�'e��կ��Z��c��ȁ�n^�6MŦB�De���&q+l�R}��ӓ�Wp���Y�k���
g�5!�<���{�#x2n���W;�˜�?����}S�����Ӻo:q�m �d�Op�u[��n��5}�%�bo$�n�������d#�Ae���:�(�X�s�W;�˜(�bJt�DO��k�P���yl⇩z8��y���-����/�:}���W4�gGZ�NC��oY������H�iMj���x}���c��������2�<5n=U�G2�7�-y���@����
�bx�y�����2��a�
�~A�?��^�6���;�T	��(�Z']��������
Zeg�";Z�^&Q	m�Hv��OMd���|��@C�_@�> ����,���儛��f�ˀG�K_a%��^�5�L5"��(h��L-�7"�����#i�	��4�dTr����!�����)��DTe��C��d3=��sp��\�2G����s7�4��������T9	�Kᡳ��,��Ť�~d;t��e����� #�
�Iƶp���x�\����ɕ3��4��8/�[$V�^i^UnL�2���$�՗+�5���_�T�"�L�D&��%����F��f����bR�?mY8�z�ްd��\�����#J�ܾ�Q�}j���!�R��;X����­g��]|�`-i�f�-��c�Bw��ͬd�����{ʂ�;���V�$]#�S��>�w�T�~/���XЖ;3O�8�)w\��м�R`*9Q���)�<�=��n0@�JY~fYAI�>��=�\̈��
f��Z֞�����kU@�g�$*�;%�+��}|�<4�>��]�C�o�rKy�9f�_�y�(����Ӊ",�d�r�2�qKy�m4��=�?	Y��.ӷB�m\2>�G��ڍ�R}���_>t�x���a�N6T��u�ɑ
{�eI�!'x��A�_fVf�۝d=5�P�d��(+59ƪ,`������J�,��Ŏ��\�Y&	��Ļ������X�7W�?�;e�۬�[|Qӈ)�9�'�++ �ꌕq�>�:Ϙ�H��>�)�� ?�E
fR�Ĥ&فK�5��CL
�}��e��[
�r�:�NN:*��/\�Xu��>	��@e�VJ<+�k\W����%��}ȵ� �P��7�?��`�ϝ���������z���Ch2�s�?Gm�`�Z�9�R�zүE��"�z7)�b}���6gf�@S��y��\tb�[�d��z���R,#�L^\67�5�bc̉�xk��3�-+Ĭ��W�l8��8�Y[j6@/�k\W`܎0��9�8���d^�,١/�r�mStK(���;u��aqA\���Gq8a)g�
�٘yt
}�R[�GO%��o��泎39�I��{���F�a���C����K\�����X�'�n}U;d#Z#]�ʽ�ꑗ���l�:x��<G-	͎톋��جp�f���"=�?b�*�\����hΫrX�PG��π����h+GUW�Յ�խ������%�R�9s��YE�#�D{iWY����n��U�
��ܾ���f���y<G�W���k�����&KBq���jx���*e��Ux�#�/��� Kh��	�_�ef�y]rib�w��덭h�\/��X��h��Z�5��Ns=20�5o��aq�S�W�����D�/M&�3��i�r)4O�m�W�e��[w�5SB��!z��:B��g"��rpi.	��k�VX��-�.n?���x���!F�}���������
X�m�2wdo�@��u. �9Z�"��
k��_�N�F2ϙ�V�ߢ(bO�?Q�)+Hd��}�cGF�_ii�;��޿,'V��>��/����L"E\�j�~S��0���_h�a�L�$)�Z�MO[�O=�]�&aRQ"�"cZ�ڹ����g�����5\.
�LQ�-�qE�87|]��zb�?�����jLv���;Sa�DP��LT�m��+V���.�Q�ت�m��hm�.�ү�h���#(k�k�If�uY�Y���C���)�����g�{����~���:v��3�m.��>�L�[$����1INS�������2%#����B�
v�E�^��f$F�~�o�X+�/^��S��xD; ���9Q3� %P�k*��U�Ãns�=�kw�n�u�A�G��ƗD!���c dZ����� �&г����I��R�1�����l�0f�=�j�񁊶FC\teN�3�!�ܹ�9�C��rE�L����o��tY��1i�$��g��9*#֠�?���xS	��[��)U�(m�;xƪ�_]d�+�0e��w�PW�[|��~��#�YJV~��u���s�pb_8aXهwq*Z�qeN��C8"�F֩#/����ד��q�1g�33���+5��
�����s%���y�ƛ���6^�t4��Z㙾��Ū�����N[�R���+�F�9wn�e�}���:V�/�%ܖ��kGSO�����J��]=�;�I�1ˊ�YE�
@ /1�����#��o�W*�=��4�倩�XrP�S��Cl��9:��>6��
�}�i�n@���}�����񯱺�G�R���DQ8�!z6��`��`fp��CW9�{%ԋ�b�hy����>��Y�~T�Ǆ�1��q0����E_�.n��!<5G_�v��i��n���x4Mj�G�pyN���q9�~�P�r0�Z"�M#�Y��I��Z����tl�%���x���h�5�r&λ��u2vq�Lz��bܓT�ʯ.:�AB���*`R�0��������%Ї����t1|��`}�j�M��]`^�uq��aG��Ѯ�j�sIb��:<f.���;V�>�2gD{��h���2��;�!{��\�KN#�d��ϚR�j,�j�b$���~��i�e��젮Z6�L�t��R��`�ǐ��
�I�����A>� I5������l��,��-���mc�]ک���n��;��JOLr�?����5[�>̠Kc�NR� G׊�bs��xG��֓�������O����գA�ӓYE��B1��$an�OZa�����C��gM��5ygWLe\`;��ޏ 98����:^����D���F�D���`[/��� �*��p��'1e��07
~��4�V��w�X��D�^������'�ox�����*-�uS�A.��в�o'�0�s�ND#�����B{�~vY�T����\"
�7��{TV�
�6���B]�Y��bS��Q��������M���B��l>[�{� ��αI�I|�@O#@!/oO��˗4�{�}6!GlI���r7��u�__�����x�u\n���.��K0O�V��8�2�1����Dq�4��:�@���W�Q~c��7�v5�i_%��6�f~�Yq��K����螡��m�U��h�	��W�rH�T�ow�NZ� �w�M��c�ٱ���ݎ�\��r�::�m#z�F�"£������}�2�ۥ�vR�S{�@7��0�ODW�sq�$�}�}*��[\UD��(�(���ｊ�J_N����2^����^�4�B`C�<��K�\G�./�Ҽ��r��k�4n�%P��u
$�����)�y��v��Q���"�����R����~�n����+3]�'Y�-/����a���T09��\�˷���H���i�/�\?s0ȥa�X���#�Q����"�H��D1����T����G����{�*�F���+s9��_�����dIY_Dck_0�Y��g���ᥱ��Ω��j��4/�����u�PH+�CkH���йԸ�c/"͜�����tD��ת�L<J�#�A����F�0��'��Q�X
�G��-5�7�f�<���iM���j�h��v7��뎕�J�nc�Xi6:S9r���l�lf� �ؽ�sZ�������ia6M�q�H�mxeo�/�����.c��� e�e���J�Rg��R_�	Y�:�����vx��<���k4(��(�er�8�z��\qS���*<}�v�薚Y�GV��(0o(��}gZ2��q�V��R��hJ�c��y��s��r�)$���G2��;��g�ew�g�|����N	�6gf��z�����u�V�pC�+��rWm�,�b58�}g�S�ȥ��+��|�g?N��YL��b8���;�̍��^�P��C��q =��1��ޟ8�d�E~�!2�Ӭ-4�-�]��V�h@Z���V4��n��R����ъ�;�;8j���!1�,���$1S_1��bDuu@�=�ļ��՘��I�z��(xq��8��%j�5�ޟP�k���--���9R8�>V؏(S�Gx'�4o�]^c����F���6m��ϴW��=vs���\c,�H��
98���h(֣?R������z'_����L��r�gW�y���
�����(�냲4���V�����8�=c(&��UB,��F-^��:�g���5�ԉlI������b_����c�ezmK�C���SWN.�y�k�ֻ6�$�#����=����)��I�/_+��7�5F�+���<�
m���#�Q[�	���GpPUO�V�8�h\У��,����;�$b�p)��7��q�K�Bu'jX�G����5�<t �A�5�ظ�T�-�9\����K����U�Q�U��հ�	�x�<f��!����<��4>�1�����ov����G��Iӎ����d�W����C��G���h��=�pBQu� �2�*B�݂v<֣FZ��?�752���*���c&S#L&��!��OL"�G�=�~���՗�nb�#���C+m�F�u\_�0���RY*=�6 ��G��*¼��7r�w�mԤ�ΝL��L��n��sN� R�d�Vk���SR�,��zm|� �<�=�-�u&>�>��a(Wʞ_�ܮ� D���*�
��c}z�Ȣ��A�|� ���V�x?�����[��C1ba��` _�y��ؒN?�]R���}��^?����_q�~}v��N9�V���1d7cL�ND!i4��Ar�L���6#������.��
�yk
[�>c�;
�xp����?�談�&Z�M�C�G_z��2[H�Z��.k�dN!��a8b���7��-#٘Y-J��@�U?&�G���o_���o����1gX��4b
��=(ŭ�AL�k#9�!���'���KFPG;��V�ıB��a��%З/��Uw&��2]���Кb=7�z���C�T}Mk�-�_���av��y����s�r��`��� O���e��+�SE�XL����V\u�k���8X��8{�2��|&�2^)��l��Y~��n�)�J�R�1OQ̊��9H�e'k�~�|$@v��ޛ(0ˀ8�H;V�B:0^���>I%F(��y_Aw� ?�(��A�8k�A�.^�IB��k��Y��U��!�Z�����z�W���z@H-�M
#��3�ANI��Z��P�=B��Y�_3YI�{�6�<$񰽞�D�M�!�Ul^�g�p�)	��6��+����D�
>��M^�:��3}��`��6�q�3^�]��ZK��@߰�2؟��0?�zt����&p���(.Bϣ'g���Q�_����0�*X䫷�+�T��}o=�]^ˠQKe�%$�"���f���Q��Qz��~s0��!�-��X=��F=�����I���S�}�n��_��ɽ}I���I��ea�z,�>�.�1v�����)V���擧�8A��h�#�v&粼�
B��������O#��c,pj;A��C!����td�#��3���`�^|K?�ea1η2��w�eh6ӌ���T_߯ʕf�+U+.�ʡ_���cL���9����U\K�	����#*�?>Lr�N�����}��%x�0������5J�/`��&�o�q��Z1S�6�[�>��/�@>�g����T9˷�J��
�<4�:��K��fM�$a<��;u���k(�4g��s.��8���Y�<�xNC˛�A)�ً�$�85�Σ�V����U�{9c����Wx�淼�	�l��x��z��{�.�<)�ʧ�I�!~m��4M�P"MhW��7�ڗ��`���׿��'�|�hs
8x2�Ɣkm�%����83�Su纼۬�����}܀�64�4\�ݖ]U��AB��JO����QF����w;����z��h�r��L](iS�At<kp���V�g�����t�C�?(�R|E��sr�"�ڋA"�G��u��ܿ
Zb�����1/e�Ջ�B���C2^c�S�3�A��8��@�$�Z�z�;�k�?\2�,`��]��՞Sr$x�9?+�<W�<5��dǾn��D~�o����;V�
�fYۿ�m���LE��ȍ�Z�m��Q�3o?�+�������NS�쪔�-/�'�l0����{�{f�آ�G~�xVS�i<iT0���ˇ�C����ָ���p?f�|���"h��d��I�L�-})�����t�&m,ogȇzi�,�#�PW����oW��ك�[K%`��m���j���ѷ=fU��i�ثJ
t��Wr�@ҷ%s:t��ĉF�f?li9�(6}MFvے���B�r+��.���*��I�w���˥*^y�p4Kśěi�U�%�%&e��:UJ�9a1f��o��%��\s��l�)>�Qcb�{=��d1�]`ޒޫ�`�Kp୐�(��e��hFC�Qy8��
�'Cݱ�HS¾ɥ��8QϙQ%� G1�;�D<�̓��X�feN,w�9�m^�7Ƙ�<H���;)�~`o��q$�b�;�%�2�"0��m��������	�w�FybW�U����8ǜ+�[K㙎���?+\��~j��&$s�O���(�j\���2�Ӵ�>�4}�:�O��)�lހv7��%���М@��ᤏY�7��q�5��O}�����^�,���k�¡'q�*�B�F�9�4��>�&�b�������i��Q���G��;�5��m["[�D�X;q��,������L�N�հ��y�2g����X�.�{c���ɑ 8��3e#���ʅ2��3#1��Ҏڄo��a8�e#�k=�V�\	�M
_���Cl�N��Y��`��)@��&��A�
�����y�-M^7Y�#�[�����]�'CңU���Α>���>uޗ�8'ѻ�ɲ[Rf��v���~���ܷ�ge�s�3��]9���H(Ob�ћ�'�g���⊨9\��Ͷ�'Xbfc��pD�Ҽ�e|e����&������km���q�Y����k]Vv�	<L�`6�@=�s��괏~�:��؅�|�y%*E�b��p_�����߱�)��Ueg�c��d�g��#�Oؿ�dz�?&�� [ג�����DF�)߭�3��渱��e;H����Ε���Q��
}������1���V�؝:�M똶��'m�R��GfA	u�!b��~ǐ}��S�D��O�H�1+�)ދ�ס�YfNIe��i7�f)�)Sj���e��G'%@�����,G���Ƒ��c���43Í~#�+Jp���͋JА�fu�9˭��sE��vU��z�C��z��ʕ�>?ms���'�����S��}.�ut�S�yrj����z�4�yB����$�����@b���t�~�E�1��b������5p>%L�>�ո�=�E̜�K6���_��S���/��1�[�U���h��#�$�8/~�)��0�4ҥ�Q���y"\"�4L����v�5s!�r�8+�O��"�hđ.����~ɒ�W��.θR}�Wz�*�t�4���T�� loF=Ƽ½�O�9sh�tF&vC=�fpԜ�!y�ɔ�S�C{�l�C�b";��wg����ߩ��:���L�OW��>ӟ������m�Pʫb����l��W��I�����{��08�C�<�#^�e��j�r��A��A?[^�QF��F��}O-_�ds^#LN���YH���� ϲ'�W�N��f3��<��C�^�J���G�����R��<�S8{1��a���n=�@}�-�e1��]���qu�z"˳��+���8,����s"��MY��SZ�1R�S��]_��sb��1�6�kx9�,��#U�P�h�Ǭ��9�`�̕6޵�8�T����WD��*D�'�lZ��)Ql����u����d�؂���Y��,�u/?�ϱ�o�3����B}�<)�W�Vu�T�q�Z20���U��10 c����(�mN�+4,u��t���:�bT�*�tV8�\\E1N�m���~^�a!�?�)����螦�挸BB�;�����F_w�E^��)�]�5�D9��K^��
;ӎ!�9�3����9��o��^�Z"Y��[;��������?��n�`4�*dyn���USI"�B+w��4@F��*��JQ5���"dvn~��W�q���ΐ��h$3��8��
�sL}2/uJ4�C�r�t/�4
U�zQ��y�ͥ�@�**P�������@s�ȿ��I��{�r�5���/% A��;ȞSj�e�!fI�ݐ��&�-�{��]rq)�c�UW����F��|��o���{��TY���^"���Bc{v[0d�L�z-AN\D͑� ��9�FJ�J?R����?6q8�e����o�x N�c�W�r�;Y�x��I[A4�O�����y���э�u�d� ��i�թ�j��X�)�1����_7O&���Ƥ�[��ȅ;��ם���a.JĬ�����hU1�o\O[#9�]y��?.D8V|e�C&��5�ܭ/K������V����nl﨣6�ZB���	�����S&�S�ϊ҃���Ǜ�x�U�>^����Մ���l�=/ ��ˤ�K����v�ӻ�6�$��4AI�ldu�nЏ���.��8��c��+�6dI�ǎ&F��/�m�szM%��1���K��g�YG�����c;2�����ߑ<_�����-6yf�"w%�}�����2�G�S[I���d@�����[�b�
1�z)^%��s�[�z�ǰ����^T�5�s�G���� �X��GBK�T�-�8a!F�AO�uyyd�U�Q �Х�dЏHv����p���^+!3ޟ4�r��Q�˅�(�R%�8��ho�x�nu>�&�^{�U*���Ũ��q�JIa����ʀoqD9PaZ+�@?b8���@ߘ����I�I=Iuac�ϴ-��7�~o��KFM�l��:ѴV�>�%�h���ͬRc������J�g�)�WK�5��	]t��O-P�V�L���`�G�Γ�����T;��8���JM���@���@�F�s�|�$�N�9��5ₗ��ds�I����:��!�5{.y��S�۬�kW1�&J_�g��?Sj�)xi�|��'���[��p
iҋe]�?}Ӯ�r�����,"}̣G~�_~��`�R���%��+�wi>*��G8`:~���U�$8f +��}'�!YW �q�W���i��-
�,�Nf�W����Rs�;~��EH�D��6�y�>��~����	��\��ĽC�ϴ�9�F�kh�
܌x��X�6�N�Év�b=����y�P��yw�c�Vц�C�T@P#Rz��Pg<�}�'��V�<�pp�ܝ��$Ǩ�m؛��v�?�Qt�?;R�Dʙ7��CǒϒI~T~0��=�H��G��b��G�E��o�$%]�H�y�](�u?м`�Y��,+���&|��O��y-xg����uY/&v2�c��0s��� �?1P9m �l![��:W��1v��Y( �m,�dvn,l����R��ə<9\�lA�����Q)p�[.,�W���!?�����2����r�[�]����
�v��'+&#��F*k*D����
����Q��k�=��P_���~���e���.�r�<2$��X	U��� qA�ʈ��N���I��T#Ϋ�E��5��̷���6m�V��6òn/���LVAS���B����d3�OkT92�]��c�X�����6�����9R�3�O��������w�3+<x��0�AZG&��Y߲R�R�#��ca�c���_��� g����TB���v�B6��J,�4��ɥ���zz���!�r������㓴�"��X��Z)���r\�=
+b���ð7��~)w�?7-+������{提r��W�1�
m�Ug;��j�Et��!+M)������4�M�%���1�k��kYYQ�J�u����܃�}�� ��g�����gBB0Ύ�	ܲnzx`���w��ĺ����I{AS���ӳpt:9�p+�~�W�A�*!���'> �����ўl�nY�g�����hF̸�a"eN�z�z��};޵���,��.�X����1,E�A�0֛_b�漿W@��>�بs ��A&&w�i��рS�w��N?ѯ�+V�	4WPʋ_��ߔ��F�0Y��1�j����G�������D7��e��e�s�����W�vRj�]G�55�/ޣQ~�%���uь�ĕ�>����ho�Zzt#��'��d>�)�F�t?�#���}�^����� ��<�2Ƌ�����c�(���:���z�+EX��]��h�؄�=�������%f%��r+�ΈD�pD��4��]Ҏ�d �;�1d�^��:|��>�KJ2
�Z?���Sg��-�����Gyx�q�I.�nR]�ו�� �y���Ճp�`�٫)�j��F�G�%�j^1G4�FUJ�y�/�t�Jk�o{�Ix?�r��
��uk!�&�@\j��'�����U��M���j�����w����]v�V���w��1��?���sDҩ�B���x�8�h�"5I�4�e�|��:���~=Z�1$�>������F�t��g��}M2�kM�S�����gb�b��/�j�DT��ns(�aI�KO��q��gY����z0V��0���G�����{�.����B��y����u~�Ђ�Z�<IG����*��Xͳ��.8��6��������d���q�m\��J�<��v5�hR_�U6༶�F��|��OiKN �EЕ��6�Zn]�s%�=2�SY��am�u:�(�����]���O�4�&lj�����pd�{N��~s��c��-�����_�6�^��@��0�h�����4E���dF�8�'��^��T&`7HIr�CVwv��u�)����!�jk?40��N9>���
��oH&�{ɛ�[NM�����$�͹�e3����x��]��_/�b0��g%��{���X!����{X����8g���!�e����@F��q�M9C[?8FJ"O������߬+>e6#�b��������H�WO���Vc�����d��6�+m�޽��Vk̪�Q_GO���ξ�g?��w���'�;�Cy��� �%��7���U�O32�My�������Waj���r5d�}�jt�w�þ�6.}O]��ٗv g��ч$oA]���c<���#V��ݑ�`8I�pR��*���4d���p�Ya��`��F�&0��'Z�o�x0v�&�imL�$���CF~U���AE������NsY��ZTO����R��PHj5ֆ�dzWk��Բ����cA���ߢ}�&r��C�[1���`����~�D��w5i��yN@`�Sl�Г����8�5z�%��B`=����XC �Xn��V�!���o�2�������j��yD���-�f��\��:sv����}@���ELE�����Xz}�^|�#t��x
}�sB����(�I	��;��'� |��]���ײ=����1,��CZJ���\@'q�j�S#>R�:�� V���f�&�:��Y�1o����\��9(�6%���;/��=����Tie�c�\1l�-��/{��[)�d�[̲*�s�Y�,cgz/����`�ԁ����S؇*�������x!w��Ny���ҰHRٙ�:��\I���4#����Nv 2k��U����i�.����c_�#bu���2�`�{6r0���/9��N�҈mXO�G��נ0���O-��D�r |�ѐo6��P#��J�[?�M����?W��S�5#M ��RG#;�"۲��o���6_W�u2r�h�G����׽�1�h�Y@�Vg(Vh�5L��P:���a:wM�=��Շ�+	��l%���$<4�����?��w�&�'��*-�#������#(w ]�����DV�O�%���I�{@޶?��C�R��V���!���ܡ��yh8g�����)6�G�q��ϡg�W��)5�F}��R'����.MB�%�v���5ܭ���L�`[��bT�ke,�q�i%�Cz­Οs�)�,�V�C�8�W�� 5.�c��Pc�g�6�W4��!�9�����ᜡ�����C�>�)�G�`��66��QR�[Ə���J���*��ص��I�Q�l���1���Ӕ�tM�<&Z����ei)M�X-�7Aۀ�!?�}0��j�-��5q:�0��ny���o��N� ����C`��n[_��a,�i�5LN\���i]���J�
��?T��c����1�x���M嶂��7L+��ES��Ÿ����*̟2��c�	nl��,1����_d�0�b���|P�㶾�:��Ѿ^f���/�Ά=r�06������>��T噕������\��;OTm'�B	�1U�V�9/ר�9G�Q����j©�j��#���m��7v�'�~F��F���7!p�dn���@b�I��z�[�ؚ8c%��ԇ<ϟ"��ǒ#�~������(��f�՞hW�6��ն�6q�]��4�J��ܫX��M�!S>@��P(@�F�z$t�zwhdJR��98���u�`X�s��<���t�c6����g��9f��l�e�$�[;�����
+�Ȕ��E��Hs��ץV�ج,�;L?K�e]ɝA������S�o]�_���U���C�|:���g�kl��Q��2c�C+�՜��T�di�m[b��n��PO&4�mF[�OJ{���a�L;�\���@R�í�֬7���X,�^Up�,��ph��zsV�9��З� m�~�+-��rb�,�Dz&��m@3�5p��߲;�5�,K�n�nr����p��fә���J�R��~����8$�r��dqh��5��mn���H�∲��Gb��-Oӟd�v��Y�>����e�N/�07jH/<q/#V�
.6eF��g���nn��������P3���<k@�S~�����G���nO��|ڐ��L][yz��a���[�9�.�0����-w�zLJ�d���;v��4�s��G�(�9�A>v1�	�{�7A� ۍ�2��ψ��/�G��Pr�ꘌR��Q��Kە�i���z���P��SC�rJ_2~XXomL|^�m�~a�(h��>닷��֘���h��H�Pf-ߺ��D�$7��Y_h�գ�Y<'^y �c[��`�����`�=����WHν�VH&
sB��`Z<SJ�PZ�E�~.�nM�]w%�V�ݞab���aj�g�L9TYS�3��Ce�򣛈Pn(6�(5�4�!]�j_�o7�y�Z�XUhl
o�2���rU�V3�M�]����d�� ��*���q{���.�K��aL|�Ȳ��{�1�)�Ĩ� �i��6>�Q\83@s*��
��U4i,�o�Sթ0��j�S~���p,rG[cW�.�!s���]��KI�&�U(���^N����I��Q�e9�P�"+vu����1Oȅ\b�-�iVq��|��SoKW��')�D���0�ʷ�;����X��S�v����HЊ5L��Li&��F�'���
ِ!���
�T��ul�,�3�`�/6t��+��1�Ge�e��ε�"]�C4���0h*LfC�}Qr��(Q_m+o�ս��ᤃ��Z�_gIP(� rK{㍙�<�{���Ze.r�'&���g[r¿���$IL=s9�@�A�(ߍ�<�[���)y�hl]�e^�V&9��vH�n��"��%q,F3�6��Q�G-~�c�t6,;UM1o�2�pM���"�
��b{:����߸օ8ٳƌ���1]n}M��Nβ,�w
Ҟ=\	W=�'�Z6D_��tH���a�,)wÐ��R�t���bT�l�4slƸ!�.!7Ll�Ԯ�W�����ΎO�B��,O�:�zc��~�"V?�`�F����n�Q��i>�t/¡��C��t۾�kF��lbs�k��R	�wb��O~Ǻz[��u���ȡ�I_���}
o.��r��}�k����Zd��У?�E��t�[5�Iv�F~�;��;�񟭽��YO���5�oMtw�=��BwGZ�w��M����J6g�-n���:NZ+���Z�O�[���a���+�lU{x��
:K4-��t�Xa�ִɤ,?0��bw߻�/�fx�~{$���tY)\2-`��e�­��:�����2���%\�����x�!{��V}��0m 6�"�x�i�����Վ�& �`ݙVk�F��������=6r
��|���߈#��D1DVO�=����+�	Sqe��f�ے�I�����o=v�Q�g�z��z������0�$gà}e�tY������N��i���3�)IQ*���N�
)%0�Ѳ�0O�^k����=rR�0���ח�h���XۏH=Vh}���9����TmlZΩ;+
��qyq�S�k��&��e�{��h\�2�C|�3�����iN�
-|H_|7،�H�R�:�K����Q�p�mA�(0Ŧ����BV���?�9�>cj�q����]�-٨_�1܆�'����t���џ���i�N��1)87ꂥ����٭Mq ��=#��{du�����n�as�]Z8�E-Jh|�t��z���_��AP��a�b�beY��k2���T�[4��Ts:�~p*��HNG N=��E��~;��$��w��|�ꂸW��!bVg)zf�-��Dv�j�Bc���ko�D�5�'MJ�� A��%j�"U�kc��~Q�j��R���҅Be��w]_w���uW�uW-P?H[h��@Y��
�:!�E�M[J��{'M���<t23w�ǹ�{ι��f�E�ϱxZt���j0�4`�6�Z�����]a�A]i�Q���\�E䳿�l6u�#+B��7'ٱ���aW/?r )ʴ+���~G3��ϟ2d���q1�S�oꍱͱ��&��Neܮ���<�'����o؊)�D_�	z���&�V�XB5��)��V�?����Ԥ��}����M�i�%/|:�rӀ�<L���|�=�π�(��m(� �$�FB��5�ÕVw�ɫ����0:�w�}��~^�7����ͽ'`'΋�Muď�o�<{����'OT�26f۽�U�ha���#Uss�B��� ����Ķ��p���[gxh~:��,
A��J��t�	�J�\/��u��d!3y�J#���en�����,��Gxk�������I(�~��G��A3հ��	=�C{���ׯ��P݀��L�����}"����+G���m4�25v������]N9�bL7���H��H\��4rۣ�yJ��`C�G{{�.̚ƋF��>��>ʼ�t�U:!��:h؋�+sa��;W׼�[�=|T��HL�t]ūU�$a�4j�U������'��,�C�X���x��w�����F��d����e����ʩ����(��r��OhptM�Z�Vt�����*��1���N��:	�˫�0�[�T���2\�*5et��|r�Zۏ�f5�(g��k!Aa����Z���� ���;/x��(� B\��B����%�ަcSZ�j�j����K�@Q�������3�OO�m
#�e�f�u���߉���lR����y:���ߣ����-�nM���@��� ��c�����z[XVՓ1���T��Z4"�"�N�s�pO�J�l�j5	���]x#��������݅J�a|�����M�0D�x<a�vD�Ї������٨��1�
��TW�P-1j��S�c�hQ�,�^�8�$4�4+���DV^���2mk&qJ�VD�CX��ӳ2g�/�����4].%��O�Z!�	[��k~R~F���W���Hė�K�P/P�3V��4�5_�KU��)P�����
����D�l5h������P�����dʈD���tQUe��Kw�'�%��h+�v�	��*�Sra�U1�e^���68�h�P:�uI��I�(�2�t�����he��C�*C5a�X�]:��ް4��=�;�j?��<��w�[L����BCR��E�8�
\cZ�M��#�����Q~qԫ+��ϟơ�J��������>^uye.���x��^����
�1��H#�p�j���$Ev�y=ϻ}�`S��������������`;�`B�+�	ѶQ��<����X"<��<ͳP�bZ��$�O%ŕ��N	�P�y�I�ǌ%�V�s��ɅAgK���]�z�m�ҟJ��0���3o�!��SΧ&���S���Ô�3v�n)�~͌�>���!)�U���Z@	,|p��@�iK�
����A�@��k������v��dxIB�%���&�r@I�g(���V\1�"D%\��f4���VN{���~C+�����.a�^r�{�����kLT	A�2�4/M�>�|���\^�1�� � |�M�=�����H�f���s�ټ�A���6r��>	����s��@[I��)>�T��aKR�wI{�"��^�`�~/�5Fzb���6��Xݠ�������a�QS�+a�t��:��� z 6<�5h}J��G�q+?�%&��M$n��8�-� �P�6�+X9������͢�S�r�����!�C��8�� vx,��	]Q�M`Y����xʉ?*ǡ��g�'T��y��!{�t]�fo8��|�(��t�!�F��_��JGز?��X��j1�P2���<���~��i��[��sװ���Qۓ�Rf��S<'��r�I^l�P*pre�\�ʕ��aכ3��dM�LT�S!� �c܈^YjWU�7�Vː ��C���t�SY2t�������e�+�ŌBg���?�3jį,�C#5H?1`TN��JV��'H�/��,�F��8���0��Ufn���B��zI�u��1�Tq�JH�b����'`k�w���|�7��c����6�}~̌���G��<a��F�c�7�)�2�� *`q��V�!��Pmgn˳�@���P�KlH�l�Zt���G���I��C�SF��?S	��F�=@x��+%|T0N!�
}]BQ�1h{�S���5�HTPD�g#~�'��<���#Kγ�G�� �om�4y6��q}��g���z|�̅e1U����0g ��b,v#,嫈M�
�uYNV V"s�G��i����B>Z�W┚ƲU~�KA%HC]�����_�SV$������H�}O�O�d"��������-�I��N�=D�����
����H�,4����\�[:L�!%���T�TB�8�]E�����ـu��`㎣}7b	��>n[�;�̾���9��;_Ȁ8��E0��8Q�~�Q�Ah-�X��C�+���"�	�A<^��y�t�2��`��2��P-��<�<�Hz#��������ׅ#�&�+���+h_t��}�H&i�Y�3HӍA1<h�
�wv �����.��'�!=�O��q�8�+o�_$=C+�&�Q��%�G%�xx�R���ը��Ja�X`��V{D�3<�� ch�c�W�E��+ ��G-�B[2��;(ˁʙ��y���Q:4���'����"�&��f����G���NM�H��|��Fa!B��ڢ�e !�ݾ��I�i!���&E�"o �Ք(�A1
؈��F��,���j�o����]dK��*o�>�!{K7 �3Od3��a�Q~��"�nEM��m��1��[,|�y������-�K�i����((3&�E���YH�uAg��tfT@���ު<6.������p���Ў`=�C��9M\??�{i��ʊB#9�D��*�W����@�q��7�X��ޥ���"G:��rKw�*\�n4�r��Vօ��;�����g�F7�VJb�Ȗ�a���,,P�tb,*T��l#�6e�h���� ��܆�~���c�ľ��mP��}dx�!��i�{gY�<5U.����f�
�y,a��_�G��cF,VO��,�!e�nU^�&��A[?�
�'w?ؘ?Ƶp���9aݻ�������RgU��5�Ø�Ff!����Q�
�	�T�����^��3�k��1��r��4�|���%��ð�f].���\����B�*�-�Pf�"~}»@���꫏��F5N���I�����<�FM�|T��|�S�|u�W�&x�HE�ܥ+go��&=X�r�gHA<%h�#je�*\'�V��!��?1��0>�_�%��e�\��f�,�~��0;8:uB��]������B:�0w3������/<�=C�@��)=���R����]	5�zv�H���e,n1�,��a�Tc�r�W���!�ab�H��T�උR�?\�>oP�	����(���"/Өd;w�I}ྼ�c(�~�@��M�R������Ro��R��w�����\��<5rO}m(h��__���E���H�kp<):����S뮊!��0kG��x}
x��Y�I3�Sy�J��2�4r�����n��O�/��>:KR���Y�v#�b<޳CX���S�="����k��͠
Wvv�/Xe��=��/4(���88���w�S�0�S�4��w���l�Fh��+$���dj����/tIM�?�d����/+L�%�0Ui:���@�^'e��Nz�ć���֕�	'�X�v:9��t�r���3���<*Te,��2ώ�m��ot�m����{�e�~�,�:���T�d�d^�%t��#�?���@��P��y.!Y9/����D�_���.�v�TȔ�矯�)wwD�2]������VgL9�"TO$9�M���b�?a���t6�_P�mF�����,��x������p��6�.�WR��^�+'a�ʭ��s�@ܠ�b/i�
�Mi��-l�e�U�d��g��N1�����N#��}񮣑���n$巖XU�Է���0@��q���o��\q��U.%_|�"��M���JbO���m��0�����c�a��<Of�}9�i�Q��l��#]L�@�C-�A�������� x��.�>B����'�I'�l`����������(~�O��lf�x��P���0��4�`�;_��8ɛ�/+Qx���=��>n���Wys��	�#�S�U�$.S8ʸ�&)?mU<��K�3~�����k��^~v���e���8�ł�4Q�& �[_�?"p�v17-u=�M.&�,�D�(�6�`=���O�Dbn~�?�v����xs2�%wq�
6䛉v�H{�v�.0�>m%)~��֫t�N-�ɶ���+���糼������䞆1٢�ۧgQ����Y��TRg�����D7HOǗ%[r��J/�Lx�8�	/!�����k������FUԎOyev�<�x�/��Πs����ҁ���w�8X�Z��:��D6�Z���quȹo�Y�'1�E��D���<Ux��3���zͫ���La��T<@ߦ��R<.���X:$������qd����!|26��&g��0u�8�p�R�#��^u~N^ձ����<6�i ��Gn���#(�����y�ң>�[�w����.鏅�}I������o���XH��s��F3Ӣ��,"0������X�ꋌ���P�AⅭE1�M�^1��0�˹��of82~L���Bun/YQ퓌B�3�jێ\��
�L�\��)SmD�3buP��I��(a�zL�c�#�Y�Zj&����&'oO/`�o�����A2�\D�
1��Ѱ[�yحҗz��Yc�R1ot/�H�33�۟L��b�Ie��v�	g�
hK�2,��l�u���/�V����/�h�㚞��_11�m���1b�5�i�2b�O�6���$��$�Q�ȇ�n�Z��N�y������Y�N���S�b(�����������K-+W�S��%ڪ��qu�h�y��b�hyP;�
.�ώ��~xK<u�I1�ú�U�>]��R\��ä��#�(`nK/�����̉'�5DN����f����C����ָ(Wf�e����L��a����*�c�8���ơ���(���<��+}���,8?�^TR������Ĭt��my�7g�����-^�����z˦��lR���T�(��c$vf~�`����EI]��_���g�ڦ��i��λQ��A��	���M�#�r��8���SA�Ђ���U�˫4�}���ٕ�.^��&]��Y�����u���
d�~&�s?ѓ�J[eL�i��+�VJk�*���2o�YC��+?�c��t
�yE���Иݷ�RE!��z�9Щ��3o�L�����,�_pH��n#Y�1I�C�$Ɗ��ɫ�[��=��FY�͹��q:(�	Ro �i0��"�yr °ؙ<+.��NO�7���2�8�LR�Fv`��ĻO�@p-�~�P�z<r\S����o��k�-�y��G_0���������ZW\X�	ҋ�D6�c;��NI�C���"*9"\��,E6'��UV
1|�����:
��������Qt~�ld�5�ɚ��;�����n4*~�����mE|*׳mZT����v�C
�_�5Q��!)@p7����Ǚ�\��������z�nQq���$�Jx�`e�H�	��!T��1�#F�dO�-?���O+��F`�d~ �6���Ye	M��^��e��G��Ҡ��YB���/�-~]��ujL��3�c�dG��3���&�4y���ر����L��˷Ve ��歺1N �<�x����i���I������;��^�@ (N_ 6&��Ə�0�K�ʓ�ws+��,"�\b�c���Ǭ���������, �!�ky�q1Ehb�.RY'lڨ����ę��O�?�Ie��q���0#���F�#��:���7�,x�YI������N�Z2���������peD�-��[y+�R�7cPU���K4㾁���i�A�0Xv��/uv�I	��4�	�L�O��P,M��\�q>|H8�����ky�<D,��^\,*��80w�:2Υx�3W�
̃�`&� �~��K��l�X�?`�=��:��H��<m+o�}̰��h�8*�S`�J*���gi �%Ń�w�y�T"�b�a���nr�=*Zb�}�s�'/��9 >N�P2��ҿ���'���AO�@�J�>!�d.>��@B�F�U�S��=�S�^�-NsA�9SI���[��ޛ�d���D�A�>�#�L6.�QLTb�8bq����z�[6,�ĥujV���D�f$�r�6��� SĊ)k��g���0��(�[2܀�"�\�V-zV��	ܣ����7U�8��3�B�R��Ml�_$��"§�]�E�"�YL���̖3�v�j�����N�(�x�B�-o�*�P��X�'�����;�n�h�<�=�k60��\�n�a��|����?��[u䤍��8�~�#�ҹA�\:�/l٫�~>�,�RXjeHcNK}3:�_iw�ۈC ��G�B�Ɉ�'n�Od�ݸ�5l�@"�n�-P֎��F�	.�Ӹ�G��waB�\�Y�gjNt���w��^����/D���4����Ei}�[��.>#Z�F����?��1�D$��9�hU]r������Dc�35�\Ȳ)�]��VWl��d�`�4���p����}�jf���%�xs��G^�>N����ەU&דcv��n֜��/$�l�v�u�><�L�{���*x�u�>J�vw߄Mh?��5<�����'?�ri�fo�!�W,�`���אX�������(��
�s��>ݪ'�'�}�U�{"�tw_�ʑ�(I��,�X��k��R0���X�8�Y�P�H�G�V0�b�(E������M�3����Ԅ�0P�y6��~C�r�vG��Z(�[:8v�)?��`����H�n�!�]jؖ��r��;���?c���	OZt�4�b�P�������_ەc�+ߖ$��/60�G�O"w�Ś#z�z�f���D>P���!T߅3������"ZʗxdM�A�A��㱶p�'�Xh�P���Hc���c�Y[lb����8�[,,����1u�y%�EhG��!Qe�t���/�lC��$���ϭ	�]����ʪJ[�FT#�#�b�^��J�#�����z�"�M�Q$��e�c˂@V�U��3�72[�_�����s��2
�1��/�]��"�,�{��!��	63ssSL�s�x� �o�C�?�c6�mA��⏓�:�Ɠ�'㔫k�#�q�a2���;�&�ʨy@��xx�VRV[@D��Ln&�(p�@�L����E�z�DcU�-�K�����,Z�uF�Iơt:e��h����^!�XXߌlAm��L[�{�x%}���4�ueM�:-��`��6��Dkr|!����^�n���gY�v.g��+/A��;��j�}G���=�z#v̱j�x��˥>i�>����z��S���z��8)% �6��;t���_�A{�簴,�QcF��4�Ǥ�F�w�"�t!��d���n�	.����u��Tՙd?��/f���9��4���Ã�l�0�aȗQ�}���%�V��i���R��n�V�d�����	��@�~�ώ�����1S�VHJ��zh�%3ȫg��mFyL9��3L���W�O�eG����]�u�gWEm#�΁��0������߳�����������W
Z+��Q�O�Ab�#�^V�}�޿A+U��S#-=00�Jl$���LJY�����&��}:�}����$�D���|d�.��42���!�@I�*��}Y3H#5�_I�VC;�������c�3�f�"���L'^���ֳ�6�QFi�6��G1����0.HB�hv��3o�Ug41�uO\K�)0�H9?�ˋ	�:Ј�����TD�'�ձ8w�vtd5&����:�GM<�R��2n����;��ݤ�>1���蓫�]������@9�Ȑ�RZ�<gb6?�҅�s��8���"�J�� ����ZE�b�r%E-*�ܿ��+����j�B����Pu���&q\x�f��%t1�2�Y_��~�٣����u2�&��L��^Kd%X��_ )��v��ruɵP�k�c����!ύ2��G�|�~6d2�P{}?��m����ª�Gd�Yd�(TT-��y�,_9W}?0p~���.��G��5�9݋��'�1dH�z�� D��l�2Bb�3ָ��9��-�N�P�P��40W�~NG{�]GR� .�c&�8�d�e�:� s�7�.z�_[[�4I/=e�Uw���b����f	�R?��*(mP�n�D]M�NƻG���'KW�dTN�v��K�P�M�@qiZ�4�	@����^�Q�vsO$X����WF11�D9m���,�:����Q%P�ca�J�<��N�W�-��wuߖ,_�}�t%A�d���>r�,#[�h~�[�P�w�A*."J{��������!S�Ux�Ѫ!62�'&d�dL��=JP�,$�*��������_ݪ�߅!d.,�rJ�uS"�*#��2n��O��o�IA�
O�w�a~��Z�<7��Md�bbQ+FYy�%^3~"�+.u|&e�[��%ºC�ؓ�Z����(gѾ�TA��B{�g6�b�2d��S������%o_�P7�Q��~ ~���Q]��6M����V]�GW ���ff\Y	�,��ژ�-��4�#�W3Ɍ4G�{v��X^�J-9��"��d$�d�4�I�9w-��R����.?����W �o���@�A�r�P���+������n���U����C�%Tc�*��t7
���/ܾ�0 0���=L-��]�I��==ef,�6�i4��Ϋ������py�|<���v2��Cǟ�S�M�1�u�q��\,Y�9s�R�E�+�P]5�N.��GB��izi꼘���g�Q\ o�1����>��r�ѩ+`Z�Pc��2��4�^13�)7Hǭ��>��G��Oc4��0���mr���'�x�n�: N��#f�z �����nd��-ʲY���N	�M]�~+�g� ~d�=xM1��r�^�Ʀ]������b���wH3`�E��l�������8/����Y�t�R���t��q�ag ���A�U�R3���f���������{���?2� �yQ�sQ����c�\.���6���P�_f݆�C�_z�>b�TC��ޭX��CD����mH�*�V�=��R�� �t��"?�+eJ���W��s����=�G��������{e�F��)��������h�(soF�T,0���L^j���>���|3ݖ�|[�J+���0�i�J�'�ό�0})t:L��Q5��Yh3	Ϛ��!���'��^�!�|�6�=�Fas�o~sX���W�J!�sgj�u�е����O�=�������įIKa�8�_�~3SS��倏��G+��|=p#H\�R[v��:�c؃�`&K#is��W�k2��y��6����6�~vZ�s9�6a��,3��}]�&�𒏺t�"=ѫON����4��Z�Ã��A��v_��L;K$��[0��7L|5��l�b�ق��1�Z6%7��Z;�����|U�����-�˯�� �J�f�b�ڞ"���j�Hh3Cj��cن����������u�۞lk��ځ:��>lo^ir�;�ho?���GKA8:a�U��5FJ�U�Zq��W���V�C�(눵 �js�K>�ads�܍F�#+w�V��=p|��u{�ߨ}���!���C����j���e)S1�ײB�]�܍&l��\J��^�I�\�+�6����.�9C�sB��($K�t^51���-L��c�J��|,��>� l�/��Ky�ȑ=S�ص�J��	)��P-���"���u�i�p��*��0��gG��J��A�4ց�*_Ee�Q%�_��GH���7��`��4�c� a��&ş�c�TU ��@��C���m��X����{:����3N�הs������)�/g�u�[ʙ�����7m��M/�u�W�*n�H׊M[�Z������\{N���ϡC��S-E�}�Q�:��逸5�w��ފ����vG�}���`�S���wD��o�D��h�E0��T��_�\�/W���:�nh9��r����������Z1	��M>�8�{:�1L� !Q�ŭ���L.b`��	0�5�-�*���]��&���|�5����3��|���m���4J�_z����wh5��Wȝh��7���a}R�Q��$�nG81G�Vu�;G�#�����;JF�B�ǀnF��aL*e�QbbJ�,�Ei2�-;�-���;���}=Q��MXQ��Q�1���)?��s���g��R�@TF)��W}ʂ���>�ܭS�����m"�Z侇��V��j�<�;���ý=�$;���:��V��Vy�^�#�d#���s%�EF���{�߉EPqBq�T2] 5_649:�q����,Z�&�w���(xP�F9<]�dB54o�aXp�ۄ�xS�xܙR/|3	�a9�7Y���$��P�O���������#Ak���U\�w
�q,�g���{�;���6k��/�{����^.�\1{�l�ä��7�"��n����L/�S3TM:��u��l.���Zew{7zK�M/����ADу�) �q�~1��j@Y����o�Hd��=�=$�<�Δ�y��pָ��
|�®��6!��^����yZ!�=)��X��0_�v;�Sݘ N�V�w���d�	#�~'�^��仏/P�=,D.����(�@�ч�ï�i��k0�1v��uoІ�{�'�^�H�7���0���:�&�taM�/^�����47ZS%R��
�r��Z u���j���%�-ID��)�Q��#�����Z���#�t�� <�W0�=�p�'���f;:��]��/�������/>f�~`�f�����x�MŬ��Z��rc��Q��\u�Z������8�f(ړ�������X�K�%��K�)q�/QtR�j�X�P�8�%���Zѱ���wDǳ�O-5a��b)s�TQY�������హ�f?8�������p<+O�1d�d�3m�9\�Y�y�(��L���l[Ћ���v����n��K��	F�2�7Q]�N�]go'm�qw��R`���V(�i�K�A�.��h]aΫ�����a�0v9�պ>oʾ3��yO\h'���Pm�|�id��^�&���|��:�/T��?�J�h�R���(N�^���|KD���otO�S9��XD -�~F�#'��D��1S�jշ�F=�uÎXbVm64"-6 ]#�*_�{��b\����]dF���=ޅ�X���0+��A."k{�0�jޙ�84�(����OC�S��NC��Bjv�x�>a��f��-`�.Ȑ���#�3M.Nw�@Ǌ͚��%S޾���6��'��0t�'S;��3������� �v��d� ���j�6j<��?�du~�)����Q4$UN�?Ҥ
}�����X������A����a�.�ME�TsA��	�������&�N8a�1I��/��y ���կ,?T�<K�is5��������DCh��Y���xv��R�3d�ˈӫ��2��"ˬ`�xdz-�/�����@�=R����̀z���Č��|��G�T2B�v�0�7���x4�N���E�O�g�J�������Ϗ܌v2�L&Yd���[���l �y"嫕Y�OӢO���{a)�M���ݑ{���q����sH��>v6 kq����v?d�/#�L�B��a�ljWZ/g_��"�7\���8Q���6TA�W�o�u�BP���P�W��\�����}e����=��yh�{��9ٌ9�G�ѩ*鏙���ѩR��T��;���S�a�f7͝8�=� � ��8�ؙ����ﻇ���kpZ?�/0��N&֛d�5�%���x�F��������hFQ~��l�)e�W�5�+_�>��X��R�[6��0�,��O�&j(V1��W0f
F������E��h#��:�q�l@B�i��ͯ^<� 4⣡���3�c�T���>���&|o�I��D	�P���a��BM=UR�R�`D��r��w§Q߼Hݷ���-��'.~1NL���������T�BU1��,����ɵ�U���Q�8�@E6w��/���Z��o��M@�ؼ>܄E�'��P�ȣ�SO��W��*PE+_�x��L ���!�A�?8���0!�<$��X!������d�iy�7�i<6�O�Y
��a�`�l<�`u���*e1.��k��ur0x.l/�
�v����o���>�=�צO_$8л�F.�� t���'���J�Z�}�/i�N� �����g3M/�/�,;���dtF��M� 0�.`�\*Wt3����e2����R|��cІ}4/�o�o��i����a��Ey3�x-�n�Q���#M&��CL&���`��*#��XD
���]׺㱧ZZ��`��LZv݀��v��P M7J�ک�jm<�ZdT5a
�e�
N d��P�&����L�V�g��x ϔ�p?]�����Ma�S	{�1�<��ω�a�03N�ރ����ʃ�`��1�o�>lK������;�������FX���&�	��M�C��i۹��J�1��MxP�Ym�lҍt7���x��������c�){L�D�}h$�'s73o��תBH�*�<-�Q����w��3���y���L�7���z�5o�C��AS�aS��'���w&J��#��T����"~mx��B��1�9O���m4�����$���I�^����k����Λh�ׁ�(�=�_ft���N��ދ��q{Ѯ�c������ l��(��5���b�~-��O�I���OPg(Y6��d�q*��4���ߢZd��k�Nљ<4��4	U�M���n�2�ah���X$���r_��4���:�0n��MF����>���܍��0A�N#�ϡ�bLǢ�w_D�)D�����B�ihh�)�@�P��z��BqR�7G+�=X����5���%zB5q�"{�x�G��6��n�YC�vYj@������F��3ZT���*^ݽo��ł��m���Q?2b��C��F�<ĳ�����T���r[)��&,�%����j﷟��K��~�T�>��o��R7�"L�wF����>x��G�E��{�x����M!Q�����>��^l6"S�g����O��E^�t�12j>����;o���z�o�X3�^�7e��1���A��yO���+yL��l�n��*�9��
/��S�u}/>5��.рؗn��X���hmi�3�w0H�禹�c��̔��u\J>�f�u�J[%V�L�Ļq7�KÈn��Y�7a����o��d�R+N5T��`�(����s�h��$ ��}�d�
�q��hu�B���*5�����#����4��b?�q*
�כ���B�.�ڀ���K.C�o����z��Cˏ���Ꮯ��jCk��v������V3���'��C��U����f|�W�x�}���Qw��Fw��;��*������
|�Qyk��W��<��e��K�	[�����6{s�,����,O�{�юڗ��a�BG�C��_{B	�RY6e�
ĳ��l:(h��{S�	[�F�3\ⱀ�x������-3YBI���8N-���Cq�1�nCC�xz��ɀ����Mj�G�=h@�8ZF�a��&�C����3C�`����&<�o��y�k���>�N}<��@�*կ��_�e~g`���5��.oI�fW�V1�8�o��ܐ�ؽ$ho�V�}�;�Z�m�B�>�bhy��(H>g�#�`�$�P�9��9H�Ā\j����Cc�8�w�=�C6٢T���i��;U8�.1Ujj�V���Mx�B)j�Qu�Y�Kە ��9`��m�"�4��cY�jx@���{�7U�5϶;���R�2�!ޯ�ZSU�=b|U��"�w��-ƻ��l���ꝁw�\�p������G\�Ý���~�[���(GV�����iU��ˆ��H�����Q%.��Y��k  /Ӿ���/�GT&`�~7N��bL��Ri���!�LUX�g��;C�zڤ^�Ԋ��p�,�]�9���Ha�x�i��jo	�e)�*5 �%�D]����+uk����gƺ�2mz�Y`~4EX��D5���6O�k8-{4R/u�_c�!�;�>��n��Avq��nW��dC(g�>B�A
�k?�!|/���C�|'Ѵ���7�W�z,�����n�P���fs��җK�v��^rvm\����>�R6��SPU'TH8�l�Pg���H +���ϱ����e�
�S30?l^�鼍���Q�� �)�AU�#�EoL��͓tS)K��F�m��i��ko�>+5I��h*��_&��l�r�.�/|t�4 �L��]���L��ZX���8+5Ja����z��z�UE���c0V>A�g��7��'�U:u��T�$~	�%R8YÁo��q �w�.��ٍ��JM��:.#��8�cגK����Q-���{�)-<N8?�h��Ķ�l�� �v'jn�+�XWJB7����@��4�X8�. X�n�&�E�[:��,�x����ᷣ}y���.w'zU�]���s(�I��}>���j�ݭt��>�+��
����?&�)���C�ǧ��7��Pi�:}�8=��J��[��G����,<B�����`��/�0ٰ�:�z\x���!�����/����ൈ�\%X �����G��&uŝA}$F� ��"n"�!¯�C1�ؕ	���~#@
� �O����G��gǺR2+	O-�\��]̿�S:�}��x��g���<ǻ �ݡ(�}GxX!��xw ������w�� ������Ə�E��:���?}�z�����C�Y��,9��(���Z�/ѱa+ƪ3c`'�z<���V\#C�Y�٦��&���h�^^��	�{��qH�1ҹL�t�.Y�|#/�ˏ��P��C��������kT��i��n��]�k�Swߛ����p��P�7yI���&F���3^�;��!�����GSu���k�̪���b�ʘ��6�B����x�/W�D�Ϧv�_M�r=�~�?�xr���{��S#xn�`(�j*~�&x=�_smW�G������qwj��c �#i0غr���czN�8���:='��ہ��F��|��i60�=�Tý�Ė�x/CqV�_M���7*�c�f^�.�����YL����k�
���q�Pk�B����uB�R�׏Ģ�RQ�=-VA���L��#�m:!����-��Q�Zǉ.� ��1�&�����/����VӀ�����lz��ڵ3ΕϜ�B�m�����\
|�I���C+�ioŵ��t���Y{+���R�O~���v���2m,Z���5t�h	��G��曪�y���G��@����v�m���5�ީ�Q�o����>�+5 ((l�۪O��0�T[�\`�dBC�������@ �L]�A1G*e�b�> CE;�ig�V�|�RCt�&��:�=m��6A���'"؅j�V�Y_��Z��z�>:�p\L� eX���3P��l4K�j�����hK�P>�$T�'b�9t)�O�� �P C��M^ǧ@�<��(b]
�!�J�:SL��g�5�� `^ht{ �g$��� %�����ΊY�b�` x� 2vD��@|*4�D��w*#�� ���K�G�\ƾ�f��Q����r�~��iC���xC�)<��9=��/�WK�,��X��dN�P���������j��7�8V͢��_���	�u��d�#���l�l��f��O���m��j��OD?X���Bl������7\�MWc�����i%��I:�c���)��K��B�r�?����Gu�8C8d�U1������'�c�	��Bhn��I�#�U8ږI��DFy7�s�D·Rx����M�N�����e1cs�A��_��Sx�.ę���A/��~��O d�Js��-���Z Y���|=���?�"4��3�F��R����1��OǺa��UJ�͐���1�l#Q2���'�Y�n��Υ�'�\"�:f+�		
k�!J��4����J|Ri��{�{@�sm%@�Kڐ�,��@(^���1Ȩ��%�0��C%�?�<s�@{����]N5���
mS�;��~Z_���ԡ�z��=�\���1�����ﭗ#���(�O�`K��+��A<�.$�D�7>	�o���!��Kn���a�r�%D}i��j�x�Tek"VYBU^�SU�V���U�O�c�]�V2�U��D�>L �??�ބ�0	c{�b����z��������=;P�v��5�������;[�>�|�U���O�:��z��~��X0G'ez ~cG�"o���0J����;.`M��c�>����}��'�7��I��\Z�o��[h@`ϻ �s�#�>h��y�������X�i.O�c��u��!�̾oK@�a_�K�'��=9�ħ}��A����/�gl�����HN](�.�W^�����M 	�o�xx�Oãb<�'qx<E(�������a����_���>���:��_5��S��?�Pu��c(��G��J[��~-2�k�4�?܃���_���%wâ9	4�t�%i��/�t��.�3����(Ԯ����Oį%���+�	��[L{�2�ǯ��K�/_�|�F��%�Zם4
_+�4������ý����E�ǿ����a�P�j��C��4�c
)�;��uG@���f~| �CbQ�	�/�%Zs�W���G��h1ls ~�(��D�	1(�L���U8	�+��>��̩a�b�x�t���w_������jT�Q<�+�B���rm)�P?�-�Q}��H����Qo�9s5�±�_C�:�z��lJ�-w���\�$:�푎��Kƴ�)�jL)�8�Q�M�M� M;���Qqc��Q�g�w��x1-��/B�WA�=�xC�_4���z��~Q�2�oXc:[�i�1W�3\���7ݯ��º�h��o�f�Xt5큋�]�+C���v�9�p;eo;\��SMO���i_֢ʅE}�FߚmB.���3��t$ϧz�#���hr�;��M�K�FDjh=؃��ô��d<m����Sd2��wH<╘��k����ıŇ鮽u�YRꕱ�>qx�D<�n�05�ǐ��Ia��+��7��m�-��_����c���#�i����į3��<vkPAt+���u�ã~�0�n�5�G>"M�^��=�i��O��C��\&.��T�5�=��`|H�����؝���1r����mp$>�~��՗���I�T�Wץ�
�!vƭAl��J�?��P��1j�ʞU�����y��.�r��l�/��{/��������������}����\~5�_���4~_ʯV~]į�������#���_O�k.?�_K�5�_���/���[��[�������_����;�u'n�����Y�GCH�.��E�*�k�V�k%�V��:~��ח�u#�n��7��~�Ư�_w��N~��_������_O�k'��ȯa~=ǯ>^=�T��pQ�˯��j�W����ǯ���k�:����u���T�S~�˯��u1�V��Z~]ǯ�u��̯��k������*]����i�Ӥ�*��z�O�s�J�i�R�ҹ6�eG��"�B��ψǞ������O0ߗf.Y�:e�;�u��/O���䇠Q'��i�����΋����ј1�P��Q{�p��6��U,5NS�B�>�����*.��ZqR��^H�̚�8S:8C��lJM�>�G�Eo��.7]%_!La�'{������h��q�n�$/6�5�|s(S��FJi��#��0�+��$��#9��rG�1�J��(���DJt��d��srU�j��]���a	�G��/�����%�yrN�<3�ycZ��V�9�*�ߑ'[e�;� %������xZD����x
���'��`(W�['��h��"���y�M���p�H(A�)�gK{p�{3�9��.��8���W)ԔrOWŝ�DA`G��/-���۴RA��SF�-��SL�fW"����rZ�4̒¨��@5���&�6W���K{	��,Y'O��Ef�c����bC>�($�rI���><��_�k�@�"��}�H�핾�����ũ���Ł�L�f�Uy�st�-�7SZ��Ҋ�I�)�_�q^��������
�?��)eQ��31�[�7���X��u�{��J�F�T��_�=P�j̀�٦�p��YpTˢ��hfVhKUF`E[���6O�I9�rm7j$�h����{��ô����ιwk��x�"[ih�\�>fnyҽ¦G��a<f��+�-��}�t��I�V�����Lpw��\�����%��]��.SU�ͤ����U�#����;�v�����%�<˜�is��~ve�h<�w���l%�m
�c͑t��$�Ⱦ�����pZ�Q�B�[��i��l)�H��mJY�5���׸L �2��6���ݍz���V��Ľ�7S��\���|B^��V�n�j�@�{��]��Ia~���ID16B{��4ڙ�)[�k�L: OQ$�� ��7��}��Tx[�#>"k��8�}��;��
�0a���6�G�����R@�ХRC�1��ؔ9�(�;����a�*h�5��C/߮�1�&��ޅ]�F�Nʽ݈q=Y3���(o�'Y�=��ԗ�,�I���(kɏ�U��B��ʹ��H�H��Cc��z�N���4�f�TGSR���Y�{ڰ<�f�Ԡ��ӯ�7�o�y����u���H�
R�5Ѥ�U�ŧj�����|?�������q�ߺ{�
��;� V�����d��ay
W���/s�2�wM��6�0
#���h�b�Y�TM,5�n2�HL��n�.���J��W�Z=����m�1��̀`f��w��5J�f�K�ghq@�t�v�0������ ��ۄڼ�;Mʼ�q ��S�%4v����b���ײ<�2	[SK���h�n�����&l�Xjfak��M�28`A,Շn�~�(/A�G�͸���t�7F�&�ǅ�sCH�^�A�4S'\K)�6�1��FC��E��a)��*��+���������Д�5��8�h��68�Q.]w]�d�m\!0X`�%�d΀i��y����rz�:�e<4톖��ϰv����1.s��TYͿJ��0���5+fT�����E{�_�l�b�#��JC�wz]�	�����>˽0Y�F�k(��d��,�(�I9����u�����R�b�������»Z`<a��pð.M�a1K�#r�㦛��RF<[���霙Qn�Se%�g�S�􇹃�Q.&
֔k��&R)E�4�\�0�����a4����s!���	.���\0�0y4���I�FI�+m��c��&�5Y��gd6����ͷ(v�"�b��+�tj�.���:�5@��m��<�F�N�3������J�!�lv��jsc�l�@߈.x�6�F�`C�ϔ�z��r�K����P�h�B
�]O��J��{X���߅��S�
�ap!>���òA��K���ѐM'�8�Z��0���P�{�i�Z?�P�UL���M2����*��]lJ`*/�;d���l�*߫�f�w�[� �H%Z&���
J�M�J+<���87����H������V�Ao�!BHn�´�0b:wOG$̒�S�~m��N�B���uz[0bzh���c�X�œ?��5�a�E�oG}��,f��A�_�P0b�C+x<x���0Mr����+)9�Mֿ���Tu6���RI)Ϝi�-��QZ��Yw����F�LIŮ�3l��vSN& ���@C��эnf�����#pdq���鋞�5ܝ:�pr
mYu����F�#0R��1�e�~������������'[�}���Uѕ}�֕���2R#׭UO��p���E#u�#t�gA�	_,M�H�A�i�P�H��*?�2�r�MNUj�s�j��ȯ�5f7�Ș�}:Rq�\��x�<�*%?���"��wJ���f #?�4q��t��٩�l+j��XW�6��yZe��d؄8�<� �>�zܽ¨�xX�"34�C+���}�F�bO�k��s�We���C��m�z�����87A�%�T��X��j��ݫ�@��S�ⴈ�1� �|��N^�n7�75:�=�գ��zڬ���EBIj��I��9Tq�<٢��>�ҾRH��*Z�Q�.g�U|F^����]!A�"��7S���=ǩ_!�Q4�l� 19���ht�u?r�@�δ�lJy8��`��ίaH�C6����g��$.芽�cQ$ ���MԧѢl�i���I��i���1�t�]�z�{_��n��V�h��  *��q�UJ�j��������J#
j���Ϥ
/��@�  �i�7�A*����̀��R�r�u%E~ Y�24R�j�,�ݍ�3}�J�*�����8�����2,�e���]@t�a�À},�gZ``(�A����A�H�ɝx���!��W�=1���\
��b�?�����6���<��'0�ް4r��j�%@��E܏���"}��&�kT�ͫkĹHW���K&l͹9���i|&3�㴞����D�
�V���X�"��)$�	�X���EUI� �5gP��?���U|WRw�>˲�E����ܧG��X�%P��T#��P��6�L��v7X��z��NJ�hwkl岾�e��M	991�;�x�b�;LE�M��y9E�l=���i;U��)Ӄ����TOC"q�)D�ʙ����l���#RG)��C���Pj�kH�K� ��V��N�cAʔ�E�L;�}�*| ��)R�U�)���D�Oir��i�R�� ��+�X���x�	��}�� ��$cp�o��2[��g�֑+ ;�
�h�U4���t�
Yg��\�؜,aG#G�d�7'��_���K��U���4�Ki �˥R+�>���8�=9:���e3X?WF�Ɯfi���a��X�g[�H�e��%o�B=P[�V�.VO�D�O:�7�3oK(��;(���x��0Lu"*M&56mm_��nG�F����Gvȥ���&&@Ŗ��H�O��$F�@#"0r��8pLC���V d'	Iy.<bd��G�J���$ߏ�kfՊ�4"W�x�m��d���7��,�>eVѹE�c1~Z�g�I��IL�ƈ�U�u�Ep�~�ڪ":g_��j�P݊�ȧ;w���E��@0�uc�R)\ߡ��2��b�d���S4��T�mB�B��$���*�ҋ�/�V����77�#��1�fR���R.i���~������W�T�q%�z�X�j�X��P�������|�:\�2⦍6i��E�y��B��6�Z�ދ�s�M�U��y|[��^gh���u,�B���NGN3���≽K��.�a����ª[�AwR&�F˅gl$��˹Ĵi���G�,;��Wj�Z��%�l�H1�%�y���F�����9Cb\���eo	�F\v�Y����DX��{[2A$�T��xk�^ء_$2��d+���q���6�
��e={���А����� ߇����6�������kę0�҈w�,<j�1� "ζ�\��6�bH�pI��)<��X#N$���n���q,A��\����V�bt�823�*xBZ��we��9�%JV@8��{���H�<��h�^<*��A�R��.TҊRc�O�Nl2?BT�J�����sZoc�l���,���H���+���mLH��0�w�� ��S
��t
f�3�^OjcЫz�*�ؗ6�F�$�{x��O�e��x)�"��i�JY�#N��Ҥ4'R��o���x�%�$v2
h����C7M��c�U����0�F�P��C�"��|ȶ��h������RE+A�J��	2�$�` y��]����DHs��֗q�8�3�E��^�����u6�`G��#�>A�_�	>����/�W��oq���K\g�FWg0S�C��!w�8�<b����x"�d�z��YN�h*��:�I,���xR-�Jrɖ��Y�4� Tt�/��l�\�ÁN��aai-��݃�o�O���O6�O6Ҩw��"��^?��2	��)۹�r:���M)N&=�TGPY�����k�`\`ٳ���}�5Y���a�I�����<�N�	؍>�p*G��_�g�%;�/��6+����A��.S�SZ�[e�&��b��e#)=ۢĽ�P�@gA��%�|�%���<�v|���g3�&6�d�n����/�k!�I����̇T*	����B�R�tz��@0�gf�YO�IY��.D�"دQ�ţH�N�0�b3�E��(޿uG�S��b\0r���w�T�sZ=����ʿ*�#����7�����oUuHX$Q0 ��H�	dc��I:$�ͤî���I���nz!	��%fԿGw�p�Q�mfpQG@PD5�{ouUw:�������~�+'u�ֹ���s�Rx�|[��`l�ރ��c�~cXl)Thʢ1�c�r1�q���u��g���S�`;!�O�!�Q�[�x�,��N�/JX�3/a�a�D�?x�7@�U�bKX�m�	�ly�4����cOv-����I���X�O��FX0��Q搇���U�ȟ»����A��t~��C?$���Jn��5�\�jD5rʋt��MO��m�6��h�`٭��VSv��_��ߑ���P�oo��O2%�T>�M�a�*�繆Ϋn�����E�������6� O�������(k�lQ�����x�:R�Vf�q1�3}�N,�aF&���U%>̀S�l���g���"�h��:b�ݒ3qg`�{������]Nu�9D%�mxr����U�I8M���ih�}�k��Ƞ#<��M���/�αvZ��S���J��F�=��N�t(-�j�ڂ�"��b`S�TY�-x����n�-�2A3����.��^Oͳߡtx�'n�m�-��*Uzc��ܶ��Vl��o�����]�G���}�������wu�2��_]���8��٦^�on�g��H��#1�^x�ET3�K0�Z�pu���;�e��H��bW|�[cW~���N?P}���i^�(8A6ubä���*V�|bh��i�.��]�4�.����x?�3�n�u����8%��Þ��J���`\��V��V�*2&&�����W��:��ҞA�?����������rC��>�фBfgq3����l~re
MT��d�e@.k�«54ư�)�ֻ��{���,���UrP�����d�S�o��*� ����N�>�Mׁd��d�w�O�賣���L�≐�w�iVR"fe��'�P�?6�X�%���F�
/C��'�%Y�&��3��`���~[�T�+v�Ǆ�'Y�}i�cW��̎\�o�"�|D�~�ㄈy|�$���F�羑X�m��69�=���	�.aƎ�O���W�h���ѝO�G�7i�(��P�'��'�̅]'�?�B��SDY��Α�BV!i�]3R�cV/U���J�y%F��-x$>Z�[�'�;�7�/?vf�!�^c����'�����o��&uv�����]�C��=���jF����M	�O���l�6���d-Z�&���)�߹�������:�,Q?���/���Q�l�-�����]��i?<���h�:/z��p���^t|�u1�9�zN��]x��gB�E��enx�=x�$�h%��4��G��s�A���0[\��:/�
կU7bIԬuʩ���� �PFN�c$VBZ�� c����igL��h\�,��^��x�z��Y;��#�(��EKY;��#�h�I\��u���00l�E˰�1�<�;~�ϵ*7��d6�L�)��`ۉD���ҹ?���o己+o�����:M��l%~@��:lL�a{��@ǋe�h��X�)mQ&$g�O��i.&F�g��p��b��67Y�f����l��P�_}7p[ZQ�i0����J:�x�2�	�[�G���i�{-�L+>[b	�"�;�Uf�n�Y��g�<,Kw���:s�����U�#*�TaT� v�ϱ[�	%�H=!V���If�`J� zb۠���!1�� =����9x��ޓ�
����heS�iF�Iߒ'
t���N�@M�����;]���[^1ԑ���.�-�/�~$]2����<	�=���i�%{�\dg�_�ܕ�)N�s�NN���	��J��-�~6�j�'_h $xh��X�5h�����M�5�U"��X�6�V{V��7�d"���}F�D��?�ԏ* ���]gΆ����U��������=�N4����b�R�Bu˂�r_���]H�h��{&PC����r�д���Ol�ݒ�P�6����P���j)�2C&-�����2��\&��Uo#T����p�Fx�-b^���9�t�y����W�G���L���i��87�)O���gu�:y�K� s.D�<��/N~�\J�[���~"��@d�Z���VKL��@�*��_�!O��"��h��#�]�.P>����9�r��\˩�@��&�]�{)�$�����}[N	�+Q�=rE�)�y�)C����P��	:#
�|��̠��͐F��E�(�u�X���b���Qڂ.\���ǅ$hJI�leU������഼p��M�t+_��t��Λ�G�I;�!�X��k ��CTȆ̙�(�w��c�������\W�V�<���
�3ی��r[v6�Y��7в����(�
����ɱ+��#����ؤճ	�O?�k:�ޅ� �/LH;������v?�Y8�} �j�χU�����[ݱ��(ޑ�0/	���YY}L�K Z��^����3�b$�`0+9w0eؐ���4'M���V�� Hf����ƶ
�ej�E]P>:�
�41>�x���@G�����?#R�,*���X��ճz��;�ѱ[���j��4�������%h�e��M⬡�O�5��չ������lm�L���DL&ʟA�#'�H�게����SB#ZK�hv�g�ȑڲB~��7��F�b>D��3��崁u��[N���nu:�?��C�R:�O���t��	c=������C���C�̰���O��Z�\����:�a��;W���ήO�Jh�J��k�ޙ=P��?�y7-
������$	���z���$�;����ԧ��G9��,��D_����d��}]]GF@>u�L�uJB率N+�����F��� �7M�m�! ��m�j���z��ί֣@�Ȥ�9�V�ׯ�55�"Z+�
�r��=rI���C0_����/Kp���.���,J�mޘ�y	Һ�)����@��L�ӆ��H jo��:�?p�C
���|�^ ���'�'��A}��ʖ�����샭!��	�3wa���pve�o��>7;-�[J��P�|!���u������ۚ�K(�,y�k��?n=�����n=�c�<r��[����$���d�4�������&v^� ��[v���Ų\��/���4��iB�񧮉������DSF�8v��ʊ�9!��haЂ���t�4ݥq��!<z��}��ˠm��� Y��yƢ��G����_�c�8�ISt�%Z����G\'��IP#��CRN��_ޣ��p~Q��/-N�?��!*� ����j<���Bb��Y8���P��z\L���Ʈ����y�!��tzf0`:R�;FJH5m)M�ێD�LN1�c�'�^�c˛T1jo��稾�	�f������:����ŕO^�$���2��/��^Ĳ���)��]3Zj�W�g��j5�g�L0�#�zbM��$�"��v��-_n�N�ql�ϸ@2��~�!ףyC��eG3'~J+'6�c��,�0*K�;Re6�Y���?V������ e�mc9æ���M��7���GR+�1���A!��#�yc���Н�vt��Z����R�	R��ݭ�>D3�όo`��y��h�D=���mU�x��N8�4�8�q�s�(�n��={[g)���)��3zBg�Z2��$Y�
x�i�j��M��E��U�J短S�;y"c�m���k��-O !� �!r��4AD�b	�t�op?3=�zp���@%q���J�{���R�I�<l��}�����~Q��s��ѫ�o�~'�3�dt��i1M1����.&�wi�����a�>�>����ϐ�%}W��������9o�y��������؂ع��c7ľ�'nT��8%nuܣqo��;7�����o?�0x�����|�E��n�(�谣Wm?��ѓGc�]rlck�=��c����߿������p�w�p������?�t|���ǟ?���������3O('F�t�O=�b�;\�@s��j��k�J�������@c�Rw��pj��J��bw�����bw7�W�l��ں:G�����x1��Ʀ�u��fh�!i���?����y�� ��������`���!%�A�����E ���� ��
�	`��A\�!� `�q���)���r� ��w�6 ?¾N��w�x�G�r��B�r����<F��t�S�i�a<�_)	Y�|�+���K��0��q��N�n�7h3���)�=�yܝ�"�6������^���~��Z�s�nǹ�N�~�~�~�˸�5p�������;�};w��_�w_
���<�����V��opw5���n7�r������o����/������7ܽ�ǹ�o����?�a,sw��w���ƪutX��}���݃����2���;�S�{,��;�E�]n3w/ �B������vr�5��s�M�^�ݷ�{wo ����۹�-p�������} ��x=��jy���3jy�������N���=�rw�p8HW����w��k�^��V�~B�ޮs�]��J�>�sG���o�|��8w_�_�{���W�[����t��:���6�c8h���Uq��Nbx�w*���+i��������;�)�r�^�W��`}�^%�l���{�M�������`Zj��q������O�^Ģ�~#��;�n ����#	��;*2��?^T��!e99�O B����q���MZ}�瀃�p.��l8�'%,���tu�Qݞ׿
��?��O��1$�O�#��q�w��_)�_)zLK�}Z��Ҋ4��KK����sC0�i���C���Y4V��	au���,gz8qi�I�#�NW��s�B�(��U�fNE�,������x����Ϣp��xl=��'}<��h8J8D���	G�[��!���'�BGKzH�l����C�1���x�E�YOD���!�{Cˮ9;�(4� ��G5��C�����Z?}��z���pv�p���,���=����9���Ғ�{�g�ϰ��u���6~��g�'��gJ~d��֦�gfy^�O+Wy8q��{~�z�	GO4O��S<����d�΂���}�?�~B����2��3�s.8�R�+q��ׅ��p΋y{<�IR������p�bޏ��F�#�N���g�	Z�6]Cp��p��'�*箞pj8�z�����l�����d8q�����n]<�{�����=�\����yt�=����/�T� <�~e�K��#��AV���"�>���w�U����&x�p0b��wt��⿣N��V�{�����%��n{��o������'/z5�ly������tT�Z����6��T�\RUn�u��vo�����}��T�<����F{I*R,K,c�W�
��᪝og���Pd����Bb�����^k�;��ex���쮑��N.��ɸ�rM�e�;�.�r�ր׋~,�n��y�c,����v�o��᷏����1%4����V��H�oo�-�f,���i'I��B�n�"W=~-C�{�n/����Z2�4�;\'��&M~�'4��j�n�O&V��elD�)���j%D�K0��z�&�����I(���WZ�{�@�����n�5�n��E���X�r�(�kIr�v�������^Ks��V�3	ާ�𗖌�&��~ �M��oqe����`'�CAH�fg�,�4�N ����L3223�g�e��06k���ҀU�Un����E{�J��*�8,�PXb6�0�hZ��X��PSЎ��P~{���s{-�fbwو������n��p����Ը���.��>���,�U�!��1��2�]�WY��g������J?#-}lj��Ԍ�rz椬������	v ݌�qm�q��[ƍ�Y�eس2ǥפM�hM�?�Ԝg��%F��+�
ͦ*�s9<���kj|v���=~�K��K��:��Z�:�W9�a7�6��a�D�����^��_C�c��B�!o3�5@�o��U���)̫"�FJq`�6k����vWݿ`\1����E�;�J��g1�F��	p�x� rF T�ܧ��`�����Kȟ����D�L͝!���/����#p�,�n�_���-���sg����6��~x�߷�����a�՘��f��m��o��i������Y-�Q8n�m���9�6z����'r;�}�1H�=�m��m�8vs�Q���C�ǟ�Ǎ��{��4��'sܽ:\9B�����r�>�E���SJܧl��%�k���}J�}J����<	p�[���o���p��Ο��)��b�} ��Yx��}����&�~/<�w��d�W����-W;j	�H dXCa��� 
�8ݍ���Fk�.�N* 2)�
E��J����%y2�NRd2���j��!����(��Rb)!� ��.��N=n��+���G}������������� E)�<Z�% ��2��$�+��16�����1l��$�&%�<-�c�e*t{V?TԊ�n��v�} :�'�$fԙ���[��&���*�V��k�}�:{��b�9l6@e~O�O�.�J�S�o��\V����ԑ\|I!)ї����WYRXZB*+
Kf�fSq���j.7�d�[Z\VZ	��9WV��Mr��� �D����*��L���Uj</HҲ�o��kd�E��un/��6tz��3�ÀP�x�2@
����AMB���*�a����@-Ax�\�J�)P5��N�S��iHF�{�v�ᣴ�^k��,M��@4��_NF}���AT6{�4X\�2����W�-�̓�� !B��߇(_r��s�6���F��%��T-T�<����L�
s�/8��:�.gC����<��)>���MP��HD���P�2鯳�' ���)�6UB37|~���&b��6]��jd5����L�f�4����i����h9��67M�����N��H8r}��鳉u���js�}4*���Ũ�'�!҈�j�f�l�X��\�9���l�aoU2`IK0ˀ;�SӤʜ��H�Nip��񠨠���d��?	fB{�.lB�}Z�:���L�Q�S`*7��j$>;��	h ��8�v����%%�³0�cq��4�6:�6c��4�K1,��1�	te�F}r��Q�$���B�B�nz4�P3Lk?<_�zq��u�}��#���;��QPFA��� �
��k,H��	��Z��
�˩���/G�K����O;5�^{�R.+D�r�;���́#�D��1��H�h�4bF�<MK�A���D߈n)�k.墔~�0D�0I](��	i��.Gņ]b�:0YP��j�7�A��Zmʱ�����v��B:������i�������������q��!r����._���R�XM0�M�"&�}� �3
̔��A��K+��/f��h��Ơ�q�yi�H�E�6G�^�*��͈Tm�2��G��K��s
K����i�k�Th���&@�=�
е=�DZ��Z��͋R��h�Sm+�`g' ��8V�s
��P�SѨ`�6�(�g����S���sHE���$Q�a��d�6���=E竺Я�$�4��-�R�Ac����h.̕C��^��ͅƢp����b�g�2Q�y8r�fcN�	#����D�c�<*�L#SH2����]�..�ȳ�͕� ��g�6	cb��m9-�=P��Z�-~h$` AY�8:=�w��WqA�YdT����H����=�����&0L��	o�P�$����������+�"�q�m�q@��� �18���
� ,7:Pj�ɺ
p��,ն�)ԟjFj���x��t��h�q0NTB���;W�� �4�V�ha�����W��h:�E@�_5��8X�ꀯ9�$:��X�4�Q�N��'d�~���B�,���~]{�D'�
��G����t�w~� ���Wʟ �����r����W��U l�p����^�8x�	)a4@I*'''8$CK������k�(��	�R^a���$׬�>��ho��#�:�c8b���'%��
$P����q[�H�o% ~�ۀ��Q/iH���#�v��R3�1����۹������ʸ!�����T�����3�%��߼��G\�tY����N���s�|���^Ԑ�*r��
g�p �QT����+::���^&1�L@A5K�:}�P�Nd� ���R�	MerZS��	�Tg����U5:\���zOb�\�����T`GW�^�t5X<Ț�C�2�v�r��Vw�ɇWh4wE�˚�:(~&b���n����Xs��M]���{�����u�*�e)?�t�Y�u8&��{t�����f�bC�e +I7:�n���>��Y�n�m�~%��#3��ɜ�~=�?��_�&��'a�X�c�WV����?���zx'��<v/�?9n�y��B�`n�ua�}�i"����ߤ�?��Q��#V���?�[iv҇�}KmP���-åך�����5 ��Fʠ��l]�@���o�l��=�8��G0��PPg����@�jQ��&�w-��0�ׂ]��ҳ�D_P����.�CM��K�����8�� v;�vR�r��ЉRA�YM��,uP~���{ X�auA���ݵ�Q�vB^��oN�����6�B�� $��܄��X
^7�k�9 �g�S��8HM�I��@�c@��8u; �Vb�[�P�%�aX���'���?�ô1 ����7�W��{�����inrK軮���j����ne���Y����;�;��wk(�{������"�������%8G��u@t��$N�DfW���̪Z���*Q���eH���T�pMF���^�p�F T
-$Q�J:��"�S�F��gڙh��BPxQ9��0"�:�r;=�9 E\K�xcs�Z>E�	z����X�����~i�v�}S�����F�֣@����@��F5�u9�I�un�?�4 �����̭CKj@�q��AQsx��m��[6����������ʠ��J6�"�-�@7 ��~EH�Xp�n���������r�� .8F/��8��2TSp͈��{A�@#�T�y9�GF/ֈ�JI��mS�m)��d���W�h��J_0-�[��X��I]��$2�������4�Y/�q��;��7(��TqT�2v�$��2^D͈�٧�ɑj���04�f���0�Rnu�I�V;h�4��`�XfM��9����:�ޖ�h=�4a���6X�K�c"�h���*�Έ�\��%������P�aq dq�aJꙨo�8e6���"�3�5�HA;d�)��fW��lY&���:��*���( \J���!��|a��"��h&eM�=tAlu��lv�X�h�1�j5jtD�PMa�nNCS�\������PchP���vu��g�v<�5�y��gq�4jd
Zp�f�H
M�qT��u���䖖����fS�LLsM��f�b�`�F� ��:����bSn,�0Q�d33�VS`ܝV�IK���,x������ �\�AEj������.\$(���9�_8\�� n�e9����4��3=�.�� ��ith��~����Ź�ǐ�j��J����yx��p��YPw�ޱ�\���������?��}�Q����y����Z��A��3���0	�6��|���Td�7�ԓ���+Ll�h�,�:�
h�5~;��do4Co+.4�+2���޺9 .�PL���}�hpA��`oQ��bU5��g9I�2���4:9��L+jܪ�2�Ҍ{�ْ�$�,����k}���V7R��L��f����xu<���Y��5õ�,]RJ�&�d6�hox,�8t��p8.�&շ!
J�g�/�A�K��]J�gr�.}OhtpA
P��͝z�\5���h�N���g�NsP��Όu!�pƚ�B�X�g��Z7�m"�h�6R3G�a��4T٪'߇��,V�d�*:v��`볨ЄԄ�3���~�e���ݩrŕEzb�IYu���TAtU��5��{nё�v�W��+�u �pV���,P
��ۏJ���_^Z,�L\<����2]U[8R���*H�lƅE:�j�����2f�2�G��f5��N��|>Ъj�4a����A��z�Y{�lcnee�9㝹A�ʍ3�����5�F�u�@7�Z��OrL3
K&�u<2���
�l�P#�eˀR�����Sҳ�e��~��)�|-�8���n�ԑW5�8��my�jO
6nz��<1�,y�1KH-�]�H9<�ʒB��Κ\F���[z!�&��K�G�T�@`-,1����8��ۓ����q�*��b	�Nq�H����ʿ[��
I=K&�G��A�(�{f���z;��u��dB"�)49�b@#�p��.D�p*�EhI9����H\P�����;�[�T����1`6���ț*���z,I�ڽn\}���~�H��6 � �����c�h�(��w@I�{Pi�y�A����zs�=�,���*�.8��Pyf �������~9p@�:x@q|}@����r �ox��e�1x8��;(o�����Ae�tPY anx ��e�� )G@�������[fw@y@ 8�	������a<#l���$����3���d(L:u@ٯ�e����g�� ��_AY���p���Ca����(�A�?eX���Z�w ��d ���S�����	�f8��p�P�zP� pk<��q�*�>�L�|`�蠒�2��%�{�~���w F�s1�i���/�� N�_֥�&x.�:���п��9�,�>�$����P7��]�T�t��"x�fT* f��yPYw��IrH�r2�j&I��3��zSJ���k^'%zP�c�TU0q�P�B�����N��6$ ���?���%~�( � T�]']�׀�8lM)���~╣Cp��G�]7%���Q
�_�)8��F�l>�D�KT��I�}��s����,U�TW
�� u� 	3������p-��C/�Kӂ[��M �Q��奬I}E�n�f���J_Ƒ5#+�x
� �נ��4�0(�6���]���k�x����eUN���U]��.�c�8������מ�E\\��ɣ���:�I�I7vl�X�Xb4W���24u�]�XZ�:&��ׯr9��T��u����-8�E	���p4����%����h��է���42 ���-����!�͹q��[�D\��[I��FSE)�
w��z�����p.���)�6�m*h���Um-%���Zk����)����91�=61M���ٽl/�J'�7Y�$%RR*s�t1�9IM4V\6�Q�k��Y��!ګXYpF�����Wp�n���˻�����1����p���K�z�U(K,��v:wB�ŗA�*���=�\���u�j�^ oꆭSYH�����ڗ~�j�Zs���
��m:�{0q�a�V��W�Ǟzր�٤�6�u�Ύ}���.7�s����I����K��7�Y@�|�3�� ��Py#hpU1�Bo�����liM= �gR�{u��X��v�֓Q�F�-y���݀�嗣��$t1Gl�T�[>��P�&_�|������3�'��2V�����<��Un�f	�,���\�Fhi�j:M�
	K�$�����v�����@R���u��7Nס,ݡM�PāJ_x�)�C��Iw(��fJ���� ֌eܘ�ؐ�tQ�����2�C�ޡ<%�8.ա�!��:��v(��?�K;��!�A��e*�wv(- �  �f�rs�q	"rA����q(�	E�1��Ub�7�ʙƍ�V��$��.8�O�e�ɧ��7jH�-��1#�&8�D�l��0̌H4�X ����@%D]+��P�buq�t��c:�A���Π����]m1�ۥ[�`���u0E|n��.���1pA�W��K3lڼn���d��9AD
Z��~��0���::&]肋E��&d8�"l��fˡ��0��K^ �;�*Q�� �D���5�.��IB�H:Tbh%v���l2�᜗_61�V(M���16E�,�3�M)�
xE�lLA[0�*�1ӆ)/t/PX�,Zl�G�q������.�e
��ghK�G�ӏ��$�ո�f��Qh��%�L��� _�%6�xU(���P^ 80���H�Jx~H��1x�N�y�k ��o,�����2@��p�p��-�[��l�Pn��O��! 'l���-4ς�z�6~����n�P��`8�O�������}P��K�� �� + � 6����E�a�Y��+,Z�R��wf�~���T�����/�~�[�UiqW��� �+ W�X�gmQ�����#pok�P�44��]��bC�r+���u|�١���d��;��>W�3��Z�z #�@ A�ʋ8�@�u>�o��C��ݡ��f�w�C��]��ޕdri�nw	@��e0����'yxL�Vp{ 
��0�s��i�~�_u�2�|.�@�Y`@&�[s�m��9�8Y	��a1@j�FO�5w���cA��h�mtU��+�}��P�j)�[�p����!�����v*�P��  \	2@땡�+��Y��"�O˙;�����~g��J;�/JY�M�̿��  ; r�Y x�h����e
��C�q{*�8����[4�8@�6��P?��N���P��h~��~�ˢA8�Ȩf`����θ���p�R���߫�����!!sMI��*9p�ls[���"��l�(�)2� �a�
��L%t}�#l�8ۻ��eYM����������:\��?�e-��&��������k�Dg�ɩ'%чۍ	�؛
�Y3Ȃ.�0/����o�C�H�qG�p��+/-�%�Q���ę]h��C�;,ptx1�l,�Bי�2�^k*V�l6\�T.��6�m;�� ���J��Z#և*�c�"�8���!u�?�)j`�L�� ZE����
��D�+��pP�+-�sKK�
s�A�fa�
1�&�m5d>���9��e��+��2\�we�d�7|ݥg�U8�-];���n��x�L˅��
K OŦ3�[x��lW�mm��*Ab��E�$��>�LB��q�`i�Y�֨9�o��ƪhL��������PY�uJ}#ST�O�vJHW�FS$w�؞D�¡�v�TtF*��q�i}�!�Mđ��S�?-�qjHK	����#�#���V��>l�n�S�\/��lQr����n� Q���-����\,�O3���Zh<ȃ'Gl_�IB�m�T-�}CS���d�ME�p�[E�M%y�@��7�M:8aG�e�T�P��r8kIL��uY�n�Ut��&�)�%ڮH� y�RД �Xxni.m����m�����\$�E��I�7�vXЌ��0C����~�K���Pam�#�m/�(AOSy���U�rS>�Y�k�Py;%uŨ/d�XXT~)�>d�	�(B"j����G'�g�?�t}7Ί���I1������!t�2�>�#eќ�Ŧ��`#�c,�nk�B纵�lzƊ�U.�@�Ut���?R�.�u�:w�-g�[Xa�H�> �����;�ϐ^�w>;]�������
r������F��	
p|O�n�R-]��c[Sr��y`f��:J����|g���Șk
H!���Yk��P�HVǪ�)C0��}Fx�n�a��S���ҧy����4qn���U4�ܛ���]@��9�XϥZ��TH@���K/�d�c�1���0=�4{�G����u ��Q���D����²�]�8Srg���E���䢐��� E�3�!��䘡H�Dֈ+Yח�Qg�{�g@�^˱yG�H�-4�X����e�LO�R61�1rRzZF�<
�|$������z��'��
�⴩�e��0R�eL7�Wf���+2 C~���LJVޗ�+�������bm`��3-�1�am,��A���O�����7�c>u)#*O \g���=�\z//6K��"(�h�?[y��8m���"��C(H�L�z�MaU���؃�3�^��At�7E�sV���J
g �s�+4����r m;n�	��T�L77�}�R*]�����×��{T}�o�����<��j![H�.^���B8&8�L)����$S�Rgs��Bc

rg�ӄ���1��8AA�lqQ��cB����m�+�A�1CU���@}GL�����a��7b JQ#�㧾#��.?fjr�7,���x�&�|'�Bi���ݟɎ¡�j��R=m���S�TO#��9�Ǐ�NJ&zu*�v*I q ���;s�: �_���<�3ȈSco<
���3���P7�z"���j�uI؛�u5r�;�]n�����>����1#�1L�w��Q0Za�yE�"4����Dz��0��b��a��%-P:�����D��<5
D�:H���t�P
�/�нWЩ�RU�S#Qω 5~_f��K�8r�->k�k�#��
]S�*��DMH��&���4I����B�Z�TKR}IM�GZm���3�"7a�x�6�P*K�эTM40����"����<~��I��-�<�I��m���Ȕ�d>4��o.��8p(��2���MhU_t��f E��$MvIfcV����FR���^>4�@��[7E���K�j��|�L�ZkM�mz�&�pɞ:B�AҢ�����)�Hy,�0�KJ��<�� K �]ѩ���	<�S�	Hΐu�9��K�8�v�Il<Н�H��D��e���kI�2�8�>��P��]�붪�΃��L���W[�J�D_�x	%�6���k E+!�k;�\�� �3��v����]�=r�;��xޱv>O��R��t���a"�*�������u�:N�m�; #�3A��N����>!\P�������a������A�*,��?��t���-)�?�Tg��J�U�t`)�������:b ��NbU��a���7l�z��^p8mZ#h�dS�2�;P�T�Z�;�g����\�B�v����	�\�{�{�{�
{�ϥ����݈��}u�_s­��Iל�3������N�2�� V�������n�սO��z�r3pe���	0~m�}����� �]�|��{�K}2.��UځR�G����Q�!ڱ{���W9230# O�F�V�9z���t�dU�[ZTY\RUl2A75���2��2#Л��TQX����Lsͦ�
\
�}��pw��)�U�SE-A�b^��T\Ul,**�%���*����T<���:��	� �K �|�3@�iݷ���n?���=���G�#�:��FD�������s�=%^%CT���}��;�l��xa���:��K.����,!��Iɣ�HI=&-=#3k��&N�<e��ٖj��^S[�P�.�g���,ilj^�`�UWW-���5ˮ����7�زb�M7�j]ݶ�[�������;����?�����w�������~d�_}��'6n���SO?����ŗ���ʫ�^���;v�z��y�o�������Ï���O>��_����}_�������C��|��w�>z����x⧓?�:�˯�u�y���q�r�}�6�E;�*���o�޳~����ĽJ�" �r�� �'j�^;�h�8|F�$���-r7ڽs��TJt���W4Qs�s�ѹ�7y�?�{�X���iaX��4���͎��]�gg��:�
��y:�:|�`���h�0z��g}�����c�0�\v0v�׍'v��/��G�
��
���A�i��먆���ݽ"`������Mt�c-K`<0�{P�"��OO
%��kn��fCɄb�j(��>�h��<}����`�?Ф�k}.��a���C`j2�<�!v�ǈgSkO��!��n�n�,�(�k���蘍v>5X.�g��"Ux��s#�O0�g��SҚmi}Aϲ�i���q��H��J�cWf�ҭ�.���#<�����M.����?ȁT8�v�*��V&�h �	9����f����SS�[V��%@�X�s,?�l=\�}0�$�Q�അ�$���:mx5�{�F�G�A3h��Y���Kl�$�qY�Ⱦ?���Ҁ���|U˾h��5G�]�[l��A�P!�ͤS��B�ٶ,Rp�8�i�
�΃|@W���� �#�^���p	YJф,&�>�\I}	i$�X�x�M�;�"1�G��8"�	s�?1��@D���%����[����B<q�?�D�������#��ğ��ʘ��g�מ��DR����4��23��T\L�����;�q%��EE������m�`������Ne�~���S�@�;Z<�d���;p��rp�-ݯ���W6��8��<<���((�9��������
s��9s����@>�(�g�>��=��N���{��O�W�v�U��9���W9���d9S�������3�1�()J�K����t1�+�]
��s-���ʀggrWp?5������r���s�Ä�3`ف������~�RO'2н����.3T�q�,jLt�e03����r�R^�`��t�Z}P��>`E��N���>a(�L���0�B���{M�8���v��G��������t?��C�$���tז�����<S~Rbp�7a����oZ��B�1u�N�p.�D� 9���#ɱ:cg�{���P�5��4EH	r�mƊ���n%�e�O�:��E�o4������ _�H�
�} ��pq���� ;��?�rHy�C�-�^��� N�EC� f H��A���>
z(蟞,���bz��$8��o��q��;p�4�o B�a� p��CJ��)�c�k���IR	)'ń��WK���<d !ͤ�G�B��?��z���5�J!����d��A$�u�"B�)S��8l<Y@lC�͓�����G:��_0�-�����F�	�:i��$r1�==��J&���(C/�Խ��^�����W�� �1���K����ݫw��>�(J��.�ݫWT/xآ� �ѽ���m����"���R�y�h��+&��~�11�	?b������zzK�D�b���IH��ຘ�|&��$��%��d2���#S	�i6���,�ÓI	�����"��v����C��#����y���mdy��G>$����>r����9EN�.%�0^!$	�B�0Q�&d3�"�Ja�p�P-��-����2�EX)�,�n���'�zYxCxGxW�@�X�L�R�/:���Q��� ���~��b�8L���৾�M|�;\�H?{d��6��(��3Lsˊ�|�"j�9Ff�A�=������r|,�0��5���A�a{��if=snnQeE�l6��Z�L�[�\��[
�A�si~~�	7����%����2r7\�yi��ס�9�n�-���rL��K͸�p�)�%f&\��W�2{8A;F�Î�+,.6��#~g�����X4o��Ϳ唖��$_B��\Lm�h��;��R#V�����\�bf���X�H�[^ZQ�f�\Xl�0����U�I=|gSq� N��Ǌ�
�
�+���.
��i��Uc_y��4���,����%�����y=���֌2�ԍ�l��1b��Ƀ�W���z]R_}����[2�am?�}�3j��r���X~�+�z���Y�������7]�̙i�'\�d���ƼK'ؔ�Y���Tm2�D7zS���H���)���������W�`憓�y�tXV���=�\!�A�%d�E�(IfX�F�iV܈><\߂R`uդ��!�2����
rY{�Wn����\�%|�u3���H��e�1��&C��I�#q�8Y�N�O0�d�t��p��!\������3�{����L�x�Pa���m��J�NZ/�S��z���dp$+�V��b�����?���(�b1��(�|�|E�"��=�[�еH��uĐ?
E3�NǄ�_Z����d�d�I_�����;�ݤHx�G����������Q��>5�C�!'�]�C��������b�R�;�s�:e@�kԅ��6C�������p���p�a9����c�Wp��#v�҄��Ϥ]x��)!E
<R!�[,��H�_t	ۅ+��a��!ȑ���2�4�2�k�ݰ���e�C��j�mx�p�a��m�L���7�e��w�/�5<`(6�1�`�Ӱ��5\o�5�1�bh3���s.C��a�1���6dr&�t��g�x�XC�!�p���tB�F�Nʔ��˥9Rܿ��O���1_� Ɖ��k����.�a3�j��0R.�ɏ]���&'���|����������=Bz�x9���>RҮ�J�Ii����T�ri���$�T+�Kx�,Js��n�~��J�4[��fI3�"����'��^��X*-��K�������
uA"bo�6��k~������^1���o��i\�R v�����#�Y�--�!�����\���R��NdW�^xB?�ŧ;��(���
~逈�GԵ���y�/��!ޒ�R\~�%äD�2�у��N����5�5��7�7��Bj~<]{��OX%>G�ϜS}�9��O��������琼& \�1�N~ߡ�0U2��; �b��Mz]�.�*�"�,=/m�������6I�K��륛���
�E�QZ.]'-�2�ti�t�tL|DZ*���_��a�Z/���I�J�HwKwIwJ��,���WZcɭ�-�i�t��&��Z'�-> >"~&���W�>�_�_���7��;�7Ŀ�����.�����]|M�%n?����U�xX<$__��F�%�E1_2I��$��'�xJ<-J�(	R?�<�"i�4A/��JQ�A(�.�ΗzK]��%�M����EzXzHzPz@�_��vIoJ�R��D.�R@�K3�<�)�i�UZ%�,=+>#>)n����YZ$]%UJWJeR��-M�Q<W:)'J����/�ϋ[ćŇ��ſ Gl��G�]�M���Gq������(��6q�x��Rl�~��	����ه�ċ��5tؠ�L�_���bSҿ`��!:���,�֥��֕���t���{�}�_:lHHd���V��4o��4����Ʀ����:�jXF&7|���vϊ��)$�����K�`��{�Yk=�=t����x��-�ȴT6y�ʛ�����ekV�Y�.�:�`F�!�Z~��A��!�����4tXH������~G�1��ʾB%�=0y�K5�V����<$~��)�G��^m�4�>d�!�Ņ��M��w����������o��C'�1�}����l�֖���_,�z����q=Y�>��n����C^^��ڦݲ`H��Ïڿh��22��޸��A��?���M�7�D6X٠}������K!�˪���X2��kgd%��/���o���c��oﱚ��<��7 i��!����h��j�<��Nb�mܤ]���֞#k�o>��f
���h�P�@�/<��6n� r�-;0�XHtȠA������3i��	:���B:������)�!��ed�؞�qӫ��_��@{�2�l{�Av�۶�gd��oݸ�v���]�!̀�Sٺ5~{F��'�C���	�k��ҍ�>�������?h{�ѡ�6n::`�����/�
������A�C�~�>�}��k��M��7%��k�;s�%c�͏�o�1h��:��1��{��8��q�g��a7nL'x/Oٸ�~�!�a\}|�ab�{��Җkr4�q�:�wӠ�Aqy�^]Jz�p�4���3��w��x�yw��������6ݸ������� ���Λ�qyU�Ӏ����K�׭��c�����d��O6�)<�iݽ�g|�y�f�����=O�;o�ӛ�=�B�[g������)������ג׽�ں�|�/_�׍��֍�����o=��9��l�u���[��n��ޞ������������w���m��?��s�����A{� �8�����6�T��W�}���%��p������z?2@�,��Ы�%i�0F�K؅v.vU�e�W�)�@�'ϑk�k��j�� �cbd�8�P)�#�I�+���54i5��=�ˀ�hO�r��X*6�[ȣ��S4	���$���'�$_
�������B�1l=�9g/��f�P.����a���3�+|G�|��@W;O<@VYZY���%^Ӆ6��]�r�p��O�Vx)v�p��G�R��/��Pg_=�,NL���w�q�t����X���)�B�o0�%�U�&&��n�)b��M��H�+ExZ�*6�;����$C�Ieb��!���S=��)�i9��5PkW	'ɓ��B3i���xi$����1!^�?C���H3��	�:q*h��G�A�=q��$��ɻ��b�������d� ���d��J��
�3YG�%��I��Fq�8�7/Jo@��(Ո��3�LT�-�j�q��'�����B���T|zȍB"<���(�E�p�P
�5�P򆰃�Y�|"	o�l!��<�N�H@*�F0_.�z��i]�!F"�IX)l��q�qJ�;y�� yY)��Zq+���j���.�`�^�R��$ ��1O\�	��q�1w=��/=�Y��"9boq��p��V�"y�:�	su
��Sh��ˢ,�
yS���Wi�ƈ7���b&�pZ� ��O�`+����3�نs6��
�C�i�=Dc���5�a���~0B=�HJ�5\�&2��Y.����4 ��N�!�p5���*g�� ��8�1�Qb	��w�?�upO�{.��R��.��t�:��Xp	@:��K���Ո�ə8@O9k�7%О~��Xr
b���N�[�O��������o���R� ةŨ��� �v6�5��,X��³B*�н�]¿�o�$��������Sq���y�J2(�
���[@�$]�A*IdM��?L�o*��+(�T��0b�"�@��0��ҷ�5�H�1��e�0E���Gk�3R/�R�C����L~�!��z�>H�r2Y��t����RD��$��)�Df	� �D�	�77	�C>&�f�p����� ��Ň�oP�?��C�ۄ�ī�o!O��Q#&Eb;��K��2� ���)�K�@�/
�R���$kH�V�-�"�
&�S��o��)����j��5b_����Y(E�(�Xa��y�Ҽ��A�c��CZ�!ayE�怰��L��/�s(�F��l"�
��������D�|(�Hv�Ѻ��\C�^��W�:R&t@����H�MB3���Q �Yµ⻤]�>�/�"o�ǅǄ�;�%�u1�L'ÅH�P�da!�M�RA�+ƿ�2	&���o�Z�F����{d������,��hq�p��$ƉF���~�����&.!@~%�	}ğt�O��B?�)�V����',�#B��y��Z�<a��,$	o�˅��a�}�&�8��l����I�;B-��\Gn'��#�%ሮ�_���ar��G2C�LhL�z��Ia����W2H��1�b��#>JD��d<����p�h/.�&�ib�E����(�6�W�O
���z	�&��s�.A,�X�{�iR+\(�%|&��_�}|O�����71B��3���{���{���b!�66�wck�J���R���VT��J5R�B*eC�%�RQ��y�}ϟ҇�߿��s����{��{��߹���"���)�s� ��̼ʴd> ��}L�b�s%����yL}�̿!�@�$�q=��w��ׯ�M���}ϝ6�Wؽ�����	�����=���z���Ë�9yMf����m+cd��3�{�<�<��a�rÞ|��G�1�o.K�a!�ss#沏F.d�E�c�cdA��I�$[Ε3K���4����`9�<�i�i��f��<�⏧o���\�w�?�<{���}�}�����U�¾ĽĮ!k�5��	�U�Uf-4�k�kQ�E�/�u�:���[Oֳo0�o.�&�&�=���,f�f���eޅ��!f��Q�{h���'�'���a�?e?����ld����Dѿ����[�6f����og����������|@>�v�;�`��@�'�s��f�C�!�!�!?7r��΍�*�+nn�ܨ�ٯ��d'�%�%�<�<���b�|�Jf��|>�y~%��W�԰4��w�c���2�����]��������������n芏I5W��m���KV�Uܺ�u�>���un�H
j��ϲ�2+ع.���-�-9|���|�&�ك�A����~ ?p?��G}�?w��d�r����D~bd~$��!rn�H˟��s�_�e~厒��c�o���w�w��a��G��;}&k����s���y��H�+�`�yԝ���Af�:Of�O������rosorop�{�ٟ�ʸ�zN�p�+[�n`��7@�d�c �F���a�,��=ݚmŶd/f���h�6�$��,�I#o���e>��WL��3��o��lcn
;�]���ӿ����zq)��]�9\�/gr�l�R�w�}�5l�����������~�R	��5�2�9("6��5�KD�N#�G\�.�mD|D����".�hqqD��&#D�D�������Q���&�D����w������c��'��{�;� _�o�w�_�_���S��������_ϯ�7�o���G��g���*�~�#��������_�/���O�O����J~>/�8���z^�O���+�g�%�r�!�A�������������t��.>���������� ~ ߏ����;|o�	|:ߟ7y����5�P>����_��S����AN�e>����I~A�$:�� �܄:R���K�P�?���ˤ%����������z�1����h��k;ć�H�8�f=��/����3���wߕ�.� ��~�h+�=�W��9t0��6�I6���e9�p��F�Ɲ��1�x�cǘ�8����HǓi�݅�I�ӌ�'"/��A��9��SSeP�8o�l�J���nq�Э;�`h���:= � (rr`!ˑ�E�U -="���f �uI<�.��1�@��_5W��u��d�,W����~�x�1��������ollLLttTTTdddDD�=(wrӄP�`�����	!�G�	��#��x���U�/��Č�₌ܬqEy� ꉃ�7͙81�`lA^a!����x��3OMvK�}xP�i�~%�~Q�sr��B���D�d�$���,B}z�~O�	��\S�ѻ��H<���<�
g:��+�#�?��wh�6ɟyqr��ax��Ӝ�dR�=i���i7d�\H�ߛ�|�.i����ii�e==����l��^�y������cX=6+$���P�+^�i���������~$�"zw��%^tn����7��1�ia�R2JҼe$����B������{�FG5�y�L�)��O�SJ;������-�����L�ǲy���P��WPt�f�L�!-쩆N�;�񟬸�R9�Zr�ǒz�5i�]�F�o	>�Q���t��?F<���������Ǜ����7�#����kI\�p��/#N���jC�iJ��Q�z���x:���Ǆ�v+±������<QƹN]�g���oB��p�˓�F���{���p|<#�a�����D"���n_�p\8|M8����@�q8>��$����̨�q��,_���������p�����"}�p����:aA���K��y�d�l<f�nɧzɷȳe8��ip)���.	��C=�^����Z�r^�D|�px�ۄ�� ?�|چ��e��VnE|�p������$��2G���N�Q��	���D���|#�a�0Cǹ� ����|�A�y��Q.BO;�(�Q�1(�M����wí�#O��B���q��.Q�-�E�Q�$<ޖ��x	Xlf"���-�POY��W��//0��G���������>r������z;��<��yX��[�~ݷ�����g����שWw,K����|L��������¬��<��,o��-�.��H�4B���:��e���z�i��oCYv��S���~9E�_o�i�����'���qZ���_\�׾�_�O�rjS�_��u֢����n��뗜v��z�դ��^�!��-)6ԛ�>�$I��?Λ�O��A��^�D������t:�0_�CW�&î�}��+��Oa�2$��D�U�+/<s����y�`P^�6'+7����ŝ�ƥAoF]���7�ϟ�G��C��y���mذ�S&20oR镗3���̇!y7!27wh֍�Ox�)�d�����?aX\X�3��s+s{����n&�`�����	�E�T���>re�|2�N��?��)z� ��v`�YC��B1n*���+/�o�f84$�N�YBh��$^��e�z�/X��·�͂mn>����'���?�T)�Yřy���p�
��n��fe� ���z{������^s��L�;����H���_ֿ�� ���x>0�z��$�M}#�[Dd�tj.��z�#=s�hV�!ӡ�9����CC<�sh2�xl0d��]�f��3)'�V]�.����gKYҦ���Oͦ�@뛶�_k���%�YXx���n���C<}J?t*s81�����&�"~2��P����'���_T6{�����ǽr�2
�����g�z��é��d0�������y3�I.����А���>OѵCz�@dHk�y��=BJ	�{�A�`��g ������Y�t̚00�,��WH!k����䬱�S���@Ԥ���C���� ����cz:,Xz��砕���ɰ�Y����l�a�57�c�aa�ɬaC�U�=����r��;��G�Ҽ|z�\�j�_����@���_��@G�+  �Fc� �� ���R�9`�x�> �_5�^�8
����@����@O�/0 \���|`p;0�,�/����>�;�@,��@C�p	��(�X@o`0�r�\ ( ��`*0��� �+�W��@��9P��~�탡��K�v@  *�� �c�	�$`2p0��,���J`3�9��8D8���K�@7@�'p0���b�`&��X�� o ���6�k`p�8�.�$@���$�ƛCF�ȼEݠ�@K�j`mR��fa>��^��߱0����/�j��������:pnԟ�2W ��Ȱ!l�P��������Pͫ�B�]�굻B)@�>�&�NM(�$�O_�+��4�5��!����q��oB5�q|wM��S��;T�uw(y���	U�@)/��I@<���x�7P�0��K���Ԇꀲi�������,G���
U���\�+TS�����<��ŏ�	��B\�ݡ:����PEzM���oB�;p��A9�pM������;kBex��R�c_��f��܁P%��K�P���Bq(G5�;�`w(i�7�Jjk����Ն*��cx q�kC��@�+Tvʑ�{|����+T��7T�zo���}�P�ҥ��8��C�	����ȣ+�䋨�ƨg<_P
T#}
�\�,�eMʎ#_�O�˨�L<�k����P)�"��겮}m��]��Q�_�~<?O�v�뼠*��3ՠl_�~HW��{�({��x�Z�q/ʼ60������{�Ѩ�#�����P��( ,��G�"��s���Q_ȯ�	�-ڱ�A<��q�ȧ�������g�	�!�2c(�y���8��+p�:�\���ր6*�V�������Y��_�M��F�1h��]^�����l��S��ǠY�u9ڱ�q[����h�:�-�slĿ�/��8�e!���{I��X���,}yI�H?�D�ǹ��&�U����ܜ��7������v���0���E���"c�%c�G^j5�exu�S@���lX%9�&�3��+H�v�.';/���tU2�&�wt�PB��Wߛ;�j+ܹC�dl}���_���_V��rKy��ݺ�8�:��ŗ�;��%��6���O��,Ȃ�G�_۔�%��N�8�J��_A2&��ߒ��|���ڮ���<a���9��셼 �w����� �DtD�c�,��z�qak�lނ��u���A׷A4�"\�����f�O�W]�~� ^��_�3d���A_�������[w�jȏ��{�	dC��`��x�{qM����Pr����l�R�2	�E7i�_��<RL�H<�#��;�dy���|��Kr���������)�LD�d,���M��~�]
{#b��v,�:�6=jQTG��p�<���8E'Ȧ�M�>�?w�ϫ��0t	P� ���o<$�Y�5�S�����C�BFC/�>�[�$�
�h���`_:��;��M�]�+�y�}�]��U�����6@�a_6����wC��P1re/;�/T�6�
�O��U7�*�y4�*�>~3�������q�<�ˠ��!�7"=M���s�͇>*�~v�(��A��O�Kh�<����y���aNn����=�y��z������փ4��%��T��o'��V�&2�0qW2L�����S�l�vFb�`~:��܍\�a��3����g`:2eL� �b�0s���<Faff>�"��1�3S���blf��~�+���]�{�¸��6���`��U�o��}�i�5��?"�/�-̯�t�(�$ĳ�v,��d�0�V��e\6��p/6�$����lk������3��O�3�k����Y�%��\�A�a��\Ø�p�#�g��Y�����Vn6��+c�sL�:n�w/s�����+e~E�c�|�7���&r�o�7�O�v��V�G2o�L�j�!F4�X׳�{q=� Қ����4fQ�t��5��f^t�6�"�7�~_����l�g ����6�صm�����aַ�d��L�7#��_�)a�c��$�P����6��om
��8߱��K�QL׶��m&�mtܝm	�r��KHb�+�	3&q36q��8���DNHLe&&c�S���!L�S���L淉�#���b��>Ŵh��i(-cܛ�1�m�0S�1�3��eW2e�+��3��1mO4��l��x�4"q��
2��H�@�$��&}�`�����O> ������)�J�����Kť�J�ҵ˺��G/~sk��][�l��lk���ε;{�Z���ݗ�p�O���'��(=qǉ�O��Xx��Ϝx�D�'�=QubӉ��N�;q��'~=q�ı���6r�u��l�����D�2�C�Z"�f	��C�q`�eH%�Ұ�$j��Y}�}�[.$��	א0���Htt�݌���nN����|1�e-H�-[҂4KlI��-	S	�\J���D-���G.E����[�K+[��&1+�~;0"����nN<�XOU"�	�(iK.-�=����ߞ49ڞD%w ���G��	SבD�H�V���	�Չ�3�*`?���I G��3�tF:��-8��|}��Zu�����D�Q�%"�D\��v0��DwG��	��
�'\�{_A�7_��\# ^D�H�T`��z�>ZB��K8/㼌�� ZA��x�*�S���5�$�$��	3B'��:��`��jy$�U���ę$��$�!��-҆�I�j�\��!(.i��FG]r�$MW$�Ȅh��+f�@��xC� �'ڬ'��C�H���$6i�#�����~$asGn�u��7�DT�"l��Q�ד˫G>�~�H'�f�Ҡ4�4�������"�+�6~<iW2�D��e���rYi�'�D��Hdy4�KW�˳'�����iI��y���#M��Iġ|��<[HZ&��Q7��]e��&��B��2�pE�ꩠɩ(E)�\~;��$�A.)���M��?����l�@��7b�,Ax�X�����P���Vw���"�=��e�� �?��R�/$�]�z{�D�YE�u��gʻ
4���%2����H����ܵ�#�p��$-�+I��J�n�$ܑJ�g�E�R��ۄMz�Ďx��iC�H��U�I|�F�)a���f�!�tFO�ͲGb9e>�����(]����,d�R��"��.g�@b93����O�,y�m\�$���&��Y�f1;	{a���g)˓��K7?Ų%�؆K��L��YVx���f�O��!����z�ew G�A�Y���Z���g�f=s!�c�O �8��T�)9�1KqqU�9���������J�r�W�.J9���ǐ�w����>�E:�]��Ҝ��Op{Np�r|��o�'�o��wO���y&�όj�p{�9ޞ���٦	</$�\M������w��$�I��$aߓoR��d���d�'���7�܇���/\1��+�'����#~!IQ�Hr�KK����~Q�ɀ(��.������-�}}�h?:�Y4H�b+_�J$�Q���Q�Jߊj�᭨F��Q��ߎj��!ʮ�յ����5�**�l�b�6F�%��"+7G�ٱ9�)�0�C�Q->�j\�QT�TG1�㨗�?���|�-Q<��"ikT�C�E]��s��"��$Fz)1�oBzJ&���A�{�G��$�~?�ɭ�sG�z{�܉=�o�NO��m���ӻO�>=��[�>gn����{nK��7�IW��<$��mg�&b�����;���yܦ�l��3/;�9��.;W�����pg-�?��T�N�r�����3�W�_y�2��aK��`h�8�������������y�J�D*�?%/�_���Ne{1�$3�.��}L��_�E_�dd�dx�
	̈́�16�<õޥޕ��&Y%�$7o�(�|�ESa�x�Z���(����f��q�yy$?�{gC���/��o�t�}�卵���*�_@ׁ$�������^���Ϻe��8R~�6�W�Z���S��~�6TrZxJ8��KmhZ8��sm��p��Hm�,�>�ݡ��ʟjC���kCφ��?��PZ��Ն^	�+�����U��q�'}W���}T���ֆ�*��x�6�i�3"�y���@mhg��Ն�ԗmm�@}����O�Xm���4�>�~�@����П�<k����+�a.n��Y�;tI8\�����#�m�bw�k8\�twH
��vwH�S������v�z��u�w�
�2�&�It���	Y�V���i�����ޫ�S��oI#�w`u�׆R�>�Wn�]��_S��E���)8v�q��N;.����j��6�������:��[�����ĕ�7������w����?���.��#"���e����|i���{�W}{�O�k���:0������(�7��G3����ҫ�$���$���Ij��AR�>��[��8��Ҋ�}i>��6}t)��O$�C:�?�&�薜�{��AviȮ'!J��ޞ���/��|,x�l|����_���+i�v�so������w?���Ԅ����$���]I�C�]R��������q��$H���'��yK��ڛ�3q�MD�{fn.IK����
�&�M���fR�X��:W{ 4��v�IS��'����ʹ�Yf,	�2�!?>;�[e�[�[a�?�'>~���[\=���#�Cf�����
�3<W��\�V��&�(p�7�&� +7�}}ry����d�=�׌�)�}G�Ӓ���'M@�kK
H�N2�w�t�QH?D�+�ⶍ��Π>Lb��4�?��ܡ86��i^�<�h���wx��p��̒���Jo�oTNE[�W�T����Ӹ����ĉ��v?�����-U�t�}�?{v���ɺ[��z���Bo�E�T���iϸ߸����O��=N���f��?�S?���[T�7����<8%*��:��{���w�zze}��/p�6!�(	�M��&���a|b|����
��&e�:8��~'|��ytRxE���{����i�:vqnl�0�_�#�A#0Cn�M��t��C�<�3I�Ί��׻}*����K�C��6Eޠׄk%�_EH*������kA����)>!u��C�(��L�NE��~0tP���#��7/������W��{�o�|:�CBi,9
Tݎ�nhKH��T�@j��¨��@:��i׎����Ǥ�ž���&	��%��iI�a_F���m��{Х���J���)'!�8�4\��Lĵ@)��y ��C�
 ��a��F��x�+�|`.��	D�Kd�:`���`Z,с끙���.��]���������6ӑ?P,� �wǒ+�a�4`��h3#���ǀ�����%��"�a`p���X�� <|/���7�?mJM�IC��sc҄\D��f�9��� -�%�RҊ\FZ�q�I[Ҏ\�*�o�;��:�.�+I$� � �D���2ǌ�4֕����Hޑ+3&e���O;�=� +�w5��3-M��<W������LDǉ�#�%S��D��ޗ��I��WL� �ORo|�y��� �+�7D�|��s������E��s$�����T�:m���s���<Q�(�9S�vΧ�ꓞ��ק���K�v�o��!����&����A�I���ӄ�K� =���|����&��Iϣ��!�ib�W�s$��G��w�����y�S�S�S�qUA���s��8:l���;G2��dq�E�'x�#]nΘ�q@�:!L'���LE�s�i�9������������^����^�)σ�ꓞ���Oz���ІD�S=ϕ����I��W���Y�a�y�~8�yU~8��>��<�>��<��>%�%���K[JY��p�c�$wv,){�T\�"ةŒ�٧��W:'��m���G�����f`PG�ύ%-��� ҁ`0X�>� G��bI;�R��@0�� *�O�=��8���.0Lnf �%@��|�4����	�R�L��x
�6;��@�GbIS H��4`6�$�x��Ga�?��gG��0�J�;�{�y�"�`-����?���9��@+�=�h��R��� ���s�E�S�J`P	l� _�#��@�B����,��I��M�������b�������Yz��<��ҳ9+%w���t���KɆ�̸^�+�،ܡ�w����t��Mw���&��%��7?��*�>1qnJ3�oJ�2��8}����S�����g��N�Mͦ�& ��c������'3gq�J>�{,�qI��=�;�ӽ��a�����k�:̜�%����2�s�*_��X�*י=ӥ*!�ؿ8�$װg�Y��=���u�?�ZǞ�l��g��J
�3\��;�3���ɞ�w�Y������S�cO��J�gOw��{�+y�=�#�+�I���5����]�N���:$%U���1�oф����J"�3���F�)?�s'=���i�\I+�L�ݸ�ytȝ��(��X�w<�O�_o�Nz�%{�3�����_���G�5�=���]26˛������>�Y]Œ�|*u�8�[φ$�O�-��LMR2�O-�����z�oKF�y�%i��hI:�W_�����6(E�-KJ�ӿ�r6���-�x�?�w��S�m���	���U�SD�*t�(��<@�2�AN���$m��Z�ɠ,<�g��S�_ڥ��G�7Ŀ�a��P#H��t�>������L�j�K_Ai
!K��H_6-\��ٴb��ȭ\�M9������Z���A�⼡�m��A6p�X��9����l�Q�c���R��&��ƅ����y��=ݗ�_�q�N��7�0#7?;�������	�|���&�� �����R�i�~�#�>7Q��m���XH���9�Y$�G�y�]�{#?� �0�����}��������i87k"�(�&Ҥ~IyZE�7������3�nEȟ�T�O�|h����)Gh���O��C� K��tj!�&N[P�?]���{ȩ������wj�[���̿���[ˊ��V��⃡���m�{;�GH{��˄v�`a��)< ��^�X� Jb�*�Fq����������W��HM���$]%�&͐ޔ:+��D���U�*�Vm��RE�J�P��>�.U�S�R?SY-Nk�uӮ�fh�jOj�h_jǴ��D�f�N}��H_�W�k������H��1͘m�?-����wq���s���������l`5��Y],�J�2��Y�S֛֫�6�����m���*�]���ng�8m����i��ҩr�9_;?9�bw���������N	�\\���������C�B[a��j�q�xPܡ�֯73�k��d��]�Ղ��;���t�T��BKa��XxIx]xG�B�^�E�(����H����H�5�Z�V�Q�-��j�������i�}��]߯�4��ƵF�1Ѹɸ͘n<`�7�0�3^46��@���?�f����lg&���Af�9ռ˜i>h�2���VC�Yg���j��ҭۭ�V�5��;����+�a��ʽ�}��IG�%����)�&�'D�W��F�R)^)7UEUǨ/�5h�Jm�6C��wn�7���.q׹������ۂ����Z!����B���t����g�h'�I:u�M�ר��Ro)K��zG�F��;Ƚ嶊�l���v.u�+	��)HK�g�5J���L��F�� �i9�9�;�k�;���tG���e�#��A�����_*� �~�Kq�8\�[:!u�_���-�z�5�+�R�W_S�R-�zm����w��֟ӛ��������%t��2BhӅ��B+��H�K1rc�+�W�B���q܈�bm�vX��}nL0���!H����O\-~/I�I˥��*I��eR��.�׺j�fi������*m�vD�է�_����A�����c�8��v�!��$c�1"�l�`�7�7��_�5�A������K�K�����l���g�X�X���[U���N�u����݊�[آm��S�a�(;�ζ'ط�w۳���R��{=��jB�D~��]��a�5�#�1�x��!��R�Y��u�mc����8d�h�n0��@�@B���p��S��"���%[���Zì�)�]�lk���Zb��VY��'�n��G먥۷���P�'�Am���/��6�g!����K���g�sЉuۺ���h%ŝ�>�>�uI��^�ς.�k/j��}���4�Wo�8QG]r����֜f=m����@�R��a���a��ٯڗ:�&�ʖ8���.(<*�+8boq�x�8V�'�7�����Y��R�%�5q�X-nw����%5��I��˥�R� �QZEƈ�"�b3y�|��T�T�Mm��0�����ƛ�y��X<�W�֮�>Ѿ�z���7����o�$�@`�I˟�x��_�������}����������X���<�$ts�Ya�4~���Zh'@��t6:5��&���ָ|�p�p����Y�(I�+��͑^�vHM�Dy�\!�--7QXs���}0�D�#Z_�i��jL5>3��͇M�ϐT*k�^��H�K}H-��yM{_ߧ��_f�7��T<ռ��+��Q�z+˴��Z1����Gs,��;88*�����s2�e~ݾ,wҞӾ	@qV�����2�GF�UnIp&x�[���/��$^��g��B��/)W�۝���p���=�B�g�1}�
��=*��_�+/��h#���V��c�&n�*�Qw��?X�|5�F���� �d�,���B{���#� ] �)�!�,��L� u�������o�����RmZ���B���A�~
m�W�^?���PS���dd7�+�4fs�e�2V�ی��~����<i�
����jn��XXx%P�E�
|8��Ff����L5G�Y�D�&�Լǜm.0���A��an51c�&���V7K���@WCK���P۳����؍�fv'���B�E��hO�g�����e�5U�{������4uZ;	�����('˹�y�Ug=Zm�S��s.w%�v�vG��n�{�}�����������ֺߺu�ont������M���i�9�E�e���h�?���!�h�&B'���Wi�M��h�%����a�'!���{*E�K������'��o��Ú��=��6Jj!��%M
¾/}ͷҼ�!5���&D)���ꥐ��Тa�����@;S1e�ʜm/�q��Mv�`��'�gH��>�j� �]O)Uj"��'���]�������lP�P�C�L����?���x#�V�=PiI�6������s̡+Y�u�g
/H+�7�z��D]��x��$uzc��g�V�����>b7^�����LVX(]-�AS�S]5v�E�eZ�fjc�\�Fm�����>��8x�|�N�l��A���
���p)��w�	�2�A����jЫ�:01�8�=����aK ��ꤸ%�6w������d�O�Z��^Z&��T������M�a�9X5U�.�����_�V�4��Q���k�iE�[���b���^�V�����W�����YOa�0��ja���N�+.���aW��5b���/R�z��6� 1K|])=/}"}'u�%ٔ�))JG�E퀶Con�ظ p���/8���nr_t�p7��{�>�X�Oy)��]l��p�p�p����� ��ě�Mֈ(��PZ -�ƪ��o����U\T�?w5[��~��V�#C��`U[�a<iﴇ:��n����W<y�z������l��<q����S�,o�)ߠlVڪ��a��V���Kk���@JdZY��/ٛ`�!�Jֳ�*����u��j��I�̼�ޫ�?�T�,})��YӲ���G���|z�Mx��b���
��^3�8��'D�@l/v��'�q�|����N��.֒��F�1�h���� I�C`�Y���z6�d��4�hwq�8��7y}?��B��8��R4�����p�I���0e*8{����E;�]����օ6�u/�Au_C?e����:�<��I 4��h�[TM;��o���X���M���|��
-A�Aq����;"6v1zp��Q���ܦ|�|���t@�ߠ�F���z��V�M��k�!D�=O�\?�1�=1�x�dA��ǁ�f'��Z�P�����n^_`�;�}�h=9��J��O���,|F��!��%rP�C~	��[����e���J����;�~�~�E��>l�H�4YC+�����|:����l���+����n��]�j%O)�zBo���\Ȳ��x�ki��:�nO�I>�����yO8*tm�e��*�1Vj.u��"5���Ż����>�=��J9o1W�Aڧ^�E�����i�+A7��k���װmI�@��=������Z������u�Kb61/FON���V�#А_��%V�g��.������ �f�З�n=h-F�nB�b�u�����v�f��S�k�L�&{2l�G�E����oڛ�3ی�4v.�Δ�vW:�8���'���Ր�/��f'oN��~,�|�.�9m�2Γi�BA��*��.�(�,�T:ؗ�����mT!�)�s��h*�!p�ЈI��z5N��֚n	ԙ}�r�������,H*|>�*��������m�iDǬ6�?�ݪ�H�O[�4Z��{�g�wpŅ�EVK�#z8�[?X�v�}�-��߾ھΫ�Yv%4�n��n�tsz8ׂ��:˜U��7Xd7�C�5���?�	{@M!�wJ?C[? ��S�e�rL�@�����>S}D]���~�P�T[hm�Y�ic��6E�W{T+�j?h�h��z�2]���[�[���@���c���y�Y�'���laN\ �'���E(	�ō��H���q�WO߈�t��]n��������"񼧛�`��.�!핮�;*z��j��G���M"�^�&MZ&���8t���彶XG�B���m!Δ�Ux����ߡ�=��!�ޓ?U*����7�
���"y z�S�?���$p�� ��˝c�4�Z�}���Muا�C�y�Z+�u��w���sre���Յ���(�[@	�dBx�Rȩ�f<Z{��������W��i���?^*8��h}Fxǅj]`�4$.���I�0e)lE6H�#�r��t�X�
6�O�xYs>�����@Os I�;�����~[���u���<7&8����i�K��~ZO�~��O���kd���o�Ѵ����`G� �s�L�0���*�C}��V���HvOp�����y=��t]�"��
݄dX!��|�lM�.�*��X��m���I*�����m�d�T�VV��z�q��(|P�h��-x:��AB���.Hj��U1J�-/�i���Ǆ��֯�~o�Z��L��Js�u)���Ez��-��=���J���O�7�EO�G��H'���b�k��ٝ`[Fz�wLئ>�m�Z�:�`�}I���`�,���Z�]�g�E]�h��dk�����Q�$�v�F��tW��7�JǕ���}���1�}�5���`��t�<��7���g�N���<�Ͽ'}��:�V�u)�
���(�*��O�V���)��K�5j��-�烵�+�?-�t[懟��/ҳ�O?c@���U�k�u�E-���=�U����>��
��k�+�DK�I[�����_k�σ�����(z����^cf��l�H�N*���U��yy�Zk��G@�͆�}l�A����Dz���� ,�j����}�����1�y�"6��ӿtH\�g�_(4�4�%?~�WJalU~T2�bȦf� ��.��\�XcJ��'��c���h�4x�K�<[�!�a}�q�x���������^F�q���Xi�j���>���jk���5���v���)q_p��
�Ey2���	C�|���!�w������� u�:]�_]�V�հU�PGi[ ׷�y��M�?)��P[^�K�R�@��#�#=$u?�ߗY%Vi�$+�q�t�~e9���j�&X���>�P�X���վ�.���?��M��{�e��R�Zk����ϰk_�h6����r��_�T�h�G���۵8}��
�sI~�G�͍��'�g̮�`�����p>t��a����A�����n3g�e�w�p������=OJ�Q����B�P*�v	���h����jo�M���G�6�efB�=kwvL�^S�k�c��ߔGy���n�n1^J�b�@�+p� =�H0�W��w؃�Li��o�ta�p��T\!~*�JzPy�nK=U�V�Ћ�K�Y����l1��Ak����η?�Ӡo�|Ơ���VzX�G��>w�A���G�stј�I���z8w;�:ۜ>��Ӄ�F�Γ�QR��ᨨ�%_&��4e��2P]���1��Z�'Pf{s2l��g���ӯ�ׄM���(���fik5J��B�\h&���R�ں˞�|�:�������fF'X�w芚��%q��r�* [�X��mо�~3�.5I\�w�nb�Z f���x�Xm�e���Ӽ��i�g��+���� K��G{<|�86�[�v��K�H�t�����՟��鍍�E��CX�	�I��2o�.�5v������MFy���0@�*�!~+�$v��I_IM��r!�핑J�2B}@�\e����z���hZ؄Z"���mȷ��^��������0�㇞��+f�UDuHJ�'�,������hO�r�,�}ԕ�>�Y���/�jeZX$?ړeQ���h��j��Z{�I���.P ���,�?��ʒr�2O�����6+�β�@��"WvG����Ö��K[%K�)oU[��&�~� ۥCR#y��2�nS�4E�����H�S9m�6F{J�R�B\�I���1�U�A#>0"p}���H:���T���Y��C���y�6w���L�������d��B�0Y8&�)t����b7����T-o�c�x�TV��r�+P�Wk��e�}�s�Eh�;��SF%��
LE;����%p����+P����l7ǘ;a�GY�YWX��������VkX�����=�+�^�s�� 7��ug�����s��G�| ���P�����d�:�w	�
��O���OBQG�����b��J�%KJ����3N�_�'�I9���������@q�q���N��O�/��ͽ��&�~D3����5�d+�m͵�VX/Y�-��[D؍�k =�_�?�c��wr*�7�O�}�K4A��v����w��;����z�vw��O�G9)xW��3���>s��|�Q�R�J�Y�n����	{�#��v�$&C�="�Dou���xD<&���v�tɆ�K���!� �(�"͔��*�������Q�O��|��)��y�d����/����#��b�2������bh��ʃ�ἠ��lTh�f6�6��_Ԇ�E����j��d�N�k@�l��w����	�7����o��r���>8(x]�08�t����%BG��Y��h���Or��V��O_�/A������ �v�)�{����������t��	���o?۩v��n�;&�b���N�D�.��bS���#>&}4m�J��?��I_�otX�u)7��˭��Ki�+�������8y�<I���~y�3O�+����w��m���^�w�@^E*��Jk���]�W�R�)���'*��)�Ɵ�,R�RV*/+�w�ѣ�Z٫V~Q�T"Նjs���Q�j��4H����1Q��N�yh�� �^Vף���M�ZݫF��FjM�,�H�G{N{Y�Dkg��Φ�0Ɠe�*]m����j����a�t�8]����}�!�X�C.S�s�g(Br�X*Ng���2����rq��Z�B\-�׉���J�,V�[�v�����Cb���x\���ˉ�;���"�ʣ�t9[Ε���4�ɳ�2y��P^"W���J�J���C:�Ao�tz\�h%Ni���|JPE1�$ϚJQF(��L%[�W��ɠ��,e�2��J�
X��J�R����FٯR�(G��j5Nm��R۫	��*��&��`索#�t5��|�D��NSg�e��?�!�W��a�W��Ͱ��;�=�~�j���h�h�5����Z�����i��4m�V���jK�
m����Eۮ���=��ף�z��To������z8L�=E�����L=�q�^����R}�>C����RY���+�*�Z߮70Z�a��J�i�Bc9$�fc�Qg4�;���(�*�K��j��g&��9�a曓ѷ)7ט��~�X �<S�\��Z[j;zRǭh;�N���;�.�ͷ+�u���>j�N+pj�3��t��ؚk��;�#q[��!�������2w9,�͐�Gܣ�q�E�U0>h�����`&����������`Eps�:�%�'x��^����J!Iȅ$-���WB���b��I��.E��������HqRS���J��dM�a�(� )[��n�Ρ��P*��H˥����5�:�R:��/G��8���Bn%S�O ��ڷ�$��x0��L��=>��q���x�P~X��c��Z^����3�=���q�~�?�xB�#<.i��I{�S�Wl�[�y���qL��3�הx|3��2�wzܳ���Uz<������8����7E{����x�(�,�����u�Ty\����sy�s����@��x�����l-	\�O NJ�F��ҵLpT���*�N��5��9w����k+<[.���[�m֪=nۡ�@{������֓�d�z#)�Y�����rp�r�c��Z_��_n gnonw��k�=�~����#�Q��Nވ�*��M2��~� #�;��4��\#�W�1�(G�0fe�c�z����o1�;�p�~�8��q�8;�D�M-��[��2OK;�H��<H�=9*��dr���@I`2dĴ����@Y`N`~X^,���:���2��cs�v���ȑ=���%u�#����b�f�� �����leƛ�!cMr�0m3	��~�8)f*��(3}�l3��,�*5��3�Yf��|s!$�s��¬0S�{e��fφDʇ�_bM�J�i�k�Ufͱ�CJ�[K`��*���k�����lUæ�n����¹k����(���������5�������lWCoG���}?zu�H��6qx'�i��9M����N{��DGpX�6�u2�j�'��r�!���\��"�ę�:� �g9e���N���Y�^ᬆl_�T:�*g3��g;$}����+�2��sr�w��n����-��&�����A���0�MA�`��t7�͆��w��w�[
]1Ý}1ǝ�.t��%���@�����-6�`��[A� ��������R��(�?bl>��qFS��VF���H0��>ǘ=^���rc�Q����L�/#c����>�D��D��3<�/ٳ�R<�o�g�e{�_�g��z��,�����i�2L�m(��n��]��ָ��Jw�[����l�[��q���ܺ�=F�|0:� l�m����`bP*Av�_�!pZQE���"��QQ���`>��@ �@ D�@D *""**"�@ ���"�����2D��0��}{����F!�~������/o��nfz��;skۭu��x�n��r���~s1
f:O|7��D2���n��w$�?M�އV{WM�h؝k���iT��]�U�o0�#xkn���$��aN@1h��h�eڞ@�sh��B�qh6�^A�5h�M~����{��`>@g1�+]��*tԂ~>�2�N�G��\�U_�/I��c	�tһߙ�G�m�9��$ݦ,m�Z��Kҽ����bU�-��i-�����`]�-W�4<������U���ıN�i^9�S�����=(9*��,��$A̗���d$+9�KA�r�.I$]����F`ꖴ���PF2�מy�������H<�Y�i^Z�_kI�Zњ��F��]t�ׁu�c��Tg�C�I���7L�����>�W���b^�r�k߸��k�x�G��yO��x%��yj��>Sps�S�3�������~�n��3������y`:`�_�_�@���z�3�ߥ�e̂90��w�=���e쌜q3jzZ:Z��$�,`���J}�~��C�O�����I���j�N�N؝�F�:�3��n�=_� PK
    �\Itg�1�	  @ /  org/sqlite/native/Windows/x86_64/sqlitejdbc.dll   @     �	     Խ}|T��0~�f7��w		0�����P�&w�.l4����U�)�T)ޅ��lzw5�۵��o������W�jx���@^@4	�u��!��}Ι���`�|���_>���;sf��̙3�93�bQ#��0��#�Y��?�����?l��a̻���ֳΝ��/y��e�����_��c�=.�?�H�r�c��>�/�9/�Ǐ?�Ȕ�����J;�<�L�q�]�r{�)�d�t#�%&���e��7̘����uo�3��uf��_3H�&���'>�޵�eL ��<0"����3Gg'��3�B�蔵�~��7=��e��)�#5���&��}|>S�������^q�2�&#dc�OYN�!�ҷB��!p�)�(i#��qB�<}\�mJ��4+���n��CO<�ύ�ؘ�˶Ս�=B�#}}�dB8<���(�#cc��@x�8���� ^� ���8��"-%����V��:��W1t�a��sڐz�.�������700ɂ��&FTZD%�����E�0iND&C���$��yU����[���n����Ͽ랻I��nQ��TZ]O���s[c�{�k��c�ů�z!b#��+ro�B��~Q�qӊf3�i47��lBm����!o~ �T�G�_�yL �a,��,0Q,	j��>��y�%Q��#��_����ŏ�M~k�@��U�n��c%��+��[��3�!��b��C2N�9d���+*,�����P�|�p�N-���F\�X��-��޷LX���Pz7"���H�l���2vp;��n�_ї���ۗ5�6�(
!��&&�kլU�����xJ��1�-�8�U�OE뙕#D5�?��N�Zq0�P��f�v'�vx�V{l3iO��ݙ1����{(x)T��#��
���kLP@��2�B' ��Z B����QO!R�G�.��M��7�-�
�P9�0|���8������L��*�O��yJc��6��D�+D�Z��	����2E_�֠p1�����	��MQ��t��W�Q\!�2�M0�@����Y�7��gFS�É/G/D"���Q���X���yf'F�-Z�x(���@�h!��B�@L|�a�����L�~
�Qҹ�#vK��Dx�[йF�R���h���/(gA�S

�YPp�撑q��*���"f�Y��.(mN�pK)2����F�@TSx在��r��A6F(�ȑ(=���gxr��q���@Tsۧg0�F#��l��𿪹��h��� ������USDe �յK`ٌ4�`-S�Nǩ����@�Ր#=0����R�ᛍ�~��ߐ��c�UG��R'|��Ķ�"І6����9"�i7n$|�V�խXA�.�@|�O��h`����@�q����F���Mo�9@z1Pj�QB$"�eMX����	���
k�ǼUQ.2���y|Y�c��b|ܚA�A0�K$p'6���m��UD��4���BP�3��?�,D�Ԣ�&Q���Q~�-�����ҟ��_$�S����b+R	r�=�Q�Чm@�d~��?�e+��>���Y`��E�|�w6R�!癪#�t�$����</b�q���}�����L�BR�,�qYJ,.����iP����W��D�������k��VA�����wU����� J� �4eHD�+�U�#��F ���y�6 ���TQ9��!F��AGo�:h���D�$�̄^��a=��`�J�"�6����b��HѠ����v�ǉI炫:X�]���� � �k���eݾ���u�,�ܢ���%�7�0"r�̧���AF�!��@ �.4�� ���ӈ�t��% Eʯ��Ps��u��˚�~�����	���HB����v�	]{)��͗��E�;Ց�Y��H��I��"�?+�e��c�/7���H5�����M���Q�3��̐�|�5j��D��<���6����ΩA¨�vH�@�9{3R�/�BA~�ǰ��UDTG��[�P*�O�˗{�=�ߪ&�o8J�+SLHK���-��V6�Q��c����X`��ŵ��F���6����)GE.�&͇c�Y�6��Ak�6h�y��V�7���O8(m��l@ۦI=����q����{�߿G�95q�1��ͩ�0=�����MT�=$��5����]�R��F Ѕ��TT�����*�G�$�Q B�H�ޢ���ܔ�;��H�Ɓx�D����J�Cg<�.i�{�&6ܔ��e�~9Y�@l��_��w�񢼜�l��~�!&:}}�����bK�\���H��_�~q#f�����d1(������l�4��w���`����6a��*��!]��^����t�=~�|,EcM:k	���ձ�:]��e3�Bu���w�o�T����A�&�@WK͚w袻��N��`s������� �*�0�"�����#� ��A�u	 [��Da+� �˂D�TA!�Y�s�#Q�x�2m���و���N�6�Y!`z)%Ô�	��6!�Ŗ���� *�K��&���F�HP��>m@o4�紐�N��S͈��B��}�<-m4鄎� �,A><Bqze-�酵���!8} Q�u��|6�M��&
g��AT�Q� }]���u�~t/��O�>��@�4��,��8�m^Tv��AEckthOǆ��#��a~=�������'��kW]�S�mD��(۽GA-(qO���#ACJ��� ��2Y���@��E�h��*�.C} ���.�r����K�\*�K�`"z�\Dg5�������k�e�~}.�����)7��4�l<9y�i���� u-j-�5g(�U�1��6;H~B0=ߙ�CQ]C�,��O�|����|Dz��L�~� �H�	�jr�S	�~a`ߍBj�������L�{{ɠ�i�wAَQw-G�4�����A�-�RF�y��2���A/�"EJ��`W�%�ש>���0S��_W�C��[G���$T�_+�%j�J�/��O����Dz�uD�����!no��Ų�4�+��&rK�	��&����A(
�"�n�&��J3�gto*�TTm%�bA[�8�D�yG��O�A���8/au��w"�U�E80���L�wՍ����6���˒���u�^4E@|���ߝ�w�Os���s=߽�����:�B�>�z�)m�b��B���9'0�����Ybc�6�+�e�O����H��6��T��(@ۆv?�6i�1觨����F�7��4(�D�-�O��W28������sE?ί����(>��1�z�Ci	�5��z�IL2�LZT����2�$���g�@�ot�'���6�%��.��o�)��>$-������Al�]g�/�����Ů���Ft�A7c#A�vq"҄����_�S(��Q|�W��'��}�o5W���ݝYo��r���I�;�w�qN�ٮ�C��;�ǖ�r\4~t��)�������&S�6���X���8���h�;L���t�H�/�J�V�&�+��q�E�f& ��f����td�_���>��gһ}ob��{��o�w_��w���&HK�ѥ��Kw��06?��?���
��8<?>�?�g_e�ߠ�/w�@�fC'vW����s&�'9�՚�i�;�QK��	(R��cAc��0��YF��F��H�K0"�4^w*V.M��#I�#FǸ��|�`۝����D잣Nߌߟ�D���=���NN��~'g�	�~,�7�	jQ�A* b
�J��ة<�|�[����u�������oA{�_� �����=Hם12�������� z�����w|����c��������by{OCy�Pgn�����Q`N\UH��P~�W���]�8�P}���ʺ���I�1{2�s[�H�9�ITh��1#$A�M2"'O�eԆ�2�D�[̣�̄+�e�&X���H�}�O6a�w]w�o��!���O�Q�/w�D�)�h!��?Y�G��3a9n���d��FS�
W�D���υ``��
�ڕ/��c��S����uP[�p����XN��&j���y�e��ΓZ���S�7����+�r+[�vF�	
�'8ϯ ƅ����O�<��m2p>�Qև�h�R9��#��p�����%�p,�*�pV��ġ�Z ����-������Y�0�%pMP|(�X�jb�L� ��&i�h��G�@���G�wZ��$��q��7���yS'aj�.���i�f�z��S���1�H����}(*�bu�n�����,-��s��.���q4����P��H��N�����|v���'�d�/�?W�%d�����K$Ŷ�"����1k�ܖ�]F�u']I�kl�<�D�~!n����9�&UpT�!�U{e�ƇjD<�!���
�E�ę�
��w���-�k����]:"lCÁ%;��&}��GbM�k�Ek��op��'Xi�L
>�Z
�]op��h�NԒ�c�|.m�0�gX>j��U}�����ہN��º]�A�v�����ҭi�9j���O��fUf��3 ^1�!{K�߅�A�CX$��Fь��Z�(�}yNt!�>��]3��ĖV~*��+��媎�W�q����!���4���%��$�+��+p�@�H�&�1rD�}����ι&�ۍ��� r�Z�U�u!T1OTr��Q�:Bc@��:D��>����>ie�6Q�aa�k0�I�Z�!�I�i<3��M_�_��k��#�^���~_o$����;�����K��W�u'��d^Ԁ�!͏�V�Id��ܫ�ʙ�!��7�#�� �oq��~�<�2+��R#�7�iJڡ���m$c�Z��S1����sX�bxqLFB���gu�HUv"�P�	Sg,%��30h3\?&#6*�˟� �RĲ;��.�Έ&�&�cΏ&m��AT.H_�`��m�^���5T�D/j6פs��@�cg�nڊ� ��ƥ3����o �\����2�>.���k�(7�P�{n���J���BG3@jT�D�[���bF�Qi�?��G"��>�q�It?R��#��.A�FL�Iؒ���Vz�k�Īn�/3��wX;���s=ݮ��=��:�O�n�6����g��9슣�F?>��n^nv�v�r���c,����e�[:FX��L���W�s�>��]�}K�����������p��BCf6��b�TTu*�3���l{�~�3K��f]Ä��"���Ӫ�V}6���_#��H�-�����W�6���c���s�C\��K�Ӭ-���,?�{;�%~il�F�i.t������i�<���5� ̅r\{�$4�~���_`G��v�pM�A6Y�>@�Kp���SR�ڽ~�g���`��s��p�o,d�b˹����%�Y��pq�:JJu��A��Δ�#��-��-^M?d���4`���]Թ���Q}<Y~.���X��-����A
����(�u�V�X��v��t�+�-�0���t/1.Xw�~ �0@��n9(X��4�"Ͻ��ˇ���C���� fa=�ĭвq��0�t���>����9�v�����!�'�J�Z֧gX�*�
G��/�ka��ɻ/L�<}����D~KZ1AOދ9o#JmU���!�O?J<{(<��"�%d�@�:��01�N��]��&|z���{��\>{�3*���y:8�{:j�]G��䋬����Tsޯ�۫+������ӧw�'�
�)��_{ܩ�ų�x�\�Y��<�8߳��+���}��o|f�y��1�?�?60�Z��h�T@кW�������a��N��t(�����<�#��C7-�|1rhi���T@�}���y�H�C��Y; �=L?����Ϟ:gQ�C�$9�����bQ����Bd�K��@h8
B�q�����<!h���8t�c�v��f�F�GE\�d�@+����+�tK����F;���l_���G���LE��
��	b��2���I�kވ4�D�#��hE� �z�j�[m,�e��2N�k�o���y�t�.e�-���λ�쪾�w�A'{
蜓�CTPĻ/�� Dzq"�W��LK�d��O��G��_��r0l���ѿ�F�}����~�Tsr%K�mR������p0/�J ��<w�Զo2C��XQ�)I�x�o*Z}!9���[����<���<�8�� ��ܾ�+��MxB©
(~�<^��9���[�#Ta��~����G[����<X}�~R!Ͳ�	�?	�I��$�4n��>$SO`O����!��}��܋o7�;��@h酘?K�n~�}�]���i��]8O�3��tv<�4���U톜ᭂ�� S��
{�I��OIi�Ђ�A糜�XQ�q���(<��+a��`� +� -�B3 �>rΜ��Ȑ���:���Hx�9�?Hf������������w�F8�>���<�!����=��&����cȇ�)��I�7Rwv����$O��y�iH%��y~ɐ��r`�w� ��"�qY��P�5&�/�I!��7Н0�ڄ9���uX�C�"��N%2����P=�6�O$6��2�@q�p�D2��i�Ϲ�\P�v�dDf[��q���چ��ug
]���9a9����g�\ϸ
X�ʴ�"����tA���zv�Ou�ƽڊ���Y¶�z氶�����17^4�d�}����WV�7*��? l���Uާ�R�K',�����v�Q���ik�t���8:�����m���a�>��=K�I�!��}x��#>��u������yA�U7D�=�����&`T�@g>��Q?��̂d#�K��K ��g� �d��=�ǰ�}�P�m�n�``�`��[�g����2��vT�|D�t�v�a����/9���	Vޫ���>˧�v�=X�Hzb'�_�!&�bK_��B��=�����|7BU��]5�'Lf�#n��j�l�ꮘ���=_Q��W��/����{*�#(�&�]`��G��fQх^��ᡟ]�������	�lߋ CRZ� �_K�i�	}p�GH�8��'��~B�K$��ǀ
B�	a*Z��[���)����iJ�#�G�cFe���;���i"��]��&��l5/nᕀ�I���|�@���̓��:�.(������f�à�D��"�-���n�!�����ݮ�rO]�'M0�8���Ti�D�.�3L0���vM��n|�t�8�OjO�������H�a$���N*9����
��<?G��R���avS�*ەX_ 8\���M�)��@�S:b��@����}��q|�a,2AAi4c���_�J2�H�TZ�~R���ҡ�f��X/�L*M�q�*M��Z��^+�7�k�jy�Z^�c���:������=8��L�4[f3i�`~�8�5׃D[{�����WG���r{]��mF#_6ڳδ ��"��@�(
]a���K�/�K[�X�?�+�M���gŨ��.��ͅ��^�C��bd,WHnNǸ��@�/wbQ:#N����)�YgZP8Ǯ�[[H���H�߄;���	����	q�|��ѕh��{J��Ê���ob��5|9۰n���W�-��`�x�'���/=zp�?1����+=|-�/�4�Q�;�D�@�G��X�+�llAϊ؋��UzKw�߄��K�>�`R���,b$�����`��$ٟ�p_��	��h��,���7��DL$�����x(�e �hs��^9C3?�����WH��Д���/��@iR�p�w���P����Z���h��r*� ��l�����,}� ��w�V�V����)+�'xA������&s$w8�
���&��&��F-�m�������G�Vn�+�+�)��"�7CfE��e,:#�O[�K,��$m/��������ٴ��!�﹯PIk�{6��
�O-ڡ������S���A��UriG$����@�7q��ϔ����8�ae�v1p�6��1X 6��ey��@�X�]�Sv������/���Q�{\@!1;%Z[�=Ĉ�0�]>&�|��ϞR�<��0��+��0
�$�'�V7��2�@P�1��8���O��1�V' u*͊_P��f�G��Z�'�vk;����Z杂okdV:�����.Ai�4U�7Ew��m�Q���I`͂ ���_�a[�C@ܿz�6���q~�~bK"> @)|q_3+��V�,�ĩ�%��l��9�Bm�:5�
�/�xm���a��@Ou�ʜ�~Q�e�3���;���O2��EE�X�Dc��	�.*�����\�+T�<��A�^�b3����c�5�P�h�^m����X�� ��y���Bsqs��) RT{��
?�U�핗䱀����l��C6@C��|)_�v����_�.�!�jB���#�'��t��CJ'U�M����b�C!c�j}Pb��[���/&���%������7 �[W>Iy�P�I��ӥa����u�`��ɗ������JO��Q�4��JA-+�|�����VI��:�\�!Y��$&_�� �/�T L��y�w�~H�|QE��n	��V�T�
1�q�P �ͦ�����-��-d����O�򝪉dU���(_�'%ٓua�C��3�t\��-�r #�����Tmy��:�P� [(J�-LwؕY�x.�,��zAq��������7�/ϩ�V��)����#����g��3&����4�4��n�<��o-!�'3�S@U�q�-&�d�X E�6bZF��l�֬�Q�Z{j�+û.�?��g�A��DZ}�#�@���j�v�J��؈>4�D%5�Lv���}�AD��ȶr#�r3�9M��#ֱ,Qz_h$����h�x�	a�[`se�o����c���f\l�i��E�	[pJ'�nwv�Q`�tG�����k�(nF�,ҥ��d6#e���5Hz[��Z.>Ri����Z�G�Ӊ	d/��kJ��q��^x�r��G��n%��|K���I�;-�0뗦�n���V��&`$n�X���RW�U!a��|՝H�J�ܓB�\���������aAh�3�
X<�>S��sL+������ah����$1�D�#�m�k�KE ��)<�t�]1����.���F|��� ����Ш?�_w?�wI�߷�,e�!	)�t,����yh3�$��S���Qvu����P���j��v��u��\������k��/%OP*����/j��ݥt�AC4�?2 S~`i5!�gw�P�C�
���8)�r v{��}�/�ʕ�
{��K��ΐؕh��O��HY�MG�/S�߀�+�J�z���2�8 z��ݢr.�Hc�Z��������f�=�#+;*��f8��N��a�Z;|`��'�1�<`�C�7��؋>�c�F���ڈ��w�	E_A�|dD��P����WTu��;�/�/%�SJֽ7�b����^�\}�Q�vXg�H����	���SY)�LKc�:k��c��E��=���V�t���1���� �~ɻ�u��a\�ռ<k�M�7Z��Ǣo��u�����'U����r����Hª��V�i״4��F��d�sM:��nE�ӷ�(�ԅө?���cP��f�}8�� ���3�*���ٜ68��+�@m3�����9!p��@�9E�<�'� ^���\��c�3�YSa�*�'��gO	����se�0�O0�5��W��ڲ���K�E��2OGM�X��2���I֟_p1�&:U�M�4�ƪ/���;WTյ��G:Qɓe�gi/����$���y�BO�7����P�Q��@�+��@Xǃ"�=��4Z��_�5���[iUoEs�[�����w�N�U��u��t`'�E��>}ŝ�7k׊T��%��pf�?�!�ҍ
w�V|/��U�d
t 'tZ���Uڭ��VAŖn�A�k�x�������g�����Lg���m�p;�Չk����a�:���P�X�����3d�h��w*������vN�C�w�nGʜJM���ǼQ�:coF�+�&���C�H5�t���u��<n�~Y��2d�sV5�A��\��K��~�U��v����y�,	��×�؁�Z�/�.���&(�ӗ���W�<tv6���+�튑�
��j���OM�/��Z��+�RF������@���a��~����{��.!km��|�a<�9[ψo7�=o�'�_��^����j��0��c�U�{�S�i�>�RT�ѩ�i�spM>��0+�\2�7�7�~+b���|������+]����~���J��c�U���a�#�9F�j1� fihԿ#�kb��mi��<�Ԏ�,8l֞���
e
pM��8�O�:1�RS��qE2u��l@H� e�ܩd��� �#�iΜY@6 ��ܔ��:)��^�+6#5��[�Z�S�X��P5�f3�i� yX�X1�ʜ��~E:�+�F>�r�r�t��L(�Ҙ`�}���af+]wTe6���	�_���ǌZm�C1����*.���� 
��Z7�-'X��S��-���#����(�sL3����6�`��9)�����Z�:
L�E#.;9G2��hڎ�"A�6��KZ��r�)�i��գ���ۙ�� ��(�r�mb䞱�Wt��Ðq�6c\�ą��%!4w>n����OP�|��B�A����+����J��k�w&�7�>�j�lI��iܺ�B����U�LB�P�Mբ%j�&��H�槗	�N�Lro�ݚ#��a�E��8�@	A��E1ev~d��v�*$�L�7�#����"j+�/�:s�Н	�'�{������9(���Z��k� �:n���ݎ��>�_��҇].}��hH��kc�^.�J���?/�^�6�����ϑt���c�K�K�cH:_=���!���]{5��D���ksD�L������8���?#��+F�C�D��?�*��g��8R}�MH��M�*�����s/AE���<��uH���$��@�-��/@M�D�X{0)�7����#���n�
�^��AJkӿ�h�<Q���:����Z��v���8u�h��4`j�x�d���PgpK���t�?y�����o�Ū�5d&��=�J���0�\����6��x
�P��z�C8	m��E*+Ɂ(����x�\fA�;!f�-
��5j�=oh}O�z'Q�Z*�b'< ,��pP*���4�Z\
�g��+'S������N����I#�OB	��P��	gD��E:X 㧦1�W�V��W��%�Ѻ�z��׮T�/dʦa\�>�|X���KN�ZS:�����O�5\Y���?<~i8�d��'�[��.�t��X����G�P��G	���ݥ��c�o�DX��L�i��O�1@z��區q暄1���í (0��v�H�XX��K�f\0��.چ�c ��3{)�R�Fm��,�����S�O��_ �!����V���j����Ė�뎨�k�z���Q�9�3y�OT&P�x',V�
�F��2�P��^�"(� ��z�oe��I�5{9��$Iİ�SV�驵:%blCb�dp�_����f��s%}��4�.�D
�Y��j�ك�jv��D�2�d����	Q!��	k���B���Jϯ����Z�܏d?)����-�:O��oTF9�w3/Y�*-�D���1D����R)%m#�|��p�a��gS�2[Sb�Qʵ���P�'�Q��6��>�"���n!�p�� Uo�.�vK_��_9��*it鳴~�d�^��� �"���h�$�N�]��V��}ezVz#K�RV���,�(}�c������50;k�$�o��T7�\�]�?����*� �2'j�0��V�*���P�3+�K=�s-~X�ZJ_���6Lp|K����'I�>>�L�S<Z{q�����T��m��d.)���>��{+($N�!�I^� �J�L�_�u�_[U)��Z�;i�z���>C�kFx|E*�ε��eP2�<(a�+(+�h��?���Ӱ�f�+P���:��m�l��������z=���0�D�r�^@�<A3��@ݍ��=5�]�ʐEk�X�}>me6h�y����B�±��T�͖I(_��8���G�u�G�����t�2��Au,���6^�*8�s/�2e�P�ch~׆���Ĳ�i���2[Z�����Ҫ��G��'��T�	AyRLP��k�v���UW�4��;n��nj�w�IW��s7��&
$�^��yZ~�զ��
��F�&�({*��voG�l�q�|��/�ܝ��W1��|\@*�©��"���zg� r���C��]��6���ºI�$�7��9���l?H��-�_�e���&���՗���N��<D��+��N��pJ�m�t(Zk}�?�O���9�f�[:��#�Ns��`y�s��ed��Y3�����˱��#z4ό�mcl�+pX<�)0:�|�e�w���h�dSW�%L�H�8�a,�05D��l=/]#���W��}�)��I��x�x(V1O���W[�.��g�Lѷ�h�g�����0Y��R)�!g�6���r�V�	�?A%�I"�,�������<���}kj��WTn��br��\���G�!ie����*\uE	�p=0�dz"}$���<\��0���V�&2�Kdc�DM�]��2�����D��+�t����1����k�`	D�p���
`=�y0��^�<W�c�
X�<~�a���ōo�rk�4_�ԭ4�=�D�z�5���Ji����.9��<��t:��m��4״�qM��e%�:WS�m�A�V����>��o���ټ��4YT=Z��S3	�6��[OJ{C�K�A�°�S;�v�gUKX�9�_��eV~,ۘ�b�J����\"�/�@%�����y�ⱃ���{Y�'�FP�PD��!^��"k�����X9)���A����]����Oj��z��-m��M��ֶ�Y����(��ZM�o��|�=��HR)0��Ġ����O��!�+H��*B߃QA.��/(�<'/�G�h�t!G�C��s��O.ѱ�*�%�|z�b�}���8v6�9����qs5"����\!]�,�?�*�q@��]&��k���ו�&F�"���q��R]B�qDg 6�j(����~�aQ����)��/x#��Wj��w�^����EXƁ8:xn9��W����d�=��A�|p���^�	�s^�4}��<�(<��|��v���<|���qM6�}nˊ��?�ǁ	�]�&��NL[*�ѼcB��]�'c��i��c��.������~���g�ǓQ����B"/�\l�oa!]�ڻ:��ޘ`W>�vs���!־���X�����g��A$��}c}�-�j���i� �v��p��=�4�UuiA��%�|�C%AX��(���������VQ�V,��f�9��ݫ��-�J���voD:���J�>�DVj�^��|���VB�t	��w19CL�-��W��&5�;��x;\��PJg,AA�ݚ��j�"���A�Hq�2Y�O`�E�(���"4��F��G�0^kއ�S��a�&F鏊N�=��٪> (�� ����`�������/y��L�]���	�ַB���0��G�����P����jH&Gk+,ǣ�A��/�_<}��r(����"�E�6�ѣ�%rq�]�E�~�2X��e��3�K���]^>�:3Ky���Uq3H(��z��&�<[Ϻ��\-(US]�����nP?Q��i�X���t~��jf	�$?�\�*���#�גv�����_Ӌ�^-2ĉz̩|��)@F��b��5�.ht��@��UFx�JG�.�m�K_�*KW���n�']���-��Q��5�r�h�J�&�sM/��F��[��~7����H�����9P ��B�]�@9{��Νd����+�}0#b���2��R��5\���N�ۘ��G#�:b��<hY�9�m9�y^G.z�k��7��L���Y��_� ���!�ń�BYk�n�@O��Ng����#>W�š;�P�壘q�b$���z�J�2ЪWCn����
:���0�����:/	������k�@��
&��U�@���3(X;R*�N5*���^��$����q �lzh?�R�V.�*@{��?���Z��(��Q1}^���7/f{�MV����s����	�WoF6T��Z��B�B����eI) ��Cd����Wk���
��B'���>ȈA6�_�o>o��g%���j��}ˈ�z�n�~�`�2�~)X 6����x��6΃0��G���{��U�kn�>D&�a�󟚍<�z��Q�ۉ���n�/w@��tH.ak�|ȗt���
��f����j����Y�p�ߕ��Xs�����D��&�.�0�7�3���v���%n��%s$m������u~b'�I,(m�p~���]���*k֖�1 ��Ek��s��(�S�%�ۅ�O��r}f�'�S�rD�b�KP3�Civ =Vϴޛm~:}�oi�R�#� DB��ܺ�tD�­k���^�b�v���p�҃-5�?ĭӫ�EŌ��Z���PT\Z�of�ɥ�Dp/��y��=G�����ŉU-�XD�����[xkw��l7�v��:�Wg^����N�&�jӻN���>w�t�����V��6��$7ص���-�hle�
l�"�U1SC7�?���oQ$ѿv�c4!�{���,nb�Qk����>(�F�_ P��]_��E6W	4�	�Y�_1��ºC+��]�PƬ�s�<�����#�Z��-e���Y�4���V'���q��l�1���3�0��xqu/��rʯ���q��j΋^�C�y�
G���X���YS�$p[��;�Eo����J��R�}�/S�ן�g`��f�o̸C&�����$'CZ ������!x�A	���v9y�?�f^��&�A{��t���_���!�	�r��}|�e��C�sG)�H�+u�Ą�	�?�wpM&O����4�����j���1�<YRUO|-[��t��?[z��Z2�譢s&��S�\S9Ș������8��o��̔���ӅS*�m�Љ����Q��ɁT�W�8+����,�3Ր�|��Ɇ���l��AK�#{j-P��4 �$@���6�%��!"O"��U�gE����`A%�)���w��b�I��s�]�sM)���U�G\�~2�>#<f�vB��tW/�{H2u%}O���<��w����
s�	��O�C}� ��b���Ƒ��~=��$1�xz k�<]xd�q3�i��Pz=������WP�-�jf�(N�����tKw�K���vqzD��5W܈�@OD�.�C�Z�S@s%i-��zWն�xI=ݵ?x�}mS�l�ܜ*׾��8�J��y���aCN�*�ߤ8�XM
4i����.g�ܬ�B��4�������j�t^$�d�RR�R��R�F�N,H���8����@=Hs���A����&&a>F-Jx_���df��FK��a^ː�*���T�.r�d~���uG��L�g�&
���m������Nz���ޘB\q�*ACr����t���M#GG.	|�f����Щ���רr@�{�����rYT�K�O��}K.���j&��(N�w�����H�������Λ�v�M�?H}�%��7�,IK4p��R^��NE���1�x��IB'��C6��R)J޾ډDڄ�k(�F��[�j��TS�v<��mr#��5�	"�h�����|Ƨ�^d)��_hp�M��.аտu"}���:�}$ ��0���E��N�o�$l.g��L����{h��h�=�����Oa_�G����׿ ^���K�&�h���^Z�����X����w�"6�7���!�S��o�������gh��	�Z?�}�����?�?%V>m?=�)?��)C꧰/�����s���G��VN�U���;}���TA1��:}��� b�U�`��_�T z�?���MI$wT}eZkarG��NI�	lJ"���[�!�/�('����e�V)����\�.��x@��g��oݙ�>��A�/M#�����˓/���h����R.���+�{�M��o��ރ�h�ۍ�2^���U���y+�5D�=��F4���G��Ut,���G,� -�;����%�)N�/���}V;J|�(1�"�5�ĸW�`\i�����2��ݷ�����Z~�z��i� ���P_������:�vz�慬�S�>O�M-����k�S�Rs$%��f���#�1�|�pL>��pē4�
 § |d,��F��˄�z���$�m�D�m6�v
�/�s�:\���돸��i򹙮�](����,���k��ڤ��9������ ���S�#6�K��d�6;�����Ѧvh��6���m@�+z'B»>�]�k������u�;A(����.U�ll�a�ujо�v^iA����H���uxf�|�J(�.����`Y�~T�?eu~#�G�/�>������5��x�?v���&�{~�[�#P&]#�mڑ��l�v_�`{�z���\L��y|[�v��j��8�<r7�����|�|�+�cc��5z�i�+Bh33���iw���>T#O$^���f���)��=kϽ�lՎ���u=����Bo���1�I��TW�m:k	�	�vo��*D9� ܳ�i��AٖPy���RK�(4iA�������o�K^��\�ʗ"R.��U}��
Qd�}/#_��')x��>�)�#�p�r���1e����r�=H�jY�2^�0�Q,Xk;�}�4�F����;��������RV���G�����p'r��b��x��ce��:î�(���,��M�Ѧ�G���mBs�&���6P�p�E6�K3��E���õۆ]5g���f�31Xd��fq��s�3KW�o>�M���K��K�g�r�V���J6�4^e�~W0B�D�P�@8ũPZ�@0�	���|�W4\���Qt�ʀ�����:ʡ�m�fl���P��7�v�z��|�$�,��7���B5�6��?�<]��|r)��䥲��p�H�{aIt�n����t�&vKG_��4���w��y����驩v� ��oj�밝����o��̭�꾝u�H|�|zL_��KN*��,X�}+#M�CT��,�g�b�2�`���N�^�z�9x��w��N8$�'�O�c���5����S�-_<�,��#����P�#�=_G��eF��K��|&(��`u#����!�f�Os�&/e�K���,�ï����!� �n�+ S�����M��F�m�}d�h��� ]��cƹ.�9͙�l�:��i�^�3)�L�����.�������!:'��ʎ�S���pH�s^d��G�7���T����^��G����O���_��x5�ɘ�͞2��m��H3����o�#�S�K�̆N]:ڥ�5�e�����2��?���|�-^eB}�lH�+�?�!��p.��KI�w*qK�oD��ߙ�)���'�Y~o��.���F�����rixv]%��G�N�Y��]O��c��$-���-����E��a�)��)���W�O��W+���8�� 5�aV9�J�r�z�o�3��J��B��g��Ϲ�ծ��ˑK���i�p}��@ݙ����(��/�$ê<��˞�����+�8�����͂��D�X��n�)����>�_��x�&��L�t�"���Ua�^`�B޹{?���nG��#��K v^%�'Xܸ������x%|0�Ϣ�O��`	5&�����=i��p�������'.�	5 ��tH�,�[�I\ت��jfoMu-D˝(���k�n���	�/Sv��������"zB��?���lC*O�\'�f7iP���"�A�r�v�	�� `��rp��6�N�A�a�E[x��Q+�S'&Û�����;�=�tn@��f��E��3��Jo�Y�@�M�Eg�!g����m�`���+(Y����!S�E��}�E�|���E�V���*=Q�6���7����+�}��D�o����i�� ���hw���+��LL�Hx�
*��-en�?�/,u�lx����s��j���.�f��șۄ���$�n�K�"����/����z�g�?�@�w��'�*|<�:�V{��1���:�d�N�P����M�p�%i}ŕ�%8�\��}�a�+���y�j<K�v�\q+�>�ػ��3P�"M�:��<U����#K����<;̡T`�:i���0����ů1������W���F�^�/������u*smq���*�4����勤݉|P������"?zb��uT���+N�Ҁ�n���=U ����*<����ݏ[r�HQ����h=�^w����n���G�q#/_��ޏ�w�0h����ͫ=���4���5m�!�-rH'*c�aQ� &�p:>>I\�w���rd[��|�����5�X��1Ȱg���+������\ҹ$�
�G�����ء����T�g#;	^Qq+(���%C���y�fdU[%��2�C��{��3\O�- ?���jZM�e��
RQ!�pa|�D.o"�)i[fXP��L��+z����G��6��:� _��T����O[��:���o#Wbq��7/I7ѡ@'� ފ�b����OѤ���F���?q��Mt~��A{�6�J���b��"q������!��Az�x�?#��^��SЩ�(?!z8VA��G į�<
�n���i�������!�IWA�Cn�HxDG��~�j~!�������@��Z�ku���~� DC�R�@\ �R��+�C���' �/�J��k!rҕ��=�jOj��jp���8��qFK�FK�VC�O�묖ޯ�{NK��<��wAk�E��KZ���?ڰ�|�J����v�N�B=K�1��tO��i,m���ci��t-���L-���aZ�i�Y+? �/5㐍���^�.�,m�~yZ8���C7e��T�m�����ⷮ��B�B4E`?���k�~�V���C��	,���z�EZ\����5I+g�?E��Akw��>����Z�ޤՋ�ǫB�\����.�x�2_�5��>�[��[�?q�7+IO��n]νJ�|$�:J��u�ۭ�u�2n�g41��oŹJԗ�~��G�aF��Y,��x"�c
���G�h����hY<���w������1��|$(�<�V�У�
�SJ�T>�{��V45ms?Y�H� �4U �w�){
9���vAI��1�ە�����赊:�]u�C� ����,i�_]�G�V��n�qM��@��m둢��k-P��D�MO��DT'����4�dx~X���B�����`)�&�%�����<���a���w褩+F�R������!��t]�yprk�'U`�P �\�"��h�l;H~�������+x��_p�ҏT$�B}�oR��#�#Q>��xI��o�i�'0���l����iN����^�Sڹ�!`D�"j��3��:d�|��$|_O;�����A5붨�!$�k²��C�XZ"*]�>/��B�%W��Wc�Zȁ�5���$�s"��Q��A�n������~C�K����t#b���_L��As�����*�
y�o9A��m�(�/�-j?{Li���N�������}E���(&��t'U�ƈj�YT��e�!�.V�fһ�T�!��@X�z(G���GX�¨�yg�T�����x���)���ݛ����{C���/�*�uP����2)�������e�JY�_Asm}m����ߞ%8�eL���� :P�H�6���ͷ��ƞ@M���"��/�k̏�7���ԏ���M�|�UԮ�I��EN�.|�"V�
&�{7��:��������)��S��;o¯k�ޜ���q'��A�<��4���[�+j���� ŗI�#T��X�%`i�v�}A,�!�X���W��B�궄'��k�B����F�e��qq�'Q��Jo�W�1<��C�_��Y��r��~��<����`�6�x����>=��dԡ������b�;6Y�WHH����or��`R������V\\̷���e�!���,��.�� ��?�U�+��p���ƉUF�JZ�7��N���҉�7���X�y~C
���e��L��C�5w��9Sݝ�5���!���ʻ�1�����4����K�+�q�t��F��xr+vi��M��Ս��f��kQ �:�#X�.����������Ը��*���$}i:����9�[t����O?�(�j����b�(�0ȸ�'���+�J��ܧO5J? �'?H�w���������v����L�I0�rǳ-���x8/1r�lA?���Ag=-��hU>((�drG��~�Bdj�uD��o���R�y Ў���?@D�dt���P��;�@�p*��� ��iW���:��-8ǋ�>�'{��ڻ-E��?ƅ��	�3��l�C�%�����u�;�1^���T����N�Tp�2ѻ�Dg���?��x�89���=G�߼�>�}�Z���!�0�0�<����i_�Y�z1�+�5�+8l�Dls����Tq� �x��U�<X? �<"q����QS��|9����Y�yQ屣�ۯ���n���FL�h׳�k:���ZS�:�l<	�=ݒ���W��u������߉ҍ3c8�ID%��v}������c�T�C?2���N�R����Kci�t��=�����c�2�/��$ �=Q�^��p��}��$5輭�>����m>ǿ�J���z>O��W�m��:��[?��wGsCj����Pa�?(t���9/~�ֆ���H���s�~�V�}9xC7܍��͑H�͠�Y�Wk�����������<�����̄I�	�5�DP�6#P�d�$gd����*m4B�-�.���d4����Zk۷��m�~V��+72�d�/@��p��R�%�_k�3����}����̹��{��^�T{������܅�W����m�!���=��^�_�����j�5~�}��F�y�q��{f^-�7l�/�v�N��:� �{�6�e�A��o�4�*s��-��DW;LJ�t�?H�g1>%o<�`�#��H���n��~k����C���9�`W!�k6��|#a�m��I�ߔL܍����d�
�ί�ݘ(oL��y�:�:����@�����_Ҟk�6�R��n�hq�#������Q4����ψ�{����PNIO4��Cf#�70v%a�i���L�,.>�AmؐO�и�GvK���\E�>���Ɨ����*�
��:����"6^�.`��V������ʈ�U���+**6��:w���F����D�$����N�����+�[<��˕���[Z*�%���U�xn�Z=�U��s��2Hz|_g��r�>����������~��wys�q�f��zE�T����`����A������*$�kVU|��ɬ��UZ��/p;��Л��\ZH?E�����Cu8�_`i�Fm�rŭ����r�U*�q	uÒq���Q@JR��&����˖�[;��7]�bB�Ze����e�%/��`���Ñ���,j��u�!l��oG{�|DG��%�����ui�j��%���h_��SU���G�:R�����y�Bf�0ŠD�����ͻ��|o�Iq���u�Ov��$���$_ o�Q|/n�l�������^:�;��S�T�������J{�þiI�����-���C�t��3�6��&�� �L�5�C��x�3�"�~���(%o�#3|����G}���_��+^]��,BS{��[�^��rE���6�i�%�z\�ӎ ���N�;�y��e�����[6d�1��<������#_�b�5�0���7�{K�(Ѕ��&�f%J���"��@����p��s�W�Z�M�cx��<~؆SF�9 ]�#e��gFk�!Y�q/�[��Q�~�����?�ګ~�rꀜ������&�D��f�_�L|�r�U%X��8�TĪ���?F�I��b�����YR��}�l�����Ã��yiY�"��Nmx�f�!W�;�O�§�ź��Y)����:]�ښ�[�ch2wL�0C;&`�Ǖ��ľ���f["������[�ڌ.�<q��M��5qK<�C䡼�%��dm��L >A~f�
������f�mW#�Մ�/�o+}�����I��g�Е�~���4y�i�>ëg��Kx@mD�n�A[��D�uV�b�-p��\�v���b�[���e�F�	K^���C���J��`Pp�G����g����|��1�q���	j�P���B�އ��:�+�nk����w>�f:A`!��
A�E������G;�T]o��T�b�<9(���=eo@a�W��75�v��a�:��^���
L��%�7Uqv�S���A�k���M� ->�v�_�P4��쉛�ܔ0�ُ�;h�W]�W�*E6,�W6���fA�n �r:�[w���Ը��u49P���p�����4Q�����~������"�R�GL�Q���b\4�x�E�Ŷ�j�����tH������Q�>��}���\
Ky�a��ђgS�<�A_�;�s3����(b9��-�.��
&N�8�A3ܡ<Yc>_���B��>�Y��3)/:�*4�\�F��Ip&��6g2z��8����"���y�:�-`���V��4"7��R����"�/��0�\z/�/M�a�`Њ�4}�Ґ�o�4��D�~3�!���G���!_�MH�F�S��{]|;<�[f�
�TT,��#e,��w{�q�d�{����,7����N�l�0`=#�}`�Ʃ���@�O{Y���v�'�D��F��1X��b#��=R�×?a}|I����F�O�E�o���ف3Z\�4`o�oX̻=>��A|/�dw��.��!�6(;O�������]7��p��_ ��~�e��x07��q`<̺Y܌ 𡸹�����d��R����/"_Mȓf�O��+����R㔺��+�@]��D���6&�B�N���ډ��}���av��7�Q����2��阙Ĺ���'ƪQip�X���Ep}:�?|#t�J�o�~�nݬV+�=h�������'+�ߴ4T�W˯Z�]#�h%�YBΓ�^J�?�N��y_B����x�v�ܣ�AK0����G�&�+�V�/셉��Џ!�2�K�
�ź�җ���AV��J��}��-y�9..W2�KN"�Q}�'6V�0��I��2s�w��W,�uy%���W�����e.*T2�챚����/��awm��2e�������(].72�?���W 7�5��r�0��ir��I�B�K8��� ���n#|��1ɦL������t!K��kh����@"�)���!�����x<����Uk>�YG�|���m�eh���
~ʆ}�ݨ8�'�
�Z���qJ�͋�9|����6��|��퓋�t[��J�9l���<�r#��n��^�uڸU-S��p�qZ�W���PBY������5�+y�t$.���p<�VW+��"0��[>�N���.�>_�V)��0��O��D'c<�.A��F-&)*ϥh�޴[��gCv'c�'�h�O�>�z���K��#xշ�z��U9/~G�aXf��!���ގe�SJ8��jQ �w ��h���V�`�_���.��\�ޮ���7���*���%?}4�"FAA��a�t���q���E�s,��x�d��Ir��h W�6c�K����������/9��K<ΡM�1�Jq�4��Ə�2v��d��T
�S�г#���<i��'}�^E_K�G�sԚ���@~սvyu yUc//�!���]�.f���͇&I!#s��H��P��:X됆�#�k�qm?�xn.we��G��U�W,�c�"��XO)�����l}*	?��u��u���͚�:�g�.n�N�ڬ���>i�q�� &'�G��}��~tY���N(�9,#'��d�D���4C�i�t�!���U�δo���A��N<V�[��r����$�Z��k��U��A�A6�E{[*����bzl���G%V�գ�jA�2í�9$����:�ޖ1l��ב���Q\.x�L��,�>�w���M��8%�kO�(�<<��Db��[rX���N���i�ԽO�+,��&Ӈx�'n���֝��gD���}���W_n��
{�Ǻw������� �î�0t��
��۱��y�ǻ�ӱǳ��2��3����U�)R��DH��1���i�+yC� �t_�����B����i��Q���[U����͠ʵ�'�M^)�L�W䦳���]р�>_�ZsuC`�oդF���\��L�������b���۲��'R�*�#hǢ}*Ȑ�2EW`[��)w�e��;$�vV)xs���Ϗy�����;}�%��vFP�Iq)\���o 7؃�����2α0�F9���@/#��~S���Pb7���T�%y�٥��W�~�ݒS?��O(�%�z!��0�^����z}�g|l�Z8�s�zY��K�- `��E`r���{�[�Y���j��p�U=>`�J�Jv�~H�X�6`��@/9W�+����ٿ��$��IC�7���]�}&�|d��U�p��<�N�f�eޒc��v�HWH컖��	1�p��"�S�4���SH����Җ�W�����g;)]q��É_í����J����%e���3�=m=�U��J2�V��S�H	���B�CU�������?�x��IŌ���]�b��S����2�8[����o,q�
�4�y#*rAr��y�����������"zU!�C��bbB���[J	I�VJ�YZ�����J�p�\(&��-5q J�k9�]\�a錯o��|R��y�����uO��l%�/�^%4�)Z��'�|h���� 7w�2��?#��Oy�]�1c�C�Q��lW8�r��@��3��[�b.�[�O��%d`��� X��լSZ�9�>�.��?��0��;eg���} Aԉ(��K�*F����.�o���ao.p��Qw����qU[������������������t����8��n)y7�S��ex5�ua�'��ݤh[�z]Rd����հ�\^1~�@��F�UϚ�w΅�b���Y7#�*��s�$��>X����ŗM��|�ɍ�~�������=؉j������T������A��6fi���O@�k�45V���ݩ���Gl� �e���'�Q3�u��g$fo��������>�RO���O��c��?F#�GS�3(�u3��&��Il�2N�bE�`�0R��.
8p��8��R��`�_������:?]S�x>z����O�M%��u2�+��L7J�&�N|R��Hw�/?��C��/��:����	#��3c��
k^-�.9/�C¯ihw�e���m��u'/�+�/w[�,��k����z-Щ�ڕ��)j�t��a6��ڕF�X,�^��Е��~������G5w8���ϵ;�&��D�|��R+�8Ww�z(p���ӿ��l�[?�����#������F��4���fcV�[п�Kp���T�0�(�/�&<��u�4�7^A�%;)���j����U�9�j�?�%�S�S��cu��^�m��|8�Ҟ��/h�p�E�Em3�e��K��DD�O�ks)ޯ~�C��2���&Y�6;��Y��w7��Bc���`Ef�>X�J9����HN��Ϫ���a����69Ð�NϦ�����l�Bv�I\9rT
��<%=��\�d@�<B�,���B���{�-'�[m��_E��Ѽ�1,��+�vt�{�Ⱥ�/��R�gUG�'_�H��W�6	�'}�jG�A��7��ԋ��Y�R��[*���XV`rd�J�0�'7���JH�S�e��� 6bd�u�t��ȸ�%�
a�펯X,6l5��`P�`ŔU�'��Ӳ�!	]G��qd��%{0�a���Ò�{�]~ǣ�\w���}��h��7�d�{oK���g�X��G�*���rI�I�}�-���N�wn��e)�RI���6��$^�O�c~B�2~����&t6C6�I%��7w��s�x���ud��icSd�u���NI��'�����3�N8MLʕD_��'���|6ܤ����x���v�JK��m�`�Mg�3��Հ�+lJI�����'N���{��=���������NV��j���XLZ��`mmm�!�u�%���0�hҳ:���ǹ�톜�C��܅i�TZdl�zi���_2���*/�=r?�0>�vF�Nk��(ܾ�|w�D�l)�G�]��x8\
�=�X�b\*}�0�)�;�R-
��ǚ�G�Т�ȵ�n!��"4SJ�9q�?�+��]Ė�6^οh/�d���<�E/ྲྀp2�XP��?��k{0�3�rx,���l��$H�C���^�s��.U&��/���J��~>߶���}wM�@슨�^�⯦�5�݊����6'j=	��b��S)\H?�"�	B1[/d}�?Bu_ض�2q���-�,${�8��Sb:/zJ,f�ێ��w��������f�.��3�v����O����5���T�iD��q2�^�E��g/��3�VC��鉶N�ic�;^4{�_���
�u�f7�l�n�K~:�b��8"�Ew�;�*�Y��N�߄?l�P�=?=ɯ7���2�P�IUߜ�����dj,�bk1@j��U����x�<q+��P�}k.�ZPpc����h��VH�g�[V
��dEwh-w�����KQX��?�5Ut����.�����|\���Ek�3�nN�a�ՓYw�(.��1�����P�j9xg�l O�ĝ����Υ�	�B�ْ EtfH��%�S]�;]��EE07$	=2��ΒBCV��	�푅~�(e�H�}�mV{ӟ�O2�?	�_��W��B��x�r~J�J� ƿ����\�+�Pମ0���������R�0�:!1sG	i:�����)�ٜ?17�{97'¸�<z5L�+ĭ��	~Qa {RDY�O�m�X;4��]}�jGM��%�('Vv��՛��F�kC�$�C	@`�h�B�j*V���*N胦�� u�q�[벸:�nR��~�DG�o���L��tx���<'���}�(	���o[+@j|$6'�R���ጹ݅���z���-�7޿�лF�Zk��e ���A8r]J�U�\l�xK���V���M.(g�V5��mE��.�s��Z�~S�cyY�4쪴�}����� 0�	Ej���k�'{��;�ш�h�N�8l�(:E�QX�^�Ta��F���*5�ݔ�*��f<��3v����<�sV��'!U�_��'BG�ʄ�����Xp���z<�3� rS���$jC���:��0�<�
}!��v[3`��\��6f)�%4j������e�Kvc��C�OǸ�\H"��c�w��Q>���"!�F�"T�<�����L�̋��d��{�@x�l���m�Β��l{O�M�!|�t�i:�AV������$���Ƿ���%
���5d|3��(��_^�Ns�4P�Q�-/N�t}����6[�Tsx_`m���k`�-"@+�����}�
��.5�$��!���9����4?V���s�vh���J�)�,[�2a�u�j���]I��l��c�K
g�P�����J}f��QlE�@�>��[���j�������o��l�U`��V
�tm,��r�Z%�@B�"7F�A���3�V���U�Qb��xٯ��xn��^*>٥�ގf��a�����X�uP`����pU1�u���2��ѢX�-�ͤ���K��v2`���0��k��@��H>z\���?MEz/�A���7��Y��m�ܐ��-��"�&�M�x���rp�hm4�;�b���БI�����5�:j�aJ���\�.����:�Wi�߸�FK<���x/�{�wߐ/�b��X�i�F�*}$��p�	6�Z�j�����t�
���H���(�����^<~d�qŃ��{��>5�玻��:'���82�p���ٕ�l�}Z�oĮNE�u�Bp��ޮf�V��Ν��$��������.���i��/�z�tV(���,R�]����_Kĥ�N�xS0�����o��+���΢��mI��n������$�L�=��j�Q�q�=v���=H���������֖*��r��^�o��G����>��9^�~wQ>�]�o-���wY���w`�ya��^룍��6٫�ô�%��x��=r��ＱC�^m�QH� ��8����)Cu�^Y(1(WB�M��"^�>FUnn,���EX@we�Y���0ׇs�֦{MRX��a����^]EL��⪛�&s�Hj��GMȮ_�5#[}��f�V_��a}e.<A	�@	�w�㯦�3�jO�i8<�ٔ�J>�U�+�D���^����`&����~��F��-���e6+������&�)m2e��(C[USB8��S\O��)!n<��@1�����_�в[!i�+�>$�߽fT�8�~���s�wl�vD�&�	�V���Ng4�O�a�y�i���m)�)��Q-|�m��١��Q���N|��������]knl�P@�F
ȔE؃�3޸]���̈+���2�ko�dm�k��p5��Ǳ����$��B���?��q��ϑ���n�:���~��`NvqJ�g%����n�W�l<��� }���(41�����y�K4���?�������	����L�ԥ��)s��[�.2α����w`M���د�7���d�&�B��vU.$�0S�܄W��E=p�O?�m?�	�0�c�/��2[)Y�9�N�3X��UQ^%�o�B��
�U,���+����ʟ�&E��n[:�~��ݛx=�vW¥f��(��)@~*�X����b=�d�BnW;d�M�W�=���m��3^���nBC�V����j�n���VA��1��b4u��O6b-�VJl�ܘ�ߴ���\m~\�� %��ʕ�)�mix�6oJ����E4� |1؊��D+�F��� �_�-��ǅ[�����i��!�}�Ē�`�����sc������蔢���S�J����p�w!��Zl{�!$�8B��p[r%Œ>H��}��q���9Z�^���NǡX�
xX2J��o<D��_=D�W�O�=P������)��D{9/{'�)|����c�3���y5��hn4�%j+������>H�ϸ�����%����J��M��1^��l{6���[<���dn�W�mg�~��U�F�����L���0E��W�(��"�M�uLl�K)�e�`���N�>��0��1t.����&�i:G�,�ߴ�1���@w�K@�f�f��{7�ꃊ�Bi��Tt����b��5+�H����f�,�2W^`�#�|4�=_�sS��d��~�kh#Y��y�R��:�F8�O�Վ�a�Sg�����T�UD����=Oa��:\*S�a��p�Ւ,����5�k�dG���y�w��	�̖��()�y����qs��I��a$�%�*��{=�3����؈�
��M�7oD"�f��T��K�7�,`X�E덥XL�M���u^��S�E�=��^[�t��,�����T ܏*��ڨ�x	9�U�jȎ���f���-)���G9��D�cI��D�����q�:�xz���a��<d{|75]��M��v,>�܈�;�W`����.P���1m�%�&��1>	L�i�{�Fk�<<��tb�A|��O�a,�����N���ߟ�I���K�o2�_���ǭ
�ob�uq��L�����+�a:򢺫 VS�`i�Ev�z��$���A1�hn�H��?��V��+4��S�8`_�=�\4�&U<(%�.�c5�h��E�r�c�~�`��{�ˬ�����sc�h��x��/޲�T,�"����H���r��
t&U/HYߋ��H�o�S ��6\l��`���L���K��1���Xb|����}���r��Kˈ HJNb�Z�dO��Y+-3�^�ϢR����e#|
����ץ/��	�r���ͳg�za�+�2��j5��6F�G����%X���O���n�2"ēG"�)��T�h��=üN��)S�\�����������v��N��%V��d!4�>����h�P6�Ń���͋�B����ĝ�9cI����{yV=J}�q,)R^�Y�p��r���L٨.,�R�e����\��Ma~b��MT�,��?���*�	�Ƃd�/+���y��7�W�4�>�ꗕ��D��[R��Q�Ձ�_w��Ƣc����uv�1ڕ�oA;R����kж�x�L�
����5��������/��S����.|��$W܄x�Y�&�}�=�Q�2���.%�w�y�������eV�X���)��#듨�	c�1�s~e�?���b�,���ϧ�R\]��S���`^�/sI�W��~t�Dԗ�#w'���7�c7�;Llm���B�a�����۱ѕ�����Ys#o�L��h���huq�D�e������O����ȶ�I{���6���Z;�<0֒9����<]�&ni�@�� ����R�6�?c-����@% �ao���"���0��y7�0ڝ���<6e�5������YOW]R,����a>���.I��,��-b�#�X[��d���T[շ������^џj�d�=N���|���+�O#7��8ػYZ�;%q� ��������g�"V��d���-wЙ<���gw��/��~0��1�1fCH�� nF��}�O,���&6/c�=�r��Fֿ}��6��Y*������2�;E��A��J}�x���>�<�#g�_TćbA�R�
���%�Q���P��M�uRs�%�'�SܢaUC�m��{�}�v&���4Mi��	i�_�@���ېV�ϣ�[�� ���%��35vKE0�3Z_l������64�$�b|¨��H�#Y����Ù�^����A�[�6w_���%�7(Ul�u+��o�1�`�V"����u�E�}�x��|���+����ʽ��,z��	��=�	t@Q���h���.�O`�Afk�7�J��-��R#�����%�h/��3�$J�(��Z�s�G��X�k�F�Q����������Ԏ�wu��H\��� f�S2E_��0�i�-��x�I/T�5=��1�݇F��ƹ�vj�w���C�͛7�����X3Tg5�I���B�a���N9��i� Qk5�Q��g>a�=��ܛ���p�6�E����Xv_X���z�K>g`�-O�go���Z%��F3��x�PO�;j|�>n�<�������(�Iխ�|��%�,��{�B��|U��zY�����:Er���Fq��~����gL��b��15}�	�xs���h������
�>���#2���`��+t����SX��yR�I��R���i��8Ï�{1e��B��L�=Bo�6�{Y8m�r���GrϤ�OI�O�W��XO��Y��������Ō���y�sV�z�7����?�;����A�����,��מ8�D�>|P@Ѕ�}���џ���݃�ڑFy�����.�z�V�%eÈ'F����J��a<_:�7}H�����+��&��<:�*/�����! �'pv}OYod�h���?}&tO'���A��p�Nb���β��Qtև�n��5�Y�7�r<}s�#ش]��8b�|C���P(>Z��?�p��z^�����w���1u���;�AK�Y�e��+���'�3?���ځl/ܤ[)pqF�/\Y�G�0@nQ��v��kS�@��A��얊Η���',�|[�h6�� �T��(��?������kk�۽�rN�&,f��B�	�?lN�ƕ��e�`��_�}���T��a=��@��;`j�v�w�j���	�y�^���>�Oᱨu{�`�p`�)+z�W�@���͜�X('H��r�q��ؿ��p�G%��{������M������	���+�+�,~|S��;M��o��͈�	�L�sC#�����{c�W���`�|�l`�3֍.y�L6���`���)YO�w�D�8n_�؄�2;D\I�h�vhR��!�|�#-a��!#c:6nG'��vH�^�}�����X�.�h�@|f���!��2.�%�K��q�~�~���UdJP�p��)L����f�ۄ��`y���?� ��<)���F�*QQ(����D.s�,&x��CP-J���A�C���ʎ�KZ��V��~C9���ZY�aD;�*,.�ڽ��Vo�X�zg���r4���6�dwG�� H�����S�>������k��h��:��a�ݭ;�ۚ6eÄ7;rY�����iz�F>�;�{"7�:3�]R���[�S۬bd/V�Z��d�q6��	�Rf
	H����i��TQ&R�w��K��G>��3J�2"׎S�^�|XP�k��yLUq�tw:���k�X����%J/�,��.�i;�rSpn��=l�ٝ�5�*�{1t�"�Z̰5y`�J@�= �K��=@�p�,ԗ�K:���cMϗ��}C吭l 2n�f��[��3؝��u���U����x�� ~�)z�\��Kx�T�����/ѩr�_B�2�e)\�K0�� �#�x�|�K�;S�tLӉ�U�cnԘH�xa�Ĭ�`�]��v�(NPę�/@w?�^��d5�Ob;n.�F�_��JY��It�C��0�!"g`��vB������q��V��Qܸ���u7�P4N!�NT�7� &+����J���h>����3��y~p]��<�����J��X���ƋCV���_.��9����=�)T�P��ȫ�^f��!�_K�LC�r-��
���Rܠ�̓�*�$���|{� ����qWC�3.<���9����U�&?�/�Қ�@ӌ����v�d��4�����s�ǆ�aE������uW$;�ފ���ڸ��dD_?��G>d��[���!��yUL�7-c9��!#�,]R.���9���z��D��+ v�a���2�#J?O�mo<�<��x����4{�٤��mMpn����Q�4���+�=E��L�ߑM���ޢ�|(��趉��k���|��W�0i[����A,>�����1��4~�: +�aO���/<h���)ʝ��P��nC^q�����������7�m�j)��d�mf��J�]Dæ���]���ّ�)�F�j��v��/�uً���<�1��qn2M+��n<�M�����?[�k1�bn�<1Q������a��$+����vK��q����e�`�Uا�̇�0|�d�Y��0��wN#��JM��D��4�$�P�d%G��+�NU������XL�Yv5=E�_�"s6�'"����3ѝ�q�T6�aK�K�v�ݹ�����%;�8�>����^>��"�p^���.@9[��{�\д?���Ӱ�ˑV�"z�=�,��k�v>ؕ�d*�*V[�:�kֵ��\�d��y�u�wd��V�4kP�,:]I���+���K��],��!�]����+��nW��@o��U����0��XW��xӻÏ!_A͕�_[Iy6蟙���?L����I������dҟ��rb�-��h�u�L}���lМ�`�E(�*zU)���(��	��yWqӑ�3�}�=�^pcQծu�ic筝w�Bz��9��"y�}������H�������F��"�R�g�0Z$Ö�Y1������@Sz�{<_��?��p�4��'�5��oI}o{�|�E�7�&x=\��[1G�N�^Nv�����l�7>�=�h��$�n;s�؂Ρ������կ�:�}��[�^�ɦ�I�(�WF�JI;}Rlũ[4�+�Gc���/ܷ�{˦;��qq��K���蓫�C����>t~@䴪��'����꧄&��|)H�?��-Ў
��	���!�-�/����?&�3���@������D?��*�M�����)��Sq���Ba�R�+�A����Ժ
�M8㝟?S�h��oF�����?^��B����^�O͒��?�<�=���^]r���Ȱ�ҡ�k>��t�����E�)��'}�JG�~�ū�H��E�+���nԽ� �_r������$��'�W�q�Y�Ɛ�,%��?֋=ir|GQup�X�½���Z_\j|�އ��k\�z�xPl���0��7q�p�����4���67��i�K��7��.�m����܅�k�/Л�%����p��r{s��4h�2���s�s�R &����	�ָ��TZt�H���W$��`5n5WN�w�ўx�����_K��ȫ�E���K���P|m�`4ٰk�k��1�߼Bt9m��{������] "�L��B;<�V7Sܲl�v8#���=S�������w�Pr�-jzʗ*Ӛ��.��Nk�����a��&��McXM��[����x�}b}����g� �<l2N��F�@kH~<�pO�ئ�b~�`�SVLPW�d�A��<���X�?u%��7�tJ��@���#;���j��&�g,abV�Z}l�rx���<�&�M>�I9�Ĕ�{�Ln;���~�j)/�<<9���І>�k@+����S�F����x���@�����S�X�����}�c�ʎ�d�A�(�0�#�.�e��1��b�I����e�84�ײi{5S�V�r肉�A
�fsѿ�������bk(����և3pߚI�8͘r2 G�M��);&�6C����ˬ����V��R���4<=3~�S�,���܊Q��>�vI/"�|�A��B2�7A+�����}D��!@�Pـq��v�~���������������<�av��V��ʎfw6��_1�2��B�\�t�f�u>�2��S!��ݖ@W�O���F����i=�
/�|h)���b�"�b����ĭ�7�+m.�G4`f�0�ƃ�h��<�14n#��� �Ώ4:,�K�Bi�\1�i���c��Բ̧1I;򁤅�F�����0��Ƅ�xGސ�f!('D��=��Wׇ�>s��y.e?�ֿλ��[a�����k��#��t�/�&t�ؚ�͋f���V�nSν��8�d����|�Ԝ�T?s,pr�ߙ��ϸ�D)�C��x`"w�I�G�FV��G��FFSΏ��]��Ў(��,�i��ض�:�:��~ ����䶱X����*����E0��*k�%�`#(����&)%}�`^�OR���t��N>��כ���h�#���f�ѽø�����Y�{쟰m®�Z��y�=��B�=jCg�ļ�\;lM����
Xad�W$����JT%����t��5h.ء�e�|�3�Fh�����]l4y_VCN���#TD�~���n=����f��$Iӯ�5��m�o�X֕���nB<�ZA�in(<w�|�mǕ��G.\���y��_�^y��Ř�,��^��Q*n�dF��l��҆�``��X&���b������4�/��^��1�:��gNLO�Fւ!a��fW=�6�9C���΋�*Ϫ��78�6�w�����T&;;�n���p�x��]���Cܵ��y�
��m�P
��v�7�KBJ0��lX\��5�}��J� 'YOψ�Ĩ���7��ٍ+�]��g���� 4*��:Bc%�A도���h���nT0d��k��2/�����M��] �H��Mg�}C]x	O(fUI���8ՅP�/�yd=,�QL{�g�Gf9�7�����`���^�|��1��0��$�i��!����{M� ��SL0?=�(E�� Y��s�{��ѕ�[��n��=W��4o�8�A���ȳy�;��|�k�/��]v��
C��f�*���7�T��Nw���`�I9Xd���Q�6ͻ�!�yXl�Cێ��^�����!tk7���Z D��K��cib�)bf�8�^�uy��W,�CV��0'`���`�$�������g��J�F�<�v���uH�i����e[0�9�AX1ó�=���~L���z@n9T6P���p@��!?n�	'4��C|��_�[�G}F� �_�C9ũ�&��11e�l`�kh����r`��u2ZJ�:�%9�'U(�s���	Q��V��<$_�����čqʿT�Ne~�]�F�R@��w�Eġ�sw��[��6�AҊ���{�y��d��mhO���A��]�*{Sl�}�?���A�oHxH_�l����Ȃ��ᰒ{��O���&��SA�zh�	o��y�DN=JPY_�=r��e�]�
�L�N��v-�4��J��& ס�nk1��0:���؊ f��
�F�۱XY,�]�� 4�ڳ��������"�^9�u*��i�;�^+1u�^7˧�2yn`=�E�4~�ș�~���)Lx�t)������EE��~؞s�J��Jh�Fe�4�n?[?>��K����{�L���8ե�܁��#�-�&]�?,!�^��o�Q��]H�s��Z�Рm��w���D��y��-@t�+Գ�B?'ܽ��g�\ܯ��QW�z�9���7��| ���k?5�+b��P�+0�^�g�̱[K�L�s�_L�+؉Յ��/������?���[^�Gy�^6@ޒ�^Bv\��������/оEZ��`݉�:�.r>�e�04H+��%q��8 a̟2Iα<�.��b�jE�b�M�W,h��g?�莸	:�p���r����#n���?@S����F��~7��b6�=ۍ��[�r���S�	�+������\�>��5�l=f_?��\��;�_6�O>~�͇Ḿ��8��v礼�	��Ǖ�����~1���x��]�՟�Nz���'�:�1��!�[�KpX��-r�򠪓=S[�gy���z w�Cf�$]*�%������ե�zM9 �v O�=�B��]Q�.X����+����%�!�<�P�a�N�#����[w�O�(@�y���`�ua�(Фb�5y�������,��(�M���@���	��f��	����ev�\�y>�5�
���=ǃ_E��v�\��I͍y�Z�N{���T��x^";�K�mK==6D�&�����^N�7Wt`U_�+��ʼu��k��" �+!�٨�/P��tk���B4z:�Wͅ�q1��
N�|���I}�,�U<M�����?������ܗ���͂����9��̮u�t��\��a,�磊Q��.����N�9���g]ʃ�e'�	�2�$��s�Y2�N�W��u�����΂�"m{��W^A����LV[y+���ۣA�j������M/"�h$�ƞ�O��;���փ��O�ؚ��0�?�[���Sl�N��MS�:��l0����Y���IYY��mM~�yv�h��rh��►����1,@
��Վ��ؽ�`>l,쟦�:ڃ�~<�T���.M�0׫����a�oD_�����{�͊����z;,S��������;�&���T��w !�,�?���!�w(�A�^����3���-��p����i��SY���1���jjPP*����J��,�fȉtid~����I ����Tf��̅�`��BI�g�5���@_�
�x��Quk�Ƽ��]��;-��Ѷ3�U�:Hl��K�o�%�Uǌ�5�8TP���c8O����E���{�EʣGɄ"��	Ìar�Yl4r1���fx<�:�����S,-*'�Y�~nl�1��ǂ�Ga���÷��ȇ�aA� �FP�s�W�xtq�a:1z�������f@7`�u���V�����	�pBakVl��xg��w5��8׬T������f�������5���b\e�00��~�.��b��?�1i�y�ܔb�M�Db�;ܫ/�Б��=/��#�c)�p�{�4T#�>��
D�[A�;f�y稚�7�Y���� =�����U}jB85�9|��5Te�C�X��A#-6[|���:^��5�Q�7��b@��[b�11�z.,x����\;���j���v�~L&�1k�4�Ci��Deb`���;�V����ۙ�V��e};�f��h��j.<���%�8ق|�"h��K*N�0?;=��d�SD�i{6� WC��.���Rqk݂`��o$�R����{A�����J"rԳ��PF]�n��݉��k@�n� �`&�6�jVG���7��.cq'���n�Y��:�0��>�7)�<�^7f񥊉t��P������	�����k�x�?6`���;��<������g�M���$�P���\�%[�i��:S��#�C�zc�N����H�, �Y�n��Tt�MȷE���'�nD	E-$�<���$KA�E�~�-�6^]6\f� �`J=��p����K�ʏB�n���śS��'�Gxʆ�7 g�W�i0_	���^"9����-���)J���"��n7I{�غ�v�f2�k�V���������=˂.���/���>�b}�K�T��]afl0�H�6��Vy#�.�s��-��{�0<Tkwe���!#46V|$[`�|�w�40h�?@�N	x�S�u�a�$�5��g�x�8�'�eDu����4���8�����?���#�~],��h?���P�sm;d��cqː���G�`&:�Ӵ�mS�a�AE{h�E���sk0m��~��۝mù�]/E��+p�o��%�ҍ���kqW��P��3�+��n��B�$^�Ư#i�����/���NBlZ&��0~�1^�/��_�!�I��u��ҝi�Pq���@X��D���y���,Ȧk
QtpD�6��Z�W��[�tJ\6��1c�sYw�yP�!�3��X�;$V�	�������v�^It	_�ii&�s7o �6G���ӹ?�3UK8�{рD�ƹ䘒�����9����P�h�s(Ř2��)�ϛ�%y�����E�=���Z�������V~��~��|� �N"�_�]ň@Y�����R�R)��ơ�fQ��?��fTIlÒx�7�c�X�-�%��v�x�k�GK{R`ا۪�^zy�=0k��J�0D���-RF�UB�б��j��B~�u�4�uI��n����Np�`o�sI>
��ˈ)n��B�<k`W�/A>��3V���nC7q�̼h?�z��2�V�wC�+���ⳡE���3~�W^���[*/)p��ğt��L��S=k�6
lF�&�RT^�j�e�OV^Zv,z0��ī��2���o�������1�(�; �H������^ހZ�a��Ye��'�H�Z�ӳ���!�r14�I)V[#��q��qK��ʐS�������)� �7/����ILx�X�����c��*��D���e��ԿY�k��1�Y���JW�/a�j��[�H;�����vz�T�b����-�MJ��l\���D�p���.��*�?��SӜ������eF�u�X������|��]��zy5?x�W3p+1$q��d�����sX��z-z�����0�c�]5��KqS-�y��m��f���,��[�#��h��5O�zPbe��^Iw;$Ͱ��F���.n�<��u�:��^]��ϗ�N+^$��%v�Ab��E���W��/��F�֖�q�6�d�<�X�G�2M
�?If�{4���=�l^����9cu�V��G�����n��M|�S���v�ߖvy��$op���7{�uPdh�u�X�F5���(h�7t�^��G�zs0�y5sH�U��v�ٳ�*o�>bM�1�<I�j�®��V�<S���󚂄��V)ק�*�D̏pX�Y�4~9?@5�P��'�������G�>��ފ}�j�.Xs���I�ߕX'��w@�js���ٷ�ZoIj+B�V��V�'[_�_ޔ�3���s��ds�|-bU�dC����C���˦�mn@
)a �n��-`�������4Ll-B���h�T	�ј[��-*�[��J�:l<�	�����c���_�S�4���S(U��䊌�	�c9��R|*93�Y}]�u�"�-h��=��+�Ǳ]2���8�-����>�i��_?):��XH�����t�f&���]�tx���j	�OY�vx�zgL���y��K�J���������Cy&�}吏�Ǚ��p�e'�k<����v�c�G末}���_~�����-j��<)N�)ꃱz88�Ճ^���z�_�|���T��뙆lJG}v+>�<�p��0���.�+QoK�/:=���ѻ��ګ��&���5#�[3��q�ꃽ�M$���H�OB�ϑ����աK��v�E9�K�o�k�0���R:~�78%o��@�e*A�>��1�1l���%�`��uwNWg4�nW32�S�-vV��#����R�6PA���5^[6�Y�sA� vzv`�P�cA��&���'y���o��{�����*�	��>/n��=��1��zG�+��)�=�Bo�Z �`�=�iM� ���E���#}޴Tr��f����t���^D0��qx~.n�T�_��^ᄤ�ڪ`̳�U��`Uņz5�Hn�� �������Um�C|bd�{���#�o.̦��hI�X���w{d��{, z��f�W4O6�������Q�ի:\�%���ķdY�T��S�du
M�e	�Z��u7�y�L�"@͌�'���@�GH�OuX��J�m�Dژ%u[�R�5��U��7��;0<�3\2Tyu6��Ït�K2��`F�fy�[E�I�䘨m����5��N���z��[��q�Ř '�IW�7V���n����k�4VA�fy���I/��O�2�w�`�����{����k�6��:&�	��}/_�,]����1���_'��W��p��LѬ��zh��Csu}���@���*�w_������&Ԃi�Mӱ�F�E�GW�������\�vT9��C}=5ʓ}u.!6w*���g�c��1W �>�2�O�;�T2���	��S�8<!9dq	|���YWʵ��x�Jl�DImT@�z��|怄�M�&5���V������?�ؤ,� �����h�Y\6��֕b#�?��ME���Խ����
�_Vw�d�@w��Hď�Hz`���%;�\��N��B�>�E}-@�E�`�F�;����d���
qۺ����������@%�o���J_���\
�������K�����x����7V�����#pOq7d=#���u<,!s��rbt��%�)c}B�+���sT�
b�V+@��'�ҖS��:�5�U��1���6���M�78,b ��U����{��1�0�W��f:�n�<���QF\���q�m.��ֵ%�x!F�� s�x���BBXu�_�Vs�˹.����猙�k��t�<�~#>��v�����k1�:O7eF	���B�3��	c.���.���הu�-��=�/���O)�)A[�,k[Z$���c2EO5���^��R�=�=�����5g�a�m\�O��[�<��5���?�7!��Nt��xA�2e��T���_.C�h��ƙ�߇���F#:�}��h������~�`��/-*���~mB6a���"Q�T{�����.e҄�^��p�ş-n�9g�ӥ�����i&����E�ef=��zl��`�kn���-�����m��2�n���m�����c��G�;ޖ�Q1��=������XOL�A�(�P(i�bb���_�!%V�5�����;'��Z���gS��W2��I濶�:�y�jCu�x1�ֺ�R�ڸ�Z|<u'��+���U=e�	z�ٹ\�z�J���$W7T���@~A����+�Ò��}�
���R�]�+��>��I�[�ԏ>�z�~��GF����ɿ %f)O	r�\���v�98,Y�D ��&�#��RQ|��b�1�lW<�9����Ο��O�,?s��g��ݲ�v�5�ey����7��`����Q��(�:���Ge��,z���(O�]�1�M�'���g5�֧/���#����?�{�H#Um"{J�6��|؆2� ��^tj�����usX�o��h��>IaU%v�]ꮘj�kU����a�vS�(�:V����z�j�}&N�e���+�;�q$R���f,���>�[��*��� ;��d�b�<_R�j�H����a�߆`�)=/)�v�������#��qI�r�����\�-g�M�D����-�l@`#m�����喢4�٥�ILZj�W��7�,=[j>=i�5J���?�����_��^�{�������-Er�w��.�!u� I�S$g��yp�T:���i)_r0�!���L�e�U���q�BYܚ-��B�>����O�w��S&��m(�lCZ�?ׅ��<>̊�d Bi����C���GE�>��NmL��Ǻ�"D���֑�.�N���-\h�9�6�c
*��Y���a�6��jL��p}�9����547cGo����j�{�P��9���$G�� B%�ia{����&� ����Ztu��Ɏ�4�Fv ��>�ƍq �ڻ͛������!��xyî�U7����}	|���N��l�1A��J�(	�YE͚���.��]�Kn]Mm���r��ٵ��b���ھ���m��-��A@p��,���t�%r�!	���~�g����_?��y�g�������l���@�?U�ǥ���;�L0w9�U>L��P>o�(U���6Z�!�э�\��:qs�M�+m�%��nO4f��u��7Ĕ��.U#�1��iB1Rj��i��K�:r`U��|y��D�.��9i1���z�p�Vo?~"v^Pr���<p����W��uX#T@�+Ue���!羠X�`��d��a��x�	z��6�HaHZ�����Nl�����#�=�=*��z:����+�����;s�l����zZ�aX�N�o#y6e��J��R+��3`���-���e��3�bE�	��"��T��t0�m4�A��<�klr�	;9��/�J����i�=���?������X(�u��rb�:,���of��;��6�=#�����]�N��!�����K�X%(��QI�kO���b�T`��H���A�Z�Pw*��'�����!ȏ ��M�ͩ<�<�oPR�㚆T�t�N�V���۵�`�(��@< ���!���Gʬ��fv���S�-a�JO��p�c (V�̔�ck��[�F�i��n��.ޮ��X�3�F�8�hvȻp?�u�m�"ٸЭ��W��8O;�r9����#��j��)�_8P�I������ݬ��?��=2�V��?�{7��#`���?q+U�.Op��,�l:��,
����t�u�b|A�:�u�
*��X�^�]��#�ͳuW�9�:�r��?��kB3�gQ��؊���_������/����+q����S?&�p5�j%< ��_uN�:�\��@E�-!+�ђ|^��S��;k?��Y���f��ɉ�h��K'+���Y�yϤL �N;�h6m�?��������#NT��9&�K�/irj��#���_��6duU�{���g�8( ��~އsϩG���PE�n�2�y�_��V�ې;�:��S�w�I�'��b%��sά���������)�+7;�]�v�5qbLAYu6�$Z�Y�
�l$	�i�f��r��!S_͕uT��,�n�*����4�)�E�a�������a-h.�Q�r��{[�+��U�d>�2;�n�#��~�Sak0P���_��tD<�B�x��9Jgb�<�g����?ƙ��8%ȫJj� ���b4hc������!NP�x�S��=(������cڌ`���Ϧy�y���f1wٶ#:.���,����?���e��0� �7*�v+�K��s�+���C�30�=گs9
g+X�3��F��k0h|��CjH��WQ��>3�I5"��N~Se^z�n��.��U�TyͫO{�&�W��L�Aw�4�U(�ֆ�ރ�D-�p���HQ���~mV��(�	ÿc��[h���H�Z"K��ww�-�:�[��d�b\�I=�ՙRO��w�||}�����>F��k�U�:A���YW�s*\N��d<\ɨC��a����<p3�m:��7�s��d���z��)Nb����f���hfQ��������[�"�ᤋQq����L�H��sc�.r�o���AHx��Ӳ�%x���FZڼ���Vx��N��sq�ԫ��Pm���d����������><� ���Q"�Q���t�Q��Ǹ�]����7@W�x�7�Z]�%�Tb��%V_��1';����IO+)��a�>�z,�*u�cx5:Q����qi��@�|h_Wp������l��1�N�5�M����к��J�+�����V$Y�ڛ\r��PQ>�xRϵ4[x?E���}8��hF�[��Z{4U?��ha�/�y�����=x�׈]���dq0i�V�Q��4�q�tt�8J�wB�5�An2>�'ް|X}�x2"�]�����}��ڒⓅ2�d��Y%bR��������.�wX�e��|}f����_!0��	�A�
n��܀YƟ��&��䠵'{��n}������>�X�V�S��~
���݉��w�w���u	n+�5��Soޛ��>��\���z`ueQ_���!�&{���W�WC���3�;���ceD�Ԓ&xZ\=�6�/_/��g������H(�O�f#v:D��{<�=-�vb}���W�R`Ȗ�M�~~��#������s~���s��9��{�V�+͸&~_L����$i���^0�Dh''^�,�������#�P�/���8��7v"����XZ6�����.OK94��<��{{�����f�?-\�C�?�&�3i�H��O�����h��[�N�߇�ٍAl�� ~��(^y�N�9yV�_���}����P�2Z���[����q=����\�h�e�t$>���P�O����D/��E����{τ��m��i|=ݚ���a�X���(�L�o>ʘ���iC���${�P����S/�N�?�/J�?���Ãp�l�N�����.[_6��M�v�q���8Um8W�8����+�Aw����yy�j������`���?�V�8���x͞����K㩏A*ۙ���Z�J=���i�3�S/b����T����_u�7c\oa�E��G@�H8#�����l_4����_$�aU��Ʋ��8�0�F޷�ݥ�v{||+��m�z<�s�����0��x�/y�C3�����8~�����U}d����Ѯ5zJ ���=��`�e��,j��v��l�
����<���G_
 /|Fk#��3�(�������N����>x4���^��H��A|����T}�g�=Yv����giD�ś��^<\G{��2�e�)<��\��	��5��-��x���S$� �{�g�50w�
�'p⧰�CޗNE����oz�nn�'�����-P9�6�*͠$����՚������K���N�H��k3i��'p��y��P�2	(��Ԝ,j�׫�W�����i�f�żT�h�� _`���l���I��x�=��Op�C��M@yAA6�9W(�E��t�s���olu�O\�����)2~QJT��7P�4H�>JP��b�z��^�,���\�����p"#y!�m��w��U�_���=�����&`�ޚ��)�tdk�y�M�����=��T����QC ���G�71���$�B}_$]�jxs�<�`W^@�4������ �vE�y�`�~�EIo!-=��qv%GT13hĥ�I}��G�����,�Cn.W�z{�N�6ΎBh�Z@'��AH����\ �������w5������v9;슲����c�M/�ChB�{:�����������8HIc^i�QS�4 o��q�4ƌ��Y��/1{C��g���^=�qB�����e�N�f��Vm����2���w�h��7���~9}Շ����."TWFM5���S��[��x��$�N��%� 0C_M�Ŝ�����$��1ãQӐX�!z����7��^���?����e5�25��f���?vG��I�S[A.��X�FMΉ�Ι<W�.O,ފs����-����3/�ʨ)kb�b�^p�����}'��)<g`��a>\��2����^��Bi����ՇP_/�M��]�0��܁��[>�7�y���S���:��6�ɶN������� �#k��[g���q����u��a-���UQ%�
J6TeШUq*�$S1GA�Bq�v�iaP 5b#WƉk��#�	ɸ��"4�ZX���C\�j�s�at'^]����c�qY��ʞ�aK�!����)3�c��f>TV���֣���_w�#'dH�2Q�"��9%���N^?n��،~��gg��Q��[�������uKp�[K3��.ܳ]�4�����%�j\r3�ި��@9'�Ø�e{�0���~��,��k,v����xߟ�N������O���c�\���s��L��b�w���9�x����;r��;�;�������sg�秒:���ȴ�M���O0�����A�N�G����x�r��]��q�ȗ�b?kh~�pa*fh�AN�P��߉�!qlc�^�[�����*	�<��ͦ��l��"\*(�.⡅�B :ϭ���[~�anGOeU���Kv���'0����.l7\�F����o�f��A��HM`g��J�Vd�
���r�U���g� ���'XfT���`d^��KT'y�T��ZQl�C���mE=��=�kB,�?Ϥh�[+g(U6趘Bfi�WCR��fF��?�y��>|<�=N��?դ��_���'� 9�Yy('�f�zh<�8�/Ӛ�6��V��C���煳(v��Y�غ�|��!���7[W�;�����oh��m i?chz��b+3}�b�����, 
�E0���=�2MY�3����aR!w�F A��S��M��o��q4���+��o�M����a��F�$կ�#I?v�xƑ�>��"L$��J���QI� �y����PӁ��˳��w�w��џ�<f͞��>���wH䣄�=��'�g��ϛ���>�C}Ĕ�?���__���ώ���n�w���<��1�l�h*[.+[��CS9�{?'�A��O`j��[}�3�y�-�q��#)��1�1��]������ "�>�E2�M�oq>��W	�%ml�}����_���,Ϯ[Q������t��Q�ˌBqB�+/��TWO����)��r�����2�ֿP�<�vԭ�[!(�@"�~W31��T��g}�10�.�y$/�k�3����m�H���� �wW'���SD:VW��٤X�9Y����Z�L�>��]����U0N�����B��"�QG���ql/��F~�"	�i��b�ʠD�=�� ���˻�f��Y�Z��?j�Î��h�J�ZD��A�U�۹c�"�e���,�x4�<G��Etn.'���c8��S`�����=��p�ƴ�ފ$���Q`���׹�`���r���R��]Rz���ǀy����޵�?��F�֭]b�w��`����[^"f��ݔ�������r��ұ���>m_�˳��4Wy��@U�kÂ�Mѿl��]��:,M��8!���֖�tM��$?���$����>y���8Ċ��NDds)��7��������-Mkl�\�M�gk
��s����<�*J'>+�\��=P�<��;����7��@D"�o�Kj֣����R�ny�}ݔLgө��+����Wl_7�c��p��.��2�]����]����]�2�pH�f���9Yq5�n�@��)o]wp/���%�4?��7f9�w���N����aٽ�[H��=柢�@H��@:���`��{��F�.���'�񍏧�!C�5rm��������)W`�;��Q#3�j$O���k\W��NHU�28�v��1$􁨳�v�;���ﮝh�2��!堵ε�/���F1�ϩ�W�~}p� H�y���;ԫ1-�/�Ȕ�����c��z��!3��,�����%i���E_����Vd����( ;V��؊/�V��w��1̻���\�8:1;f�=����ρ�ry:�jV�������<�/�%Ӥ�4K�y����k�v��S|�|?���W�B�����'�1.�g!��E"egqF�e�����_�@�`L��������k��F�i�t�n���U��t��*j�s�F�Yd��]������N<]�=-L��F��ұz;Y�\�X. ���X�hE��,��yk��J��M�������- �
����X�a��;��jQ�8�Fw���i�E��:Z���q�d�.���F��mO�YZj���~�\@?H�����
�0�����P4�-?2�ζ)N��2E_r�E�A�#\EJ��7���y�@e.։L��.�
����X4�[?5����L�|�?�?�;:�nAd� � (���y6v\�������pQ����G��%.�+�����v<�#���ߍ���Zu;6��Fd8���o��_a\��`CճEE�=�]�$(W����x�+�=��~w;�C��X{m�i����VWc5t޴<��
�iL�E	e1I ��������wR�ҪE�X4����X��,��W8�V{��S��w���ͩsʺ�b�G�;K�8
X���,�3%�W�iI�E���b�f_������V�rlr�#0b$�ٍޯO�w�cvي�a����fr{-�bY]��,'g�у�[���oY��{|��/4����8�f5^>�Qq��Xò�{��v��r8�|Lh�xIx�G�QM��/[���7V�	�I�FyG��*����8��N�1��\�W
HPiC���hY���9�&z���t����̝1}0Fp̢4�\�7�eHǹ���kF5�t�ด��3�D�`y�~��ۮɌ���>Ɯv5�!�� �p���}�KnQ��f��&�2�i�>b޾�5s���'�&vu����8�'|A��*.�&�ۥ��kǛ;�K�HA�{����@�ϐo̪�෧Cֵ��O=v�?Z#;t�����z��fi�2l��W�������=�b2
�!6�����J�V7}��»W��{���
��A�m����ۖ��G�+(G���+g<d�:��=;�2�d�����)�ᣅ�0��{�d��0��IP���Ɇ����5����h��1Y�S�!)��ت́��y��1pg���i�-�*Ay��.�W�c��)5�����
%=��wHMCd1p�H��'/�����u}i�0b����q)�s���M^�D�fN�f!,Lfx�oB���$~�~�:m�!�������:�t���V%�A�	�WP�=Ҫ�O%WN��X�ڰq3��?b���9h���-��M�kl�G���b���,�~aWl9@�.ǸC�W=
]!�ˍ���"uS��'B�w�1�/(W��+�����Cf�7�� F
?�(J�c���b��c#qx+sӇBc�9XR=��J����H���c˯Wm���ݥ�V6��.��<��5ê_U�>{�&D�αՅ��U�.^���o�|Т�Y!�J��(jG�{ɘ��]��_�*�"�L���Knm������c���,�=k���Xh4��*g��f���YH�$��S*�y��M��E�I���|���݂��6e	R��>3���6G=�Q�ƨ�Մ�'P�5�}fo���$��۽i&l���-ͫ������c���=�g?4$]ݽ�ܪ��w�`�!�wu	�PΦ�骼'�!	�
�G�bC�XId��PI��dq��/շ_��8�ЀTVt\����X�0sp ��R��ʽ%�՞w]�N���߉����Yt�n��_���r�/��hT����#�V	�K�g�@�v���A����|��	6�Ikp;�[I������/x>D�e����[V�E'�g��Թ����Z��V<%�+�`���v~�I�|\5D��7e��H���(
C��K����C9�����zV�4�z��Y5IAG�NW�N͉���v��a��L��D�a�t�YIu	������Y�n7��������s	�׽�E�b;��^g��C�� �A�k���I��	ʴ4,;���y*��f'�h��k\���(�p�ΩIr%�z��	u��q�o4�s��Ê\��pV��T�菦|��]B��b|��Z�Zy���B&ۇ���r+J�Оv���ٕQ���o��=�9�O�d�������v���Tȼ<��J��	����h�?�C����"�N��5��m%d-��Sīk�w�MVU^G��#u	���I��Za���{�3w��(
���q]��R�<�w��ڲ��]�A�E�Q��V�%����E���i����E��G�7�m��KKx��#4�%T��9t�Q�s���V�'����Mj���oݥ_�%��W�w�4j�k�Q}�=�;�܍��h�=�ͬUT�"��#ް���aE�Fj��NgmL����k�	p`b�n׼�O��<Ĵ��?i���k����|����4�SB����c?��^�>RK1|��RY��1Z�2w�R1^�4�>D��|H�A�}�������i���5g�y�ד�+�?�������>06Κ+�6�d���H�U�S��en17�>	,�� �!�3˜�K��{y�~�5M�g���3��k�Q�}847P<�$����UF��V�T�g�C#K��;�'�W��A���B8�ޓ�6?%_���X��5"p�8l�
�S.�����f =8u)����C�C�;R�����vB�D�C�O�������'Rv��)x�;�P��d������p��=1}'�K)	5p���f#d����;��j��V�8���N���[c���M�Pd17(��m���3�<��r��<?�2�����IF�\��߭���!��7ޯB�#���x�7!)zƊs�����-+�f�9�Ys'p/5�;Y�yT$��1w� �T9�Q|"�⨃�����?#;���j5�)�Au��LE����eZ�c��zO�G9u�oaX��m[�h�[2l�Ɩt�$��U����ψB��AU)M�J�.>&s��R�c���5�	��Fq�y~�|۟w���~{m�.�����E�A$wpdA�U�5Fw��{%+_�_������r�����L����-��y������L��]Z�PRp�;����๋Jo
~)�?��/n!0B�9����h9�,{3n�[uh6<î�Yd�5�,3����K#EoD�U��Z6���h�<$�%�C�t �1զ)�,t�̊�e�w;m�5���T��_��.w�:���)W�d��#(Q�ܖ}�&u�?|��H���ʥ�Rl�l0n����2����L�żt%*s*0�£N��Q�؆1�Hň'�ë�d��$Tz��R��_;T1����~����cf��^a���Sa{�T�B�B�s�����U�Y�*+� )��R�G_C��C��F�G���s���ޕI�[<<�r�9
�C�� ���J��?��]1|�qF���%��0�v�C�sԲ뉷�K��"u�ħ�_����ܱU�6nVAnM��S>+U��. Q�T���r`�}G[e.W�d� /ɇhP�� �J�8XډQT[Y�����zXh�X���v�n{�� ��?��P	7a�C�M���p�#�|�g"���/�&�:s��d��ՠ�>��!����t=�Cb��ݞ�.�]�7�;���&���d��&~�.u�t��"�)���'7�4�]�\�1�'���h�hnG�UHL�'(���x����;�
������˻ían��<��-W[��K�����.�]������㼏���v��.��y�b��z���)��25G�[H� D���I&2���r0Zg����҄Cd+d�Sme:>�!�N�n��Sd(��?%�V��<������`90xO5�]�\��VmWL���Ԩ#Yd�=�XZ�.E�7yց��%fm6L<w1�R�%?�����Ȏ\�y�T�Uv�]�a��R]�m����o9�L�9[
fu�d| x������K��e4y��tP���t�����6�9�5~ǚ�#��T��[���M�O;�Xfa��#c�W?�ă=���p�#�O>��xs��]P�<����BtJU��ȥ����
��?������2w�6_�C1bI	@1�ga<Y��D{E����ҬѢkY�Dk���v��Nt�?��?ُǧ��	5��%�}1�%���x����P> �NX1�-�o�ZD�}U����Mu}ip��4�>r��hƝo3�dQw�Ǖ��F!S��w,��P4����F���3]�'�Nn�������n�4�����Ę���4�JhfLK�OR+,IGc�9���vʹ.�*"�P��_�>�R�0F^������H�6_�}�~[�K蟬�pB}?6�3�U
�TO/$�*�ͬ��#-�}@�V1 ͅ���� }����p��9��>�慽t#��=�s�'�Q唂Yj�gP���<Xd9�����$&��rPxx�[��I��0�r��}�R�r)^��<8����\�c�)ڊ�h+!����v����n�QX��	m�>�(�V�Q�	�zH]����&�0F&�z�Atzr�\9�V.0�!�c�f��n#q�Q'����}ZX����IF��FT2ya5E�_�p�0�[ƹ�&k�����"!�31<�ɣ5�ea�.��/�*�qn�%�׶+א�%
+�DU��F9bJ�ߓ⸸�t�M���g�-K���c��kO՛� �1���t�a�@����0��9hW�Egk��:�������)APZn���Lw6�ԣK��B�.�q����Iy���7	k���.y�~�7Vg�
�}��R��9a���njZL�U%6�]Ay�h��-f!a\�>f� �m��:1hCXɎ�-�Gt+(S���v0!H0(�;�iWj
�
�=j�-��Q�ϖRF]:���Z'>j�nFl�-�ļ��Z�Ci�i
���?���>s�)��ݬ�).fkq%����9M̪�{�K��sbz[&��f�au�r��)�34���dL����>ځ�(�7��Uϣw�-()hK�9+��^��ץSz�@���ҩ4��^_��-FpU�r��=C]�<�TY<q<�����kO�%|c6���������(��sO�r��i����D��N�Pӆ����d���
�a�蛰ć�|&x~���n�Wk�ĢIO峬�����Ŝ2�b��F�O^�^�(R'��
�}�r�E����:H13��D������56�DW[�1�QȀ�槡�]�K0���jsi�������v�O[{�X��~�HzG_`i]�/A��)�J�דL��W��������D�M���\����D�.#��5��^5��MFX�K���P������0� ̇�d�ה�V���?�Ӌ�P�mlo�>��(�<�+C�(��!u� ̅(��G�Pc�
�=,�.�sĊi�,f���vc0��DR���CB~䏉�r*�l���H �������~��`�����T��ؔ#����z�>�P�V!e}�������/����9��J�,a:+��$P���e�՟b��1���a��>��]��lQ��P��,��Py�?�Sa�VZ���k�J+����-�5���@�slxZ�|¥<݁g9}�K�c�uډ�+E@��<.��bDc�t��.�0�F�jN�&O �'<!��98{Ի�õ��ܫ�@��&vMH��ܛ ��XB���fk5��g�U1����Q����3v���.e��	����Ei�����4yb�_���"�-n&p�U��}�j�g�3e���U.���0Q�%j�g���y,�pP]��1�>�0�I(�C�hv�hRK��#�vc�?l@��!J�APFw廓`ԠI�n�/K��{A���n�&��ub������wT������ֱG�?�7��կ��Vg-a�����".F�|#� �������-�TZƒ�"�t/f�OP��:N����oqr���kA�'���@�>��;̮��\+c�35��-I�P�A%���'��(��bA�886܋�@0���ũ����SV�:�w����-�}1�O'��D���E�P��aս���j��P���W�����*F�ʉ'֩&�>$�B�.���c�5|��	lK��ɩ�1ꄪ�,��&-Cb��]4�BB�|�`�vfQ�Ң��#�o�c	0Ks�ЌW�_���f��U)p�>�m-2��-ϴ"�?|�7��\�&�σ�Q�S7z�~�E{�r+9M�W��������pvZ��qS���G���x7�1�<8�h!��^�C[��ԫ�'F`�r>�����W����:����IvK�8�/�M�Ű�//�wȲ����n#��/WkCՆ���g�"���ܖ�@�7��?cO8i�9�V���XB(˷`(�x<�B��[>�@������ď��h��\�tN�s����R���~C��ꏨ�f� }NsH��R�D���X)�8�S�aU�,6~G≺���
�VcS���j��Yl�ip"��	i��N�	vq��ӧ&�|N.����#io�f�`ͽN�i��]l%����j#���0�\�+fwO� �����#����m?Z%�Ն�E�!�1JZ���7�b�t��O��
S�Bq9����o�
4���Mj� JY]���KT:-;�AH:��[��Wa�Q��	�_,p���N��/<Ss�꼢]$��֓]�r�����	E��X�Y4w�g�svœK�c��3m��g�Bj��jdG^�t�>C��ik/���w�O��i���Ʌ�����9�����՛ ~ӛ 0��$��K�G�yt�z7Ƕ���������E�5 �U��ң��ԓ8�-��O���/���Cq��r\�v�U�FC�ޢ��9F�-�
8z�o/�m�����m���V:{�a�\��NPC4>�~T��,A~D�����O2�E��9D/.�(��N�`n����=����ep�(s�dyy�ԉ�Ґ�ſ�1'WrSDs���K(Nb��tzg>���_�a$[BL^��onWo�}� &��zê>�e+B�Y���,Z�d-Z�d�+��7Χ��N�BӪ��x�N~^���p��&�9�h��Ҏ�?�6��f� ��n�G�2�_�]A6�P�M���T�.e�$��H�J��k��~���}y,�ɚ���}�Ǒ|�_��Z��y�����x�Ix��O��ة96Ŧw�S�n�q���r=�E!�
���h�3T��:�aMC�̂��ܪ�$�%�b�*���R󢺾{�2~�0����N��� pѣhx�d����v������T�����==��z��*��u`������M��=v�J;��f$|�ci����
X��yu"2c�O3U�M~w�W>����7V�J�����eW���"ܚ�u��"���ۼ�\�.��-I���Ɠ�۷���T�Zs��� Ҙ�ߙ*Ą(��cr[�e��O9�e��	4�:�ϙ�������.-${^�݁����ԭ��(��~�����4�'NJ�
u��bQVyń	�z��k��ג���(L�}����Wb�^��Ko����i�R�6������u8�~K�&�Gվ��n{k�Pݛ��!�����ޙKY+e>{��.��9\��G�J.(��k��֚�0[�Z|�x�be�U]��o�ؖZl�P�e*<.PS�Z�
����+-�R=��_��V�� \���k��B�Z|�)��c��.�3U�na�(�, �T��Jn�z�,o?k�R�㫒b.O��;$�d�w[E.�A�yG?)���?HĿ}�?�Q��P1������22��	�.���-	I��Bieq������;��
�����+��a�݂2=) ���h��Ҫk���Q _����Ϩ47wi��,��V�2�x�Z�E�&��V�
&���u�-|�A��Vx���{���#,��3�(�!uI��RӐn������s�R>*�ʁ�,�Ӽχ�m&��$$᠆��AQs6SG0�("U�rdg���g �v-`R�pB��2��<EU�t�� ��ی�|�~�'�W(��M��3����Q�cןf�!���Fd�~�	�w"Xmy޳�mڜOO>%��<���r:}#ש6�C��b�_�V�R�H��ɜ����2Zi˳v���͌�K;��+���^��`.�{0l��I-9B���u$�:�CΨ�6�;���������51�X�g���l�I��	f�0�4�B�K���O��;W��R���m��nB�\vYQӏ�����-��_�j��$-|,�M�o�m��D��+X$��TBE!5
H��0�pqZ��з�n��D�V#l�6R�
 51M=�XL��p���H�ІE`�������d�H�q�;�'�~3-�&�N"A��k#���tdړ��L˟��sJE����P[����<n1��,�-��6�3]>ޤ�0�<�����E�vc��ז�t"5�V��ք*��x�X�À��7R�;#��b����8��2�hUoz>����ͤ ������EI��z�z�=�2��[�{������k�}������ǿ��_�O��_	�~�4�������^��#����M��P�y�����Pr�:��o&3�0�O�>����SS��|�n��X�1@�p�h��k#F�l~�/��eʯf嫯<�L���6x�̰c�*^Hq&���5��57��T��Қ��B�B��(�1�J�^�ӧZ�	��ô��V��6j��t|d]Y�A��43�p�z+�L3�V?|�u(Nl���H����$/������P%��d���;`bsp����T]1���-��aI�������S
�8�^Ej),�<5x���ja�0Y�"9d�dى$ye�Zp��_�&��H_R	]���_�u�Έ��,�fa�N�h����7����\N��A�D��KLr������g�o�D�fEƐ�|����|�oi\���D	��w+%�[~��鐃B`��.�-��Þhj��Ǩ��<A��qX��"�D9�e6�~���\$K����ꘌ��J�UuI2j`�OV���I4�pnv���	�w5bЉ��\5�ݐ�rykS�¾�%�1����V&����?�cd���S�+,��h�d��f��3���/2uR4���ew�xm�Q'��Y=EB�>s_r�"� �&;t�`�@�����7Aydϐ�ĮT#���m���^����9��`�r�L�;P��59}p=|R4�����*tҒ��햎���BF	u�塑�ik>A�j��3y}y��j^ 0�横��qj����A������U�OQ���ȳ���o��M��"�fO����H	*�g�lRL�^;��l�t�$$pmZ&wAj地�X*\���}u��u(k�+V��.F���H��E��-��	���;v�}� ����<�CP�K��|[�[�>wp��tfH�;����A9Q���Qӭ�������Ҩ骓H�,�b���-^�俬0C��OG�n�vx
��F#^E��L(�?���n\���?oc�|�qA��d|6.�!rFx髌�q���5y����ŘW���\;���`�I�3w%}b|"P�-�%�N}Y���`�)���6y6�'�\B3��R�/1�~k��/�$b���M-������wp��/!��[���5�V�/�"l?lO�qqa�x����V�K<ŀ�L��1�kq	�jBV#ʴD6+�U]I"E�W˗�Xl������4ڿ oW�E�8\f�=Kx����g��Y���,,͡�7�ګL��E���}OƔ�h�}H-�C r�x��Xyg[�����"�����"�r�Rt�xo#cCh}9���y)��e��.�2z�b���ٳ�5�,�^32�2�qI,:0������Ias��t@|U;jw��6r��N�`,N��f����<�V�<_���o7d�X���
G�&��usAUJz���Q���UꦢpU���伤��<z�Kn!�2[����^ I�`��Fע[7��1�\�U��0�ݙL��l���KH��M� &5Iր�4r��[P̫��nh%��f��t4B�w���\|�(9l�amp��W���~�[�&�ʥ:�(�ڝ�$��<Z��F�oD,��Bu����C>�%��"���Q�K!ƪ��T�r)J7�B>��V��ʋ1h��m���*��i��?�U�2�H��Z>!Kg篧٥� ����30�0����Z稣��V��mX�/�����*�1ȕ%���\[W}40�B[Zl:B�Q:��Z��t)����K��[IN̡[ޥ��b<>�������.�����V�Ń�u�r�i|c���O$㡤���{Σ|�Ic��5;FK&=�R�{%�wڈ���-c3& �r�-���a8���{�r�:���h�[or|l[��(MPf�3X2�E�8/'2��4֘��u��oWwyQ��̵���'��)�������7=�G��	�@'8�Mv�=������;E���s(����%��e�{f������k얇&�~�Q�'*�t�".��B` �?T�p�!w{NOL��.���M'��Qg���$|�$�L��I��ᎾLn9�J����6g�fMd�ݥzw�3F�傷�&���U�@!���I��6a���2��~E�&�<D�hk�:��G���	�����0��9T���^�2� 7p%�+Vk����{�>�~�D��T1N��C���Xs�����`we���gR���� ��2�����Ab@�>~)Y_���?��"K��W�ϓ��	���p���lX�	����iG��)�qLm���A��]0Z��\�����K8�\�SS����q&e<T6��I:��3���+a�@'���g�4�㍚#8d��B�I���m���D3u��ԫ(�ޡ���a�}���4�+��~-)��p�e��1+#G�!��;�x��Ѐ!P)Ԅ*)*R%FE�<{B�Vv(T����Py�N�Y��&��w��i-E�F�����./�J���,B�i��$�m�N߮�ňe>�̈���F.�AW�����xwR7ƪ���T�%6~C�v�?����(q�y)�E�@��X�I���ǎ2u�*���®�^%h�~*F���4��1�m��b��*_�V���&w�����ޙ6��������,�w�'��I=���jm�&mx=K�I�m�(*0��Z��|�ƨ������.���`Ȱ^�h*����J���{��ͨ�P�1��py��О5�/֘�j�sc�MMB���*VBC	��~G�f*�Є�>C�9*mg0d�%�r+���Br�\Ԥ;����!�w�ǁ�%g����@tBK��44Z]ܧDX��?=��������Պ��IN5�7�H\�9c�(���a$� �+djڶ�tW�wM�[p�/�N�ύ�_$���|mz��=�J+n<�a�NTo4P�i`�T���v��-�R坂6��Yh��]��M�
-I����L�"ſ6$�J���ߥ��G^�>��(��b�^�b�tNH���t�U*�IXF�'��������0\0�9G��<FoF%9G�І7)��`��6�7���Mg�)b%��֙�L1*3�6��֤��s����(5e���X8�}h����ꥉ��}���|��N�]�'�Q��f!0��'�sE�����˅SR� \�Ki�t�j�
H`�'��F�Q�j�(����IG� �XB��(�<�Er5^ ��Ag!ﻞ4�a�����z!ME�M��Et7�ݍ,������z���t1�F]������sJ~(�ot,@�E���4�D�c�����!���T�'���x]��&#2D�[i4����p�+<>��9��a�@�$��×Wq��axQ=k�JQfCבu
�)� +�6�<]�QE;��V)>}�Q��12���%H�lB[W��D����@Θ�1QŒ�]��}W~�7�X��ݞ6�<N:���k�E�!�^��`�]���>��gp,|���τOS���s��&�������p���k�8�����F��aK��;���']�76��ṡ������C��xgi=%�d�5j�~�Nv̂=>m7��d{$c�7���S�㞥.��֠���Ck4�!)���;�O����"VƵ�)��	�%`�-d�s�_s��}H}f3����,q�:$W窟l��=b�y��]؂���|��a���1+z1́.�cJQn5�؛����(��9#�ڤ`�I�yE��䠟R�$[k׶)އ�UoesZ�	&/J;��=T�r��K�\HI�vɓ�.ӬX�Nz�ԣ�Y���Q�BA}w��l��{I(V��^���C�~�
L.t���'+�����֏x7�W���(N�[1:�=@����V���C���f�ꨲ-�}${�����/�Ɉ�������+!}	�}L���F����k.8��z���ㅁ�"�x��.�殠�xw�'���P�Jw�@��T��v�A"�r�یǒ�
ǖ�%�+��(Ix�t�Ƚ	8�l2Q�@M&�Mjv�b��W�9H�����h��|��8���r�� �Y#�f��� c�����b' �#�4EFr-�.���q9���?�ɹmϻ�?����F!P�����^h�B�J��6�a���"QW�獧E(�	ۂ��ol-��O�������*��Xi��Ȍv(��8�@���R�kW��R O�Ѱ�2+��¸�U�ѭ��>��ķDcr��?U�WGM��BE��hC)2S_G䦴���1@f���!�9�Z��a�3��w�1p0<9B 5lʏ�.�q��0oW�
;�����h��k�.��_S����sv(ty����f��i�U�dz^��������7������tz���Nn'pQN�#N��f�)�)��z��ety*���Q�%����n�BX�م\-�Թ}F1Ոc�P���xq�1�v����q�8�?�^&9vC����0�jk��olR)���b�ʪ��Lr_�'�˦��%��;�D^�����Ӂ�p����E!�p��f%z�^O��@oN�Y�/���݀�*��x#0�i�#H}B&���t�~<`n(�ǢpF�G�7{`��.��ΦinO�OZa"�x���r]�5��iE�cl:��I+`a�O(�:��sq�߬���ۀE+�\�5Q��"c[�F�ɘ�Y�W���¾0�r�N��X.��;��z�KN���pj$ױ��r�_� QU9�ʸ�reu���Fk4{�ɗ[	|�3�_�} ��{8`�B�r+ɫ��h��R�W�"q9�}��|��dFؘ
��<-f��.���n���|󜥐q&'NL�Y�ꅻ/������Bf�����4�c�P� X�v���Cj��
�����K�M<0���-P��ژ����y���2��K�$ﯰ��,/m��
EvE����CS��蔇6:W����5x<|�^E3�ۭ�g�H�t�)c �az�<`�/��;x����/��x?�����d�p����X�u�+��WDG8���=�iQS۞L�2�tȄ�Jl^s�ԓ/K=q��s�x��3J%��GH=V�I�A#�������Hj���C� e5��zH�\\Vſ^��?�^��V!�L����Q����E^���ÿN���Ok�a�h��+�6���h�E{ff�&b|�zi%�*����}���~�� �v��Q����TÏރ2(��7՟"%tD>����?�ѓ[�cp��@-�QS)t��SZ]P�&�74K���G/e��nｄ��4v�������*a;����:����y^D�,��~���IW��J&\'-�;\�Ͳa1�iN�s,U�/��j7�� >ٕ(�+QG��,�Ii/�:�A`렁�i�#`	q�/� W8'��(^:��Ҟ�X� �kTai��$e��*�77����ꆘ%u��np-V&���<���c�)��k~�Cn��C�U�s⹶^�V�i�X~������֓]1���|�a&�1dK��V��*s���N~�C1=o۴�	P�މth���� �f�%�p�I��ۤx���5����m�Y"K�t&Rڀ�~
�:���Ȼ5)X���T�W�!��\7��`���L��>�|MQ�f�1�����	�OQ�%>@�`jt&�_�YQ_3��
2��~Y�?�0`.�_3jq.����¼V���u�H�g�I�w>��cj��rm�h=4��"�܀��Z��.�}2b8�;�c��W�s�bZW��87�tR}?/[�2�4鼠�KnP4H,�r�a�+��E���4�}z\�Ӽ?��. P��'M�c��_����b�X�5����qx��$�7��6���	,�|���
af���7OH6/Oƫ��+p���h��Cs�|�?46�J�2�����	��x��GR5 _R�&�L.^�I 3�g)����|�m�����Л���DV~CoH�c��N+㕑{�&�.�Ը�ȫ����o1����0�Zj���o��H�2Ŕ�����#j��H��T1h���*K=���ܸ��rd�~+��U�}��O�G4^�)��=OG��,+�&:ƺBx��!U�tn��nL��6�\��5�����xP��cQ!�>l?�����D����~�8
ZY�;`�ƭ��=�?����hs��s�:�B"@���k�-[�z��C�)�7r�0,�ʨ��O�:2<��ϛ��8������e�qPIrh�a���I��+��P]�DK���`�4�������G�L>߱�@�Q� ��if�@�T>��\�fxYL��(��B��C��
�}�H]��Ӯ���1�4d�1�r������S����<�&�S�cU�����d��z���n��.�u3��%��4�]CK��5��[�P�5=�i���(�������X ��e
��6v��[�e\nb�����d�X���%T��7vY_ү��}w|��A[e�ߡ��#ΞF�V��K	}���:������e���s��x��������Y�=ޟ������Zʦk�%0JV�M��2�i;}����Kj��۵��b��������~���'�%��#��#�ж��<�->"l���}��#�d[|D�Kh��vi��?��}%G6m|�-�ؚ���6���m
��4�pͧV�2���vR�{ގ�����?�v��gގ�����ڇߎ������]Z��(���cvY����<�<�.�Bퟹx�߸����䇱	ҡ�(<�z����{w��7�������ߙ���wzk|�������[��ﳭ���MG�%NÏ٥ ���%�Ħ��n]
�[i��c��!ބf��sg3u���өW@B8r�R��@*���i�1��-��>���y28��L}�G��*���-��ہ6  XOӛ�V��l'DPb�f6�^�4x������Ւ��=2�Y�{� %���Y��b4�#��\[	�z�b�LW���2=�s����v;�W�Y`o���_"ˤn�w}L���xY�8�x�f���ӱ�C�l�u3~�:����������l,�G%�K1,��H���R���Ϸ1c(Y�� ��-��gj�ʡ]�gm[��Y��,p�\3���� d�!!d��CqH�fd߇n&�����a@�CR�TN~?�sLK#�m�f�#Zn2s�����H����5EޢI��O�e����ٌ�>¯G=�C>$�qɆ� #���C�7#C��� A� x�]r��]��k�a��vˮ)�>g�9[���Bz���\�� j�R�E��ϓٌ�xs��&hW ����V:d(�e�� uM?T�t��b�o9�Su�tXY~ /�o��!��
40�U��ދ&&K����_�3u�G�Քߐ����o����Dp����,��	>�>eI���%垦�m��$)�y+�Ѝ\P������Z�q%�T�����Iؤ�gG��}	8�dT&U��p��bf�7�p��9��m�ω�B<+����I=��a�$��~��ï�ar�:��7d\�c�lBc�E��]�w��0wF1����J�8��3-0�(�E�����@9��7�#�_n�����*7}X��M1�j�&m8��Ѥ��_Py�s�2M|vW#�sӎє�a�`���E"�y�/���,�� ���L�s,�ڐ��ua���nH�ۀ�qFb[�{_�f�s�F�/K��7iW(�0��b7�v9��@�C����� ��-GS�Ȑ���M_*�wb�F������_C-�i6��b;����/Bc���e����IU�E1��&�p�q�0��ͤ�d�c��]%�UR�g����7���E���I����W3�F��$��~d]���uI&OB�h�\����6p�_q�$�GB!;؇`�V���&KȰ�_l����	�&eM���?��z!Í�kP����j����zv�^1D��i��?3c(�!�goƈ}f�����J?�6�)1
��C����H�ӊG�
�ԟ&.�J��Y#n�!T�܅f�5��:�;T�	���'����A���Z��i^G�H؃n�E���,/VG2%��q;b�3�H��I���~B~a�Q�S[�R�-<_���@�i��[��O
�U� <��#����m �*����4�i)� E���Y�d�|Y3*�I��Zެ���c%�*P�%��]u�]7�۾s�mns;'i���h��TD��m�U(m���y�M�B����($����=���<�<�9�v�5��0��:��3��%m�\#V��	�� �]��mx��$�������y�gؑ�����	����a�UF�mv�����f�M��\+_��5{l�k#gu������2�awL�`5�-E��Ӧl�z���ov�K�ru���5�s�R+e��wK�)m�7������C�~�;����/0��2�i����J�4B��\vb]��G>����Be�#F|�TG��watG���Y�S�1�p�q PRl��d9g2��J�d��&�Bm�]�,�ߔ�ojl;֥V�9;f�oEҽa�
:g�2�(�x�+����Y�z���W�=Ta� �~H�R�0��0X_j�˪y��:D�s��b­ѧ4��6ϵ~�#j�c\���q�A���*�-�X$�3��- O�`SZ������g��\���G�[�0��G�ﾍ���Q�@�vg���!��xݜ�o��d!���[m�����U;��`���>B�а�^J����^��"������Ӗԯd|�^�%�q?�آ|	�+�䰬���|,���vz��U%�ʿ�MwS����7����Z*��,�|��C@�SxW�4�f�%6ߊOF�Y�)5W�Zx��ŬW�DxyKA���&�M�Ģ��O����D2���e�C᭰t�[����N�H�rm��04:L�9#�D[2@��<�~��Um�ʋw�&�e���Q6_A�a��&v���Â�Ǟ��I�햭�7��BI�Y~x�1إ�sZw -֏��ok�G@7_I�/��I�"�O���-�}����+�W���wR}v�o'�*R����ھ�C�G�4F-GvU�lB�Êy�K-�*cb�T�S��Z0hM��a�s,��+���������0��|�s������cF��'��f�Qj�V������@�RUk��H^_����&3Q�J�t��=�+4jݽfC<l{L*��!�)� �0�}B����`g�Չ>�����`�߭��%V��8Vo�ח�ퟤ���	�ɏt4��Y'_�����%�`%���ܨ�p��W���L�a��[��ˍV*�ظ������'�)XػG�F�T�]�F����$��������GH�����rEf�ڶegV {�t(�0�C�lMϨĉ�_��tW�X;Ŕ�eΝ�W�T�U�c�-��J2���އ�~�6~SGO�ݻ�x��\��B)�ɶ��y~�~l��o1*���J-$W���V��BQ�
�K���ȑ�c�}qL_��J�E��G���7rq��pmNi7pѮ��'�e���4�0��t��;ρ��x���h�v#���Q���`*�¥'���b��].�7e�$P#@��U���:1\}��T�j0�ow�Hk2�������Pw�@N��7��a��;Wor��qQԛ�뇟?���@���y�RM��e"X`F1TatH%�鑿$�0d���WeT��6��|R����uv*?G_/�W�&������?5�񍋠��3.�fE.��Ӱ�o���1��1�ی���:��n��H=�\��g����X��=��'[�!�t̶G���H�G�<� 7��C孾����W����VX���� ��d_�m�C���Q_������FcR�Q����T�JVG;%���K��x���U��O��������rG6� �����2i�����ATn�i�t�������:0�l  "ݹ�NLar��/�������4�z�M��Nj���f�=��r6���ӊH8x^d����A�X���U!�
�Q���cB]1ĕ������s��;��E�?�S'
���s�A���c�W�g"R.U����9O����x���,��lI�mJ��0����0 %G� |�wu(�ZH�$�X�l}��w+�k)	�<JWϢ��ި��V��gp|�OU KYy-�@u|���Ȇ�cCߧ�W�/h��|#��~��;:]u�~�X��g'�+��K�An5�ꏣ�2^?a�e^��<�хo�ǉ��k<˼�M�b��LJ��{/���?C|�$�<�+�(�%��C��gV���>����q	��,`1����j����,j�̈́T���d��)��,�
v�,���f�O͔O^+�����_{?��2j7̕����%^��]S���Iͫ�⥊�rI�9@F^?K"���^aN�ZU�T���p��?n��<��o��G�����K"ј;4���L'�6 �~�?�ɯA�Q����I�Al�������M[=
�^�ay�����~0q~��m�!^D]|~@�ܟ�؜t���.�,Z�j�]�-�+w����������R��Wd��N��Z>Q�a<�j(⠈K	_��K&-�F#�m���Gs	�([��)>����}��3�&M�㛰S��v�Q(�23���[9�WQ�Q���)bUO(�4��_��1+��\��Dy�*���oq��R@iy����BY��j�ii&�IIk�Z�4j����.hU�q�K8�·{K�]+�S~ր�#2)�|��\+���ª�S=�K	�8�����n�}��0�zXc�7��l��
��׌��e���vSx<N>��t~=�A�K�u�n~:�nҵO-�)m�;��$;�3~�H{R����U|�%���U,?��[K�WM(�7���c���{��hu����!J�T�����/��~�P��5}E�� ���u�ņ�ae���ɷ~GoA+k�RW��ތ�'���oq��k�gj��$�u�:��gI��9���/�'��ȏ.N���8�?~y������@���C��q���/燦��Q������������$��������!�A�+�������s�������K��w��闭��	�Q��lh���2|��?b^bܹ؎��ܯ_[�9,����?=�������Ǔ�A�/�34�������������!�����8��=e���|����7�g�������-J��o�?qX������!�e�0�?<��,����� ��rG�eC�_ޫ���C��E�?}x��c��������n���?{h�?3�g�������!��	�a��3���YC����>����Cпז���џn��o��k0�����!��<�O�=�C�_u�Wϥk�2�5��z���e���.=����������u�E�~ب*iCӿd�����_H�_{����@�[���N1��/Bf�y���B����h��~�����Ӈ�ߞ�94�;����M�����%�����f���/�������a�x��Y8�'�?�� �o�1��v������8���mH�O����7'��`���N[�Z��B�C������S���D�	ǰ��14���S��nx����7&�����?,��K���!��8��?i��l�V�_c1����6xg�j&���V?���������w��ؠ�*�_�:�0hj�1}J��>U14>�����ѷ�����f�KS;�E���v�	�;K`π�Mʚj�CcE:j�?>��� �ٗ�m�4����_]@����]�
l��s�Ql�����{}�����ZȌ��.�ח���驇�z�B�X��<���LC���(iy��Bp��b������4��B[@P��y��}th����VG�,CAL�vEc,kA�{g�����`����nqs��%_����ܟ&���9�)�[�37��O�wY#6��W�f�]N��F��5�:xq?0��=�n����i��ʙ�߱�dg������1��N|7:n���\=ƴ�$=�V����ܕ��!�y/�1���ނ��ٻ�a~-�_�
_�ʌ �������OvF�t�\�㪁Z�mC�X�%s��������_�ۗ�B<�J����0�&���=	��O� ���?u���������>O��	�l���R�A���!��l��oܡm�x8�Wz�|���D��J���-�m�������qM���'�~�AJ�ݘ�]jֶ��I�RK�}���c�#��5�*���2��'�Ec�7��<��#��ϋ����9�$��.��L�/ƅ�`�3)4gm��wZ��`���mt^X�ySF��wci�XuD�q|`\)2���|`"�X�E�P_�.���~�7�6:�ƒѿ��|����)|M�
�3�a8�?l��b\�����7�Et˶EVU��)P�|���CPe�gȃ�CLCÃO@y��}+���W�lVG���v�W�Q_���F���L>I���Rif���o�����|yuN���6��;�-�7�����u���j�N��z �Jsⱷq�[�����j�_ͩϐ���HC��?4����o���B"RT���Ь��J�,�O���~2�.cO���x�C�������l���zyQ&�1�G1	a�dq�«��Y��՗s�f<w�«#�ڂ0bƀ�e�!>�ܨ�$�G<��qNX�B%\]��'��$��ר��fC]w��|;ߘ9�S�7���xI��C��x�"W��\�i>4�x:�s{�Y��z�Vb����%�κÆ�X��߰O��4��Ao��`]���?=b!&ԻRDi+P�ܝ!4+c��Â�`��W��� 퀋pe��k�+8igs��8�ߝ?�.�	�(�vH;��B����V��vR5�f�g�g� 3k+<j�l���̈́iũ��1����ym���q7�t
N�����~|r�~��Z8�q�P�A� ����$�w]^�?�s��o~��H���L<N�N��oIx�zK�c�ylRd�N����H�6�'^����<5I|�[㱅���׻�ͪy������!�H@��������B�8�����8����s�Yu�R������l�\�7
��X��S�������	��av(�V�Z`�n!J��ʄ/C��X,��-|�Xf�d�O����2 20���o�p�+�=�ᰗh8�%r����+c�k�3a�=cuǎD}�w;�0�)㲽 �����#����N�8����C��O��ט���D��|&��_�w)y=����p��\�	�.�M[wۅ�cO�p_��F�kC8<1g���A�
	,�7��&����n�U�}���(�����~�!$��/���ngv$X=[����ڲ���V��G��r3���W"���̐�cŃ�IA'������7xn���V�D���o�C�R���d�_n���x���F���l���w4<`�v��^jB%��>L�]GZ.9�V��fj�)*�;�aF��9.����r:s�7*{;�M����.��-/6G5��x1Q#��%Ҏ���)�T>� �=Y@�J��(˳��W��c�<w�$L
?]�4���P�~��b�Bﴇ��+Ũ2y�Y*)"@(B��`?�뭘K�!�MI4K�b�����JB��!C.3�%p��2H�<�\���rIQ�D��PtG��a��������:��n��
�������}�/;5���Tj�j���E{�Lռ�\k���=v����Zz5���-zWbϠ�?&3qW�	��"�y�ٕʍ tH�-�L�_L�K!0���BB��>M������ES��6u�֌o{e��@C[���م�x��/�.�{��J�5�!���r!���!?���疵v�����*���v����'� ��{� Wm��������x��h�RV�2�
3NC0",�ԇ#	sU:�V�)��$ �Ds��8���{wm_�h���l-1����Aiy��K��-2^	��]io��[i&��sFʪt�o�8)�(%�$�y"�H����u�@��K(��h�j~�������)�@�2���H��P [[�Wq���w���<=�GZ�tL)z�<��1�M�_�Ҕ���^�n:�	` Wp��l��3���dem���M��<���C[�Mw�W�����T�i֑�=�)W�k�jo �
:�,E�$�K>(KVG=�ු��i�[x���6=ܙ.�S����l5Y����,��(ݛ�Zb����{��%g��_�p.����%��*��K��4/�ț�����X0�g� �kZ�D +�����/��_{���S^,C�݈)��-��~m�Un�xKc{�m1�p�o��9�?�����Kb�r\���\��O�p�N��(�=*`j�^�t�QY#�7�j��[~i�!H�S_�5@����I�2
y�	#{1ѩuL�x�=�D�䢘O��nʅ!m�ւi���3�V����. �m�W���Ar�4c�4L*^&ʟ�D��W���(��U�)۱���	1�8��D Dٞ��65�e?��'L��t�x�9H��!�?�����jZ�$*�oz6N���n��$*r)ٞ�̄��FU�wݲ��[�E���ƭ�?�Qm1���Ke�4��{I�7��f���nS���l������]���f���|��/ee�6��h�u��h��h��q����������7Ow9����܃���Nw�1�f[�5E�'=���k��� ��	1Zŗ ��n`	��g�r0ʐi;H@�F��bJ�G��fM��F�ip�e���4���&�� �q�P^�=s�:�I���Q v�������uz2��EeU=�R�?��E9��Rw��ʗ5��Ԃ�P��{N�S�7/%Y�V�B� V��%��0�By�C�q���cp?m�v9�=d�����$�2萖�ӂ|{/BbٍM��}'h��K{��PLc.��m�*��P��yE/���7\i`��̂�\�#�i!H}���%[��(� �z�(�>(ӨhT���n����8��O�Oj��L�nR�%���j���^�<�#����>�p��&|����ԫ�h�'��7s)ٷ�|	��� ��� yJ��[91S��4����ƹs�4-H� ��}�	���;�6Pd)�K! C��O����I�<Y����K��X̰gV����F<W_�)�y ���`S�:�I���:�0��é���	��E�x�(���t;�r��n$�oS?@  6m��%z	�7��Hř������C�5�Z4��)���q�u�c'�����J��V�PCڕͧ�.�Vx�@��u�2�M��JmoBl'�W[���S�O������B:@�J�u�"ß�ө�R
]*
����('P@�ш�oGa	���C��zk�6yf�[^/���P���	�vO���3�T_�8�o������f�q�T�<�&⦙V�����s'?�s��<5*�S���gf��`byu!����WL�S���zyf�(�E��x�����zf���8,�F��%�v�o�]�#����sLn �5[3.ؙ.Ar�0c$Q��E w���`�ؚH���[�*�ʚ'9��(B��4�m;*�Z���<3�o�&r��m�s�37���ݯr|=���of�|W�<�ȋ��&�+d��1q��@���3�u-e�L%	�F+�iZ��:v�q@���Tr�:��}-����| �\�7r�S
b|c��|��[3��(L#�m;�1��o5���̔� ������8K�\��?7��u��َK`�bؗ�!R�L��V/���tД�v
R��;����4z���sv�4�+�P�mOm)�f�1�;��Ȏ����p���L��������F����|�F���{?��[�K�&��w� �~��i���^~c?-�8�4ݹ��/>�Z\LJ-�:��O�|�ٖ���[�S���e�AW�H��ܡ+Aͫ2i�\��b��B�f̯06�fS)��6.M�������K���@���'��{���L�g��"�o���̝��?��ȷ	5��=�������xSX�*�U��j�##�	t�L�q�b��_��� �������Iw8�M�.�e&���\�6��
 ����ɇ�Y�3#��v�[:�o3��a�`���8E����P�I�+S]:��0���s�o�3榟im]�*���(�im��ᶊA@.���;d�Q��O�䚙�>3p=�q�~��Ǡ���D���N0�u�Y��[�ם8��_J੺��E�cR�J��i��r>�~��7Cy��s��խ�W���[�L�YK����Z&6]!��e�-��������#S�<��ێ�٢����3�m�l��w����vx�c�%&CYR��3�FG���Y	­�!�az�N�k�:#����[U4H��mv�B2��e�.��������	{�!�v����=Qz�8d=���?z)ʽ�+fS���O�u�AcW���%u��4���j>hr緈�Ƕ�n��������6�ay,΁OA�y��V���g!|§>��)§���Y���Y	�K�s)|.�O04�����p���U�N���"���.�;�+��!�3�P��yN��vz]<���l��t�#�bރ	x4�P��v��E$�����Q~�Vge����ϕ׶������D��W��S����FlVL��0UP;L�/�l?#)>I�p���w�@)i#E�c}s�O���[�X[� EVі���
��C�R̰���<�EԬNNj7�rݿ��$��\���o<w�6�k���z��MR�'mv̍kP�"y\�y���`������_���斗�>����`"�fƂ�ޫC�A�_��;��ﭸq�؆�Tx)tmUkA'��waU�.�+��(���j �B�)2�\TɯFz�o+���"�l_��|�(��_�\^��?�A����Y�>�N�z
�`g-�В)�i���@C��s���hMd����Ђ15��S�ݮg	��|������o*�����|S���-R��&��AD�q��ju�d�@�w�K�l�����˿=�a���C5,�Y�c��y��q���{�oW�Q�s�0�$�T�Ţ�Q������x8�ak�\���G�XXm��ϱ�֔�����;�����'l�1����B�X��0�c����]��ߴ��Oq5Nuq-�۝����-��Nٹ }t��G�Z� �5F[\wb�����l��Hf<5���n�(�
��F��*�x�����z?��,���'����%33ɥi��PȒ%���9l�=��vXa�q�W����y�}��� �]Ҥ\�z�i���;�y�@j�P��Fc:�3���7p�|G/��zJL���q��kʢJ��[P?���(�2���|��ǻ�6�\�=���f30�a�,F�o�&%x�Ǝ1d�b�ۮ�}e�S$���fȘ�B��"�3�� �@���Ev6\(�Z=w�cCű`����hv�|(U�Humv-U0;3�O�+U�&!����tW����9U9�Ȅ�Oj�q��70R�_�˯+4��>e�_��%f����SJ��iLKM�?"�H�d�,i�(��<�Xe��hk�����JLCP��,�/��/����!UL)�o�D�I�Cg���YE�O5&i:��b�?��ކ����s��.��^B�q74E�a�	v0*��<cYe�����R+.�R�rꂿ^J�(���g0w���\b˥%�eV;kp|� �Z�˛u����Fn���M��[�Z&��\�����0�
%���~Q��nYX���q���!y3Z���m�,&Ϝ�X&!���%;^ʡǜ"~���K�{!��K�W�X�i ���*�M��~$J{���Vj�U��b�	��y�o*�Ь�Z�B(����r��8y���X">ہ����n̨d�.�O��(���h�����ף�)�n��N��9B�#��X��p���_�V���[�U�6�BS�-MN��v�!x��0xݡ��`L<���_�����ʤmј�vګ��+s[���W�2Ը��#���Fv8fh�o"�<���F���}+ۀ�\�ǅ*��P�`7�?�ܙ*+���N����`iȴe(�@�?�{R;�n�L��T:�Ռ(UF&U�5)S�I�b-#sq�ΠG�_�?R��"N�ߌ���]b���w����\�4�޴uԚE�Qڱ^ � �LB�tW�Re���V�̞Ng�w�^֭��߈�2�6�5�ۏ)=-p���$��V2���80_|0\�&:f��+T�<>)5��;��魑zV��@}P��	���{(������fمYo�WM��*;��Q.�S{�X5;ۍ`?A�Yi`�d���Β��Vik�Y�.e�\�֍�9E�8$W6Qެ΁�Շ��ۓ��h5���l�l�˅�t�� ��{ C�?ߌ>�xFN�V�T�/��~�$e[�w���lN�$�c��b���T��E�U�a9��+�Ȃ��ք76��yYt�A�ܲ�@N�,[�乀' }�`U�[���])�`|Fn���gbv��D1�6Qg�[Ly�=��G[]���m���B�ܔh��,Fw::�|3���������+��8w1Lަq#����t��ѐ8�b[	��P>�N��R�����~�����]�����b����c|kr���=EC�b�G��f��g[�V�#�z�Gȅ� '�h_�=�gSj�+��7�µ�1�B��z�9���N;G�8��|2X>\�0���c�崽�b�t�LG�]�Ac=�8����0W�D.��o��i�u�PE���^��DR.I�n`Be�S���CwrE�`�l�6�L���^�O��獃�JK��X�=HTh�e���ߊ��K����gA,$��Y�GP��{��|��,���"����p��\��9�맛�N+��Ne�Z��a�]oX��|�2�^~�W��e�I��оp�[F��&xnr�o_*ضz#�M��!��,�U�Mz��F/j�)��,�HK{�6���������;�c�4�����|N1uIL��ȡ(r >���3�;��Yg���_a�o	|R�"�I�g���U��]O660��C�VJ�1������@� �1��S?����������,Vށe
�H͂�?��YZ!�r���)�?��B���_�}��*��y�u�7n�Lu�>�� �{��8jJ�ߌ�_ka��י��|�}�>x�8�O惟�Њ�qf��`L���]&<CY�kv�Բ`��iE�os���6�Vo3��p��WJv���+�W���%ǂ�,�]�����us�ҟ�e�p��T3&��)(�4Bkhdp~�-����q *Ĝ���Vlr�@��[��9x�U�U1��o||�z�̳	�������$b|�eH��%� ?D��x/�e��g]K
���A�YbÝMsI�����?���`(��=������l��&D*a�Sa�WC�6��F+'؎z���&| &|8��&�+M"%rE�dQM���	L�]G�u�O7�$8¿��i�Gp��=��>�ocW{2�}7�Wh���:r�����I
ɬ�2�������[&D B��;����=��@ :���Ӿ�agȨ�ӧ��e%��T�T�S�<��j���싘�_����p산����i�_5���;��O��=Z�����8%Xo���v��V�%�P��^G���_�<9��;�8V��S���n��D�@Rdp��7
�F9C�8�	�-N�C-�+�,غ����t���OsX?Bj�;CY?wr{_)���R]�3aD�%�s�����	���8�=���6Dk�VZG�����K�
��(���7�Lq}�%���U�P_:PY�5~��j��<�e�z��sɌ�x:����<�ox	���'C�q𐿟�7�:4�p��[��'Ca~�K������7{=�h:��z���Ρr�C���Bp{:��sl���&)���n��I;���#}��;�Pf��3� ��s̸��^���??�߸w�����NF�ȵ���K�@J��,<��)���L�t��Se�u�ߘ5H�������?��L��b�4�����`Y��l L��f����`���N<�W��x��/�3X�	�u��8�L)���;�FSF ~q;5�8JT���{�9d�^��q�	�`䒇���dwnM=���@Y�n�?�C,HDس�e�:wx��.��@DA�������$����Y����hb��$=�$�LW�y���ީ��@��b��aY����e�[�2̠��`ZmOn� ?hl��4#@x�Q]�u�L&A�F��GQלE�/~ߡ��L��P��>u\*��hL�\��E_�����.��(Tu u����+ܵs��	��2Pf�W���~��;�_��˺Z����о��oõ��������4�Z��w)]����/�gH�T��O��]�Q�Q�9>�*�]�z�����P܉�8���>x(��Z����7��#����=p���ߝP��k�^{;���&q���e?����5��j^�� �ήn�گ�H�\R�]��?=y �#�<�Y��K�v�s=rԼ�{��x鳫��գ"��������San�J��h����U�>�g��J��j��3���������~�NJK���h,�M@W�^g�ʿ�ЂkڏSi�� ����+u�3ԁ�2>������oN#5 �,KC��LL�,�.x��*�Ǆ���j7�H3��{U��������7���u-(�V�2������8�AȇK�c�Hj6�oL�Xp���rx��~4Hi|7G�,�͜v!���?���#���Z���\̎�oz�>ѭuwf5P��0^�/�_ g"����F��c�f�~����oԸ��K�f.W�ާ���0�
�D<f��0o��Z��u�yf�
k�&?[9+.�n[��HY�
9�����#XݤW�Z���ڴDk�#�Q�B]�!��1|�Z�Zӄ�m��f��>	m�wÁ}"�e����#�6��o�Ĕ�:��B]��z� ��&�3��/>� &]BI�/��e�QDA�2���̻�q�j��f�dw��b���B�^�P��j;�Lƻ���B	>MՖ��%0x���������26��:�9-��Ш�?a0��tRlVS��DVZ
�r}�(��bs7����E癀]ąC� <���g��U��F-�k�C�?j�@�`�녨����*a�H�%B��͊g��l�^w\=z�9��.�g��pPo)ϝ�ƘFc2���g�a�~��l+��fAP���$Μ����o�_C�mһ�»�;���n��l'��z���,gO�Q��5Z���a�l$]~1&y�g�B��J���tIa��#��[���F{���9V4�.�+�	j8�����R�{�����O�&\���C=M=�d
�>��!SP=��!�I����c�yqY)>���G��v|/�2��z����biV>�
�jU_#X���V�1�ի�t�ws��sĶ��w���T(䰝�7�p��{L}�ꫥf��]����C�4쌤�]u,�Q��W%1���!n����xkRY�v)�9��ks�Ő��ߙ��e�]r��_��6�Z����%��f�8��d�|�h�ڹ��z���V�NqHǛ�F*��e@fr:��{esj~K��*��'�Z!�C,�i���T*��+(2��al���V����;�X?�>��{��)�,�~*���ڼ��#�4�7p�42�x��2a�?h&�}��!?�>g�	���n��O��'�S�s�-���ڙ=��w���nɂ�*��4�ޣ�`� zt��c�.�}莃���\A'(�`s���V��Jn������aȯf9�
�~����%6[E,=~�p�S�Dp�1�N�C,҉L�������]T+�/"}�kp���]�������R�a�S��;Pb�Y�e���U����qUg|����1}?�?m?�hng�}(y;뫺�i;�Hr|l�7���~�r:]+�0�- ؑ[��hk+b���%�+�Ʋ�Y��0�ڠ\Ս��PX��6XY�2�5��Tpb�6|��s���ľ�=�J�Bf���9���Ly�0P����+�F�q
�����Gy�Z����2p� ��T�9 ��/��:�p�(H��x��鬘rb�(o��)�|3�b'�}���}�@뤋]�J��aū3xD��񁿠�ţ�����������X�>�!/��1��7�B1�-��x7g�U>3�E:0sI��h�uJ,2���o4�� �i��X�P��sw�Nׅ���~�0�����44~ˋi�9pI�(j�O�Տ��+��?1X�Z���Lʖs��?��D����甯�9�/���ngc2����/�Q�;���
슿K��0��xA�y�@�,�?;�'El�
:m�����jU^�¢�[o�����0�}�x�[����0�tjaL��`�Ӧ��-ĳ�
���b+���Ǵ�S@�8�mF�?���6���g�zd:��O<C��]�r;q�9�X�b��5�!j<�Rlv��0�?Bh|�oY�F[i��->�Ak6wc�T�Q�萖܉�-�E��C�s�R{��Q_c� ͧQ�����\��^&����s��X/f��D��ka�5�J���[Ft�I������W&�c�I�vM������f�P"�}g�tX2=a-��'�'��������e�����e�Y�(}~7<o��9�e��l�5��)G,�e���l1T��Z2n��:�u�v�C�K΂^R^�����ڝ�Ar�Al/v�>� 
�k*��,G)j%V�/g`U��� >���kh�V�<��ߨ���j�i�I��D�v�� �J�M��C%-m3�i�= ��P�_3��T���<QZS�o�7Ө@��@��K�s���e���:wS��o���Q?xF�������J%�(��E9��@��3�E�t�t��Q��0ѯ�a��ƙiE9| 3*������H�o�.��K�[3��K�@�o)�3�:~��aT%+�����1us���<���]��ķ6u7�=��&��Y�3;� � ��ގ�hv���'ضI���oF�H툒VGj��+���2��'���n;ys������YZǿ�q�Rؗ��0&0�F�FHb�L�/G�D�{ϱ���R5��ڑ9U�u[�a�(�^s% Έ�sڌ�s����)Շ��3��!I��ߤQ�܀�F������_Q���<J��|��{.�#���-x�ʂ_xx�C��t!A<�`>�m�̀��*L��tJA�[:�J�_ p^��2\(��r��
�R�1�S��1rEn!��Y�䰠�%EҊܢ2����� �~���A���g��
����z�Qj�qA:�ܸe�Lyc�PCD�7��1蠚��P�'�0��.
�L+�t�[*���q�CvMq��n�ϛ��J�4��1S�@��(e5HvQ�L�����"�9;�9���Y��a�E����|4,�P��-#r���g���Cn-'��p�n�!��8-����Co�[��H�.�^����}i�7T!+�^#e� ���>}��C:A�;��(�Y��cv��9CC�iΖn�<�N��0;c�t2�-�Y �Cz��ˤ�2�+��Z����Ɛ�2�Pܥ"~#����i7�Ӳz���l��J��V防�(�e(u���xo2%F}
}M�c�+����r�^�%^˵��{���<� [���J�q��F�� ��Y�~m��<��
�ڏV�Ԭ��γ��=q��Le�8<�Q�9�iEm8���
�^�9����4=����SC�3 
<��E����P�=��S�7�����R��6��Y���V�yf��bP`�{O *�5��w|	��%�*��4'`t���2a �Zr��z/��������"�@��J�[%�o��{1q�U���j?�4���~|�=�;����hѸ�|�Wp	�%24�t��- �Ϡ�������?G�I�M/1-�Dc�g�x����z@z��}�Qzb<����{l΢���J������������3Շk�$�i���Q�q?F?@����i���>L~���'�c�&>���r��Y��@�U��ׁ��*Ί\��C��OGMW ��6�U����ͺx/��R1�@c�����7���*>ԁ� �s��4h��DOhޖa�-�B�*om���è�V�|��Ip�I��IAj�2����`�FSr9sZ�*�;D��v
<���T���z��%\X�N�5�f}s>�˚��_5�G�F�k}N���F+�I�GE޿(>�h)��o_*�DaK�PVG���6���7�O�ŉ���VBj��D>�'�0�mHD7���%�v�G.���a���N��t)f'rz
0�C�a0���
b�Uz��ެ�m�s������{������NG�[)s�T�iC.2`Rz;1�d���B2��u����а�W��[ٍ٫Yc���p��&E��
`�=lF��O��{H0�.-JM�6d����%y��و'�����<�� ���M���Q�dt[�\�1�Z�L��)q�Igτ��$I�}�����/Fo�(�ʂa��Y줈�N�<���K�$��_}�}��
{�����ʞf �0�Wc�=�� 0��D2��GQ����8T���*��R_�_e���9��63���=t��{e���w"���j����ﱐ���������썜�T�HW����ļ�ZNL>�w�t�8�%�R�zI�*�8la~��(u%��o�8�rD�ۤ��ל?V-	ւ�h� �](Xt��XH�[uݗFf���5f]\�9D�#�)`D�7����9r�ɿ�,���M�=-F��#�L����2\-�m��qd%�Հ��ە�`�n����@a������?@��u �}�������N$]�N�s��`��@���gn�	��^ L�j������aD�n�(����F���l5��=���A��u�B���n`&[�mrm���{��ds��H��@��\l���2�V�]��e���4y%��XS�~��A��cu��Ҽ�O�O�6���O���&��=����Y��+����rE�&��g(^��ʅxx�	7�f��Oa}��g�U�����`cxҠ%І������Z-��ϥ��oW��R�gR�iμZ\m�,l�H��ߒ^6�tR��<�>D� &��7ض���:G��8��m�$��p��	z�#�5h���.$�i�u�����%;�~��U��&D΃��H܈̄�>]�ct���*�%��.��_����F�]��5b�0 �~e�t9���6������8(��p&��`'Lԩ(	�����}��h��1\�������l;�����D��#���K[��J�ʭM�ɞ�T|E5L�+��Sb}����@ň��Ȼ���J���������m2����Ѥ����G��E枒T�(��/�N&|fS�r���$q)�%y��0̥ �J`)�çݛ�SnV���h_e���I����ǣ����e��	���3���Bb}0O�*�Cja�ʧ��LMA��:������A�b�(����	�(�ޥ�j��`�ż�#y��v}�Pq���NRDi���dh�M2eF��;<_m-��c:�GC�w�<ޭ9��鞟��0x��i���?%�-M?2��*y�=~SɤjL�2E��'�-�U',�e����G��R�v��Uѿ5g��׾���&���~��,�~:�L$���.�q}�:*~������\_Q���1��"}X&��a	��1�y��.��,#n{�a�0����B�#v=���H�#��ޏA�C�1��Q,_-͜��J��`����b��"'�F�1���l�z��[g�L�G{_C�ʻ�^���~S�qf?3ҫ�f�2ޭ�<�K�U|� � #*�,�����D����g�Y9J�Z�Ҫ��&AyIq��˚`�~O�!B"�M��`����r��S������3�P	����ԧh��[�����C�b
W�Ae]�^������~�۳��A$ܟ疯�x� ��+����C`=�� (�͵�&�iLApf�ltc��%h�,\����:v��^N�����E�q�������"�zY �T.�mNz�CNw���vQ�7���Q��H{B�p��rf�|[m��R �G����g�(O�OJM��0��\l�ܓƘ���h��k\	0&U@����E>�vH��&'�'��3o��'[�N����B��[]�>&�&���7�J�t�-�@G�uб`�Uk�+Pв���c�_'hxd�OOr�-�9���*]l���:w�t�l#-�H%�2�����.l�|7C��A��&��acd+�I;������)�Ό��h���0�",/��u���4h ���9ņ�>RZ��ߩ]�T��~v�$�B�q"��i[����p"��sH��y C��G����V*β��Et	�?N)�(ϥ�i �z�&#���+��U9taj>�Z�5GƠr���%/��)6�w��۶��4��e�M��lt��'��zO9��x��Ô��]j']9�E`�֖�������,���A���#��C��.�S�6ڂiz�v++����cp_������1��8Z-�aSq��h��8za"R�Ct(0M��r�i���7�4'��ډ���hS�eƉQl;��Y��Kv��ڜ�
���[�`F��кr� Gt�k��)%QA���^���\�߰�H����Ҡ-k�����|b@Pt����y��3�x���A�kP~�RWL�gdvO�Ƨ0I�lk�7:RVP�$H��@>Ѕz{1Pq$�oǶ�kQ1�*����
��?�%LӍ5�1*`��fO䪥�I�Q�1���+��Gr|c��[����C�Oե<W����>�>��ב�j5|��=n�����1��#:SL>G���n|�1o� ?�J|�V�%^�F�Ѭ=�������L>���{��H�)S^��d�3uB�!]x�o�x]��W7>�{+0��/�+�>EmC~�e�=��:�xP��0�閾%.�7�:��W�\s�0������9� D����7
��?�y�!;*2YZ�>�Fo���|-6��@�^��|� ��N�W�!�yX״5����ֵ�4�8��:}j�<fE
��@���3p��B��h��U�b�En�$��� $�B>���l������n�\&}[&}Je$��ơ��}�Y�B8$��$�TiuK�6�8<��a����<[&}�����A��/MW=>}o,Gi��}�v��B������� ��O���՞�; �e����PH��Ah�5��F�\O{���E�\|�W�wi�$�k��m>H��f5<�^��+����6i�a_7�Wa[��˙x.x�;¿&�X{<t]j�j�S�'B�|&������Sc�p���A|��=��p��OԎ�0Jm`�W9�� ��"2kF}j�h�o�O!H�6��{��~.nH���wK���fȷ��"�h�"����<��'���Ə��9,ʋ�5�,@5�c����O8rW���*o�GVR��r'�A��m�r��oMgb`9FDcf��8�)5�_�S՘��W�:A��Ԡ:Y���:��!ٝ[��i�Ԉ`@�9� ��4�9�
����!��뢴Mx��ˤ�)&>�mO!`��Z�*�����L�ܻ�!/��/�׃���ེZ��U|r
2(PCA?.���L�ַ�������)������ÆD��vI��l-�{��̞�:,2tw!o��$�4igȗ�����~>�a2��r�f�?vШ�����*5>�����=|`'�t�Fm����~e��������i��E�R��t�K~�L���n�2��1����v�ub��h��U{���E�}|�+��e����cݽ��>vȷO���#�	��g�d"J��J��$q"u�Б�ItO'FCcN}�86r�`9��71ϔ�0�����-?`�>��B����S(Nb5�����"+M��#՚Q��yx�@]���$Xd�b ��٬�
Qv���N�#xz�S	�x�:Zĳ�Ja�!1RVR��$�e�Bxw���+�����V�rN���1�r�}�����`���g��ޜAq?g3��?(�Wꃃz���b*��D�OE�E�\���|�������{q�+]m�r�Ypp�?<�+���\�~o�R<�B,�&q6�L� �~�{�3�l;G�Sv��<�E�Y�b{@�iC��2�.���a:\��хN�E���s���Ey�t�@�K����hAv��I�Z.�c��a�����-�G���s����#�w��(�w�^�&Lo���E<NQμ�z�U�5��G<�m�i�ܢ��F���n��7�S��Aa�A�n�z�,;���A��!���聹�A�Dϐ���%a+��4Ux��j����ل-����haX��O�d��ѧ*��eq���,���K�|p�9�������j�8m���V����[1��gb@G�1�)���(X�y8+��`f���̳�4�f�;�B�̴��s��}Ja7�(2sW<������j�����cӞBG�5CPq�������5/��=mV��&��W�w���hD#sO�/�6Rd�5{բ�|�E:����{��v:��)aǴ
�;N=Azh�J�m���d{�[�ۭ�������84Y�3�:/&ua���v��˔����A��f��|����Q'j�$�{�M���2�&�̞`P�$���3�����]̟
��w�=��+@dT�*�#/�6��8��(�)�:�;ԅ�x�k/ za�oa������o1fs$5���}"9�B{�ϓ�*��HZ*`V��$��`gMzU�����PJ����,zʼӨ �:�I����D�]ZAtI
z�^�db�!8e���;�@�_zO��^������/��x5����|j�O��:tS���J��}I=������w��.]#d��U@�`}����4���y&Qz�-_���oL��4I�ME�=��Ţ��eѭ|��̪n�؝ ��#^�|5�t�R.��U�����F�a�7��������*ߛ����V�W,|�d����v��h�vo����٦�H�-�6��I�}���8���X,�A��b��W���&�hA7p�u˂��>�T�Ř�U��5�9Q.ϓ�bu[�w�9�(ͷK%ST��bE��mH��|0J�pw���xLN�kʔܞR��otΩ����"�[cF�w�T��"�r�)��0�Z�cN 	.�C�?�K?.$�=ϴ�b������ˬ�K���]�𧴡�,">��Dk�O+T�����חq�끩䶗j}�|��z��� ����XL0��F>�f�Y7��dh�����;[��~F�	�����@f��v��Wc#J�@ե�����Q�X�s��a$�[L��NC�*w�ط�<�Zr�r�-}Mj.y�9��`'k�����C��cH֒d�0nB��P��܀���i�7-4�wi�2��F���?���pԛ4�9-�,t�N_�-\�|O�∦y����o��������ß�Ĕ\r���x���Z���	�2�Z�uQ��/&-�T+��bXBx3J2X����vmG�ű7Ԝ�!I����B�t
��wc*kjKT۸@�H j#������Z�n����k�yu�F�m�޻0��o���o��Z���?�Y�VB�)�СU�\#J-����{n�:��J[o����������m��;㩪��;��N�|Q�OM�}���?��y��=u����wJ8��!�̂����L���h�������5B^��8��#�Gt�ڍ��1��/�.�<e�\2�<���Dl�����bR�	�I����,\�&�a'��OP������P�ឤ|0���p�w �޿�����N@	�R����s/y ���>�"������&�?M�B2TǸq�֍����ȣ��w�`�Mr����҅�f��T4�,�.���7�wQ����7���MNy�����ZfB���`v��Q�*sA�;�u�T��ŌV��Ctã��e9�W!`zW����$�_�~+�9�UJ��Q�P���(��;N�¥�S�<�}���.��=�+Q�z^ә�{�H�+��<>Pj��K:gYD���q�q����/�h7XH�������}L1.ă��`��b��c�[��*��s�[��)P���u��U�VQA�iO�	�P�b��j���$���$ҳc�m8wqw�������
s��^(EdS@�"�E˵���>�I���ϤI�{���>�s{��Y8*����!+��Q,f�8���S�C`[5�e�fw��8`hS���R���-H�A���Ք���B_0�%G�����μIK�&^��5֟���*�m�"b���	��~��@0dƂ"�e�}�կ_W:���� 5�P�Y�-x2?�q�L���m!�*ϼhS����E�z��I�׽z��wT��;6cN^S�U��h=�h��@��|-�Zc�?F��9�f�tB཰�F^RX��!{Sis���-�Mȉ��:� ��R�8��%�Nd�GpӬ�bf 6�g�M��S�����$�1r ��w%Q8v?4��T�i{��Grl�!VSbe~5A1�؉^15�r�t��ByG�,)�~��y��. ?I�EL��y�w踱�3�k�_�w/k�"�:�qҳ�h0x�Ý,�+�<,T�����V���	\�;�$3����o##���E����G֝U��&��ƘS��5� �Kz�"�64�{�H92z���&��w�=��[�4�.�����w���lva��O\�-|�C]y����Œ��.|�'�{�;<�L�x�Z���%������T|�X3���HX�T7��rha�� +�ƿ4���%f1L��&Q�襛\I���o5NZ�/5*3{6�=�B|9�`�& ܞ>X��z�fH�����$�Q~�������D:���Io����Y���Z5�i�D��,�fYO|X���8�~����?I�{��/��\�/Z(�!O�K��5[�%H"�N��8�D���f$S�}����AB$L/FI�|o�|؂��1"A�yyJvz3:<�*"@ᶗD؊��Ud�$�$-2��tv׌H�[ ��u_vuI+qi��=��un%��G��r�9+7p�~�8`�-�q+�-G��S4��Jp1������7O����=W�����b���H�^���l�ao���8�gr��lX�W'Ց�� 7����*To�Y�B��c���ņ�����]O�����J�0���pR���R�[�N����0sôA��Nr��L�dzT=C0ϸ����Bӧ;����^�^��	�}.k@��=l���'�ڐ_�\�t���:���rqo��8�*���)'��{	(;� �4��f��;#��R������Ъ��*�B�&��*2��.})|h��(G���mȿ�ɨ-�1T��)U��V������/I���:�.�W�_�/�:�3�|�U#��W�Ɩ��窂P��M���+�zqCh��7���n�}���R��T9/k�N��𷖏$ o-��KH�<+�Ϫ�KD1I��� !� v�����Zω��I����X=-�ЁK;h��{%��~�֊��b~d�����Y��r���]�Փ�l�Y�����D��b>����k*���X�6*�բ��W�%�4��"�� �#�f�B�k~���x�V#���_Y,���?�,*]�@�jZU�`���ƈ��8�'W1xs�6)/p�Dx����$�'j
����'s���`6��8�ú����w�n]�R��<�K�����b+4I'��E�����_�4Z��+��g�Epi42i�ec!��%G��|�E�9G߆���\�wu��K7h�qM?L"�<nnx��-t"��X�<lo��pd#�:hs���}�,�:3E�`ԁtq�ůs�
.J��SJ�7����q�,��9c�Q�#A�{��J��Kܡ9���O�-_�<�J��ro�љ��'<�)$�ߊ��w{#�����㴖q[��x��;d��ܢ��-�S�G�|�Ҹ�=����?Pv|�S�,�zO�8�o=�CSJ�7O0��l�����	���b���O�aQS�Ũ�h�	�d$�/��]��rs%�s_+���I'��E���� t��ӫ��W6�&�ԟ~Â�,"LC̺b��\lKV��$�gȫp1��E����A�c])m�g�$�f�]��)�]\�9���k��{�+*��g�y��.��8_������6W��H�P�MTzaB��o꾾�j��� R}'�`�M���֫��Gר��z1�!��y���T������$j'	���X�����X<}�� ��E��J�'��� �	'|�N���?���H�q�g����~��|W8l�.��
L���C�(4�Xח 9�݃��fl[_Jx��m�7��oPOpQ�)��"�1M���@:W�t/_��R�2.�ӗ����^���3}�@��)�Q�3>���O��5�_z�E��M��ŀ���m^=Zm�j|+���l�爮���G=����n��rd���K�O��T�HS���&�[o��j���'$��ڂ�CEQ���f?I�����r*N5��'Z�k8����>��)#ؗ㯕�3���Cr�l�DUa���k,��D����G�I=���bR��ve�&(���1�2]�z��7]��7�����K��
Dɹ�ϧ�|a�!�����Em��2/�$B ��&j��.�1~�[�(��-p=�{'p��B�G<bA�ÿ+�%��R�/�2�!�:�1�UI ��J�i��_���JlDw%�C8P+2�0��G	�P�O⨡lD��A�������$1���eF7����x�{��;�8��{����_��Wx����b�/֌�-����t��Lt����A�����\������.��y��"�j�~;�c�d֊b94���r��:�����v�V����VmEn��Cr�A�q�6�G�6�*�;i8icvkw��q�<QKL�УwxE8�f������^�dͿ3��	S2%��A��GV�̪�e��k\�������#~�Y�-���j��p�c��9�/ɱk�������I���j��(�Lg��%8Hlp��d|�Ңb��B�:c�e2223*����吟y�&�v��>�'2���Z;W�S������Us�{3&��0�����t��EB�(iE ���Uw1��6IA�/㾧�b2��'p�b9�:H��!: w�ȴ�������IҐ�䔴x��G��>����D��ډv���?�N�6\����K�����.��];�$]���D-iRsU��_�}7�#�E��.��U��ҧҪp����ש�ޑ*9�}�qU��CH^����ne^Xɨ�m�I3]�@
���F��s�������o\N�s	�l�"^���Zb��қ���*�]�`�� vIb�� ���L�����yp3��D/N�g��h�_X:�/��q�ɉX,�b����0��?HU�Y�p	�b�'F����r�-��ˉYﮂ1���Z�{�e�G_\�帯����	%���d ^I���]|=p����6&p �_��/Y����aջ͟ѯ�_%���I������ɵ�)����v<��O�h����9��`䗪��@A҉��U��Ɗ�j<���H7�ʛRÇHxպ7�#�z����n=J��	F̊��V"�dRK�P��T���.����r�Zt�S�Oq�!s�u[�"\�T,D���B��y�u.��g:6���\��1�R`�C����	�ќa"r�ư9�� 6�T�H�`���0t���/Isĳ��̩�9�k�|����.D�WK2?���2������/Wn�J�^�XJ%�vwT:�$�C���Zf�h9}� P)���I�b�<�'w���)�n�u�7RA،MH�Oϋ׸�k�  ��6�B�h�q�{��{(p� ���
:�����������i�����V����Hƛ(,����>?O�HX�&Y�Hw:6!.q�X�eϓJ�C|�9i�3Z}'P�b�ڌ<��7f��� 휛"7GI�y�Na	�h	�{9�ŧL��c��>͑��x���+���_�e�?�ߪ�c�Ҡ9���q�"' zB���/cw+5+hn`�8�-�!�������O۲oм'Ӽ;W��(��;V�*��\� C����ؓ�X��6�囄a2)_�l��/©��4���Y9Ǔ���M)Q�1Ȯ"�d��1;+6�ѹ�=F	ؔ�k��Sm��6��b�Ԋ}6����ҭo&i�X��J�����':a1b�1#�@�_`��3��6[��^�q/~���Il�mf������ޑ�L��(�P���j�����+r���sl�}H+}����&�NAx�(�*\j7�A=���N��VsΏ��҉Zgg(y���q�{њ��U,@�1j&��'�`������ݓ
�'�XV(������N#_�CZa����0��|�:�>L��5�I�'���+�&.�o�G���>����_�u�&��^؉hP�
�''x����B�6���إ����V���:u��#��]�ꟿT��Է�r�U�KKfD��t9����A�T��yR2KDG/��o��?D����J����e{]/�i�\�����K�&�E��Y6E�Z�
�,M!�t>}����N��D[��G{�Ct���S��E�fi��V�F��%�[J_B�!��>��6ޜ5�asP>�LO�:M��6%xG�!�����y_�)N��bφ�l�$q[:	���Y��%���f�r�ZD���p�:�_/ؙG><�C�9��Õ�G�{�9�-�2��#�|H�m善���K�
"}P�צ�U��>��}W���n��ў.�O{#��P���9�[��-�.�+m��9���53i���I>��>1=}~\�����Q�~�����3���<D�#"@�N �I7E�:c�pB��IA�ǋ�c��Xh�J�����T�x݉/�mf�$���g���;��S�R��\޴�Z�D�U{��~�ǙH�{K�'�RY�>Y�6�E�v��`-Ó�%U?��o����~��~p|�q;IDo��Ձ[:W�	>6���}����ڊ�?��m���a��r�g]P�~.)+$.A2�/����m8��$�,&�}�����������2������b\x��#�Z���D���vK�T��GG�-��nO$�yc���`L���Q�2L�k����[D(��M?Is<��j^j��w&����L��ʢ�і�+~ ˢ������6L'.���̸;�;��2ۿ�`K��K�a�G ! R��*�N�t�����$�Z��\�5�=�ĕ��I��-����=�ۡ�dP75F���;yg���`R#���<�'0,�r����4rV��oƂ�rE��`�������8���4Q��F�=���	�߁y��$Nl�Բ�ތ�D���m��'�����'3H�nR�N�d�a1��jRr������7�A3�K�=p����}��n�P2�L�������YC���7Wnv]֤8ʢ��u��$j�~6I�I룎��$�u/�e�H*���c�d���'���U�P��6��ی/���ǐ���l��io(�;=S/�$@|s�9�F׽$�r7]���T'0��P'� Le��U��c��V�ѤNȢO�'�����Ԏ<�W�3�w�����ˎJ��ԃ��E��Nn��Ѥcj���r$�s���x�P���.:�SQ���kG���y�oiO=)�78�t���|�_�'mpJ`�k20n�� �^!7�gx�vt��� m�h�U��E�Q��Nd˜����ӟx�U�rsU��ܥI�"�px������������B���p-�?�a�ܬfd��"���*x���f㧫��
|��_3[�:�!Q�K9�� Z5���]qv�+�`�1�A0vG�Eg�"Kݶ��y$nu����l�L(���1��8j���ܜy��\{�D�i�[N�΄����h��Y0̾lr|��7Z�F*�]��I�=7�}k�]��}�4s�v;'�?Ĉ��9��Ĝ��ԩ8�>ٲ��ݰ7ޕ�q
�T��&KJp'S�BΨ?"�����Ͱ+�Dޠ/ތ� ��D�����9L
̎�h����.d�eG��Z�(���z�=���-[Ti�O��ύ��P9Hײ��:��7r�fŹmٟ�^J+�M"�[�u��Z~�<��k��}L����#|�3�m�]y�{��^�VG�GI�k,��/�`9AZv
�^�k�G����-v[�w�H���,ص�xJ8W69�$�O�C��!!u��%\MO�96Z֭j�{��?D��mM�oC�����!���zQ2E��Ik��;�Kc���u� "��4��<N��(��}������<Ԟ�����lQ��IB�8��
"���_g�M�$������3��n�g2R/nq��u������6��qc�<q�|���r�AMߦ�t�ܑ��=��3Uc�D9|�Ds6Q��`�$�lC>��a�P��t�N�,˾�]n���茈wT���T�p&!!�06߬��#<�8cr�O2����è�_�AGS�0��I����.|W��6���-�l���w��K�p^7�m<5k��f��������쐟��8��6ؖ�ܺt�Z׮��c|4�|	O� <�\���^ �����JZ*lu�h:<���8w.����[:,Ci�O�=햎�#�f��/����Kp�,u�q{�v�R��L�,�Col���J�����V�4��1db������LI~
�hܑ R]b.�c�J�ͺi����޵!���N��w���^c��4k��>�j�I�_��w(z+�εM����Cb��w�T��:������&�0qݤ��fU4��4eC&)V��c3�km%H�R�k����}�=���mkg��C�t�.+���|���֟'���k|�աߨַE&_��'����UG�㳪#�����_HX-��i��A�7;��@3*��H�}�6q�k�)��8
}�$����	���ߜe���ʑ`��(��������f��S%G�(�e?ͦ�+G)M�xXAG�C�/X�g����?�o��T9�֦t��q�RI�"���(Mn�]n��M_}%]�)��iGH,�����w�}��5�4��
1RI��p�R��3��D�'F��W��Te(�貊���3#��gF���H$�|-��9��J����J�JX7T����S�N<����k�#�>s�$�>�
�'�+��.�xFF��-��u�/�[	�e,�X]�,:=R�����K^�d�V��S��kT�5�B��sz�1���tme$�T��W��h�07���8������y�R����LSr�����fx�\��t����Dr]�w������zI�@2W0�2���P%`jģ?!п�N���B9����g�-	��E1�ڥ����{���Hff��K}\���r��V���A=�j2�f�i�?ζiԽ&�ZR\����	v��T:����?�Y�A����0ˏ^}�'R{��g�Dm�>'Y�)9㼓�?�#%�9ŉ��g�����;�T��$�qM�➨F��<.�����LT��č����R儯#��ގ�ƥi9���C�H�RJ:5i��Q[TZ]�i�h���-g�E�ǔ�s|��"f��q"�:r�Sk�����I�9��V���P%���N�F��c�G�Z=m;1�ݬ�y((ޒ���/X��f�E����ފo&�9p��s��|���)�S�w"(�rw�޼j�M�@B�$���M�t��bnJ�����"ެl����r��ÎI ��(A��V������4�5���n�Y���%j�y��e"������e�=F��ڤڢ�Eh΃�Z�A�K���i���Z�I�_S���Z�)G�pF?�m�yb�Kk���F���UF��^O�!BlO�a�:�rm�-�:��ӕ��h��h;�]eT�::�hCGg�-��TF��,J�r�)i�闛�~�Cd����;! �]�G���ߐ5�ld�ќ�������a�����Ff���UJ%j���B�=�βO�\#b�*�}j4�}HA3��ۧ4/I��+b��9ވ��b��w�g���}H�L�n���a���0ao��&��GM�w���4]Z����w��/_D3��9-���n^c�ĩ��*�X.Gp�	�t�%���E��ui5}�m"o��i�S:�x�G�|������qGY�yWM�8'�/"�Į��`ۧ��g����b�����H�^�c[�e���/�%�G�}�j.jvP_�M/W�(^�!��9�5���d���A)p(6~���kh����&G��C ̉�R۹'Dih\�������8O>Tg���Hx��F]�q�Tb��?�f��r���/���y?�ק<W�2ݣǈ�w�\:�u|���UR.��M�M{c�8v��z�N��E�Z�J&�?7�}r���8M��h_bt��l�dR^�YQ�4���I��y]1�I<��z����&��?�D���>����<\{�����x5�����)2���;T�&�h��N��*�[Mg��Cr�ۖgU�	�>�Z#�-R%݄��+/e��n ����z7���B4���J�D�o�ڢ?ʹ��ݙL'T��g�D�B�����|���%�����upʞ�C��ZN/x�($��Rc�'��}9b`p��ԓ���XJ���f��=�)�
�����T�W	f�
WI��"������Y}�ث?A�����a��I��an��7�k_LH�2e�(d8��~��o�yɲ9��a�6T�0��o�����.���`js$8Jv>h�(��s� �e��Č -�&A�rd�*�D*Jp���T��{�I�b���?�l�X�{�;r�C��l>��;����XM�� ��W����ϲ�$m�̘�kl1/<�+NN�ur���b����IDI&�6"�ݠ���\?}�ѫ~�:zV����H�c�1�D���v�a캂#��ϵ����x����OM�~u�ѯ�ԯ.E��ͳ�td�����7�L��o!�^��J㚢A/�������Y���dҨ�6����-�̷���]��/��.���[ow#�ߙƈ�ݕ-<5_�ߒ�i���ǧ~��584}~{H�:�f���A6�N�R�p��u�J.�<u:�0�pc��Ϡe�ە����d��iz,�����ÿ.��/u��?�ڄ�:�{N[�ܽH�w�M\��'�KU�;gsW�onS���3�;�D6\�����)��}���l������������f�f�l��Ad�*��S��KWkƏ�����ґgӜ�oQqS�� ������E�i�^r?:����9'r9����x$��jqD���vb��z�$���W0y�]on�I/W(�c�U�h�_	3�&q�aVL�|��_L��ִ9���r1m#ڤ$ދw�~���h�I�`ۥ�c-ɱ��<���F�Bv���z`XB zm�
��#}J��p^������g���=wX��	�ؘ%Y����/+OX�0�F�`|)�6�KJ��
���;���KP�)��c�qS������(�~���L��S�S�ї�xg�ďF��ۇr֮\:��4}x����C�m�y�酦��=i�����M�����6`=�-��Q��[ʶ��|��έ?��$ʗm��tX���>y�6rk~�|WTX�[�B�yh�)���^�,�	v���_�k�+N��d��+Ng?6�J;����*�#�����\�q�|��R[PC�Z�"l���'f�:�~�aտ�F�*~���d��B�~��"�΍�������_�f��s��(տ�޿�j�cw��f�i�t*���'���z�ͣ�'as��V#z��B��>�l����ץ��)g_F-�9�������lVDGh�{4������!�d9ը:�@��`�^��"�O|��\I����S�='����tk��@H�5z�X���h�S�a�]ic\�65<O="�C��[>;�G���YIb���ٶO����ؿ�<�zWTp5��v��Ak�̎#�^�������i���J[~�8����<��p�2�����ٱlz���|SI���X���䢣��0�E�uwj�����N�#i�@%����G���i��^n��i6�'O�Gb��T�GfY��s��h�drO0BM%(�w��LB��c��[4��`q�,�	��h�4	�����=	o�z�\*
�8R���{��bR��/Ō>���2q���J��O��j���r�:�r��v)k'�)�7���V ��6`.[�QwO���l�^���m��a�ze�����yr�T�Y��K@ L���o�X�Uz��8&$V3���#Yt�W�G�-�Wn��i$gDì�M�'@$:§�Ӥ�X�����C����$�~\�*���h/I�\|3�*}�JA
�U���m�T�����W��J�t�"��)%��9-]�C�sj��rs��6�Lg��ufK���`O	M_&�l5�=+N�˽ztI1)�{��3��!N��9����=ztn��?��ӻ5�unlķ��6��/�O�<�E�����t���ɶ��T��%����ϖotj}��A��7����[ih:���Bs����mq~�F �-���k(|ڼc
�8�`ܖ�曃φ%�G��9��Ls�����N��� ��A������ۘ�(�{ΜL�jN��dMh`�Bސ[4�72ڶ
>ț�{/�ۥ�v�w_29�����Eʊ}���?�6�&6��h��,���u��/���1\yn��54U�S;"��gS{/�L��|K�������� �W��T�΃��.T�@��4��Ⱥ�D`�T��h����?���^d�J��%�U���ռ����kY���!�r�SJ*vRM*�I�C-Rm�/5��ߡ�Ԕs�w��{S"����Zn�ߡ���4��:��X��w�L���3��C�I7�"��ᢾ��yw�O��8=�%7'̵�&��\����QI������Np�q|��Ӧ�Lם6���(� �zs�5�7��Z���[���{i�Ap��g�˧+���rs�P�B�~r�y�?Th_�U&�O�"��2�8q�-r��eQ�@�fpU��=�y�'^[�uXʢ��u���?A�1.�K��/�I�u�������y��^�u�_��]:S0[��YYq��/I�B����6��W>kh�S8�X����F�������6��+C�8^��)���ȣ:m��*��3�|�%���k�d��|�e�V/^h�f��>Ƴ��}$�z�~"xq��R�i�15�R��Q	a{o�eQv{��-<���`Z��]�]�My�5���O�����6?�ґY�CR�MXiҲ�A����TcZ���f��Őɡ���1༨r�-���P�.u�fړy/��'��f�Ү�2˔�V���E�.)=m�����P�<a3���,)�җV���Ɨ��+��>��#U���~	�(����л��+�%�7b���4Z@E���%�5��x_"���)�0����"WG7������7RW�"���c�|��=��ܟɍ����Pv��i��۳
�z�Ћ=zC3�#m �wi���dF�D�mB��JD�)�G����T,vz����@�<F9GQ���/L$k��'j��>���g.�.i�l��7��O8l�Y|ud�)��H���"�o�a��K~��$��i��<�o!1@[��KB݁�����:���4�żw��cL���a.���q[�����>�{|K�;D�_�����\*buW�^	��=��H�Ӊ�Ht�g��ʉwhm�b�1��PP�=K�B>iy�����R����H	~n/�S��4���<ܽl�i���j$���4{�٢l�����<x�i�'$�߀+��s<�|7'���1���_]��cJDD�;�E����&�ѐWm���tWH���46rt��t���{�h�0��o7s��R��,�H%�W}���Dnj�pTeu/��(���S�D_"w�[�:^����wQ׵Y�b[��%��U'�Ns�f�ǂ��+�Og�+=�uc1aks�V��Z��{<^r���]O!��tɃ�n9<��u���<$&�m'ޯh����6�؊1<O�d�&���46a�x�5�)�����h�<5l��FIr�+Y�yi��ϭ���!�w�.��PBn�Ht�@�@�"1L~z�KO'u3���?�U��D2�V�G�G2p�1�H�my�����n��mn����s�3:i�N��m"���y!��a�CU?ID/�j���j͙#?{ ��3=��K���i_l�O[2� }�_��<"���QIk=�<�X�����K'�Y԰�@z+�!�?:�])4�gPyI^���$��fٸ�R��(!m�A����Ǳ;����2��!�&# �%X��!�eg��4�Ӆ1_igF\�ɕ�qiyV��{e�Ǩ���u�M�d�ıW��V�gQ�U��k�|�2p�y��ıZd��fKE������9��K���D�f�.7��j�[0��>d������r�׏��=��Kb�+Ԥͱ����^��/��E�'177R$�m��ѳ<[/�{{E�1�}�lN�Wt��i�{[��C൩d���ֽy���MtHWl3�!b�AG|��~ ����&���9�;������8�ʅ�0�C^�iZ��Bn�%�9�M�yڹae�X���H,c8�$}����S�J�0��_��'���J�.�bOo@I����������l%��耵Z���;�{����WR��7{*��}3��t��}����y��o�/��z~=�����3��w�4����$����WQ�u�ת�����	B���YG�Ȭ<���%�}��l��K��wH0��Vϖ��ՆF�bDp��Dx��,2�ÓI ��C�F.x�9�����Zڭ$��o�s����*���_���������U��X�o��zG��tyq���n	n�ʐ���-��Q�G�����6˟�P�z���8������(����Ǿ��E��=	�ɤ�Q�.+�y�Z�3��ϟ��� `��`EG��s�4}"58���>����w��^�كI��b��S=dw�i��>b��\ǹ�ܓLr]C-{��F/�E*q؄$.���/�����L,��ګ�O\�U���F��zaA���$�Z�ܞ F��s��E49<t���p�C����^b��UyF;NΝ�� �k�~�d��׌iž�c��⩊q�f,.'Ej�����IGŹݍy}	�3�5Ą��J��7sO��=��H3na�x~#s��K���`Z>���ML�'�-�`
��'���r�)<ƣ��{�ɚ*2�[�W�4�<[R��P�܋� �Ē��R%6)�o������t�CQ�=��G���R����:ĢE`�b9&P�/��ˮV'ٸ0����*/��; k�tΚ����&�����![��^�D�r�����X��E�L�������!�G��~
��cM_��[�RWB�+5�{#�]�?���_��i5r�1܎� Z��Ax�(�V��I�o�ɳ��a����7ǅ�׹?�?v5;j�.HŻ��蟦�K�l����$�Y�us��T�^��	�W�,�>ea5-||�wز9��v)0ܨ�XK+C�<,x(w{/�(Γ���\�E5�7��S�����}M������$E����`���Z�2�1���v�~v{"�TE$?~ )k�7�I���c���_p���g@?ef�r�Y__54�����)��ۼ�[
�do�Cq�O�Pi� G�մ+�i��l
�O�3Gͩ�ޤ.�T3Vq��~̣��u3��b��>�ǹF�����,��Kek8/�ɬ��w�H$�	��n��0������� $�>��q�p�27��jn����-S�yRӐ�b+ǩ�=f�R+������.J�&�FQ��J��5���~N	UL���orl��uK~����E`p�qr�MX,5�7I��/��=ʖ�<�>��(
s��g�����<�^Y[�L埇+��ޥ����?E:`���4�7�Ӧ��
�	䲃�p ����A2�(םO%��2�5X_6�����@���Mn�e�MP���r."��+*�����4�|��^�,w>��]v�`R5&�J��V~�u�cB��r:zwAE�%��YYv=qy�V�~b����H���+���[ˢJ�ԋl�����w�>���6�x�zr1dvh�yT���#Ѵ.��JI��lO=��'����y&�XY{��zt���$n�O\������CE6���D���&��*��Q�E^Ӫ�����ˍ���nZU����(e�[�ars�ȑ�L5��觱X}/S�O�0�����a���7TN���h�WО��4���������迎$�N�p��2z��rU�2�pD�E�W�+��_ABeYOx˲K�򤚂@�]������?~;�9J�`�H�'���8�A�mS#�$�P��W}\2]OEUa �q��,-�9�I�
?RN�FE�f��c���<�~t�����7$�*;�ֿ��k��S��P&�q�d������ˍ���e��2����9���`;��Iغ�n��;���%�>�o�W��Q��M�K�O�}��5Of����0BNj�B��Q-�σ8�3Ʊ��51�y���H����B|h�VH� �w�EuV}�`��"<n�sx�FsHϩ�Rm�k��[M���ZsHi"EQ��-6#���/�ņ���N2��k�bWK�P��}"�݃���l̚ϥn��EN�j(�
�9�/Hehx
=�f�2��Q
�~�n"%O�G!���8��F�x�W�B�a�pd���:&p�%�:�?Y)PYС�U:5���`4���R���V�(��ѯlϰU��(3�sYb�!�q�'�*U^k��6{����۬fX��5�
^Om�;Έ��x!��I�[�B5þ�;��}@ ���=�x<�����H�X�_g��C-�'AL���BE��Q�N�)���7��?�I�~&�Y��U=�5��du3�Bܯ�����ۂ�3O��ЫH-Ӳ��%b�FN�s�G�I��s�b��۝\�Hj��.��Q�kj���8���J�� /]�M�&�2��x�5�����p#v�I�l��=��q��9n=���26��rk��nX�}S�n<{�o�&A�6(�d0��/�mn%�j��gO&����+���]����S��LD�<.ͷ��7�OB)Ey�Z�P�^j�B��N����X�|�h����$��$�k�p��k�{�����w^(�rPy�G�k�T� ��ļ�Ĺ��5Խ�"bKU��뮶YN�`V7^I)�yȚ�f�gج��E��c��������Ѩ���G~vA"	����������~�L�꭫yS��&��A:=��ئ�� S�&Q֣~:G��爆����*�I��!xA��.GД0�Ռ8�bY,$tH��ĝ_.�'f�������5c5�;b��TtOꂞ�}��͡)�5�"EjY��T�
��'�/J��=����A ��E �O`"�cF�g�8�;αo|�8��\�1BT��R���_W�v&U�d���j�\���V�j�����n�p�.*>�Y-s�X�~Z����&��3���E���-���խxP��,�j��b�a�u�+��#
�����|��s$9|��q�����P��YWm�|�U�7�ܲdN?�A�+6ͪʑn�HY��j+b6͔b�S���Ib+���P{%�>�����x(����`�x�x1/��u�,��an϶�y��-��a�9�}3�-�/[����n����M�[��-��Q�]<psb�qZ
O!q��C'�t�?M���V��i��ٕ�6;@�S۵���_��Gȡ 7���f5<��8�(8�n%x�r���n9���n�b�e���3�ιeԸ ��9� u�lk%���!���z�r"ʿ���vY�a`�*���e]鮦�
�FM��Z]rh6ķ�w$�ER5;87�?��r�S9\��F�T��YO������B�<�2�R�0���	lc��w��ٛ`�T�c
p���9��F	�D2�l���",����9�u�w���Ep^`HAG# N�ß ��;�*-�Ch�A�?��XL�Uh����M������b��ȕc:���~��y_�iE�U��`�h"n����?��+�5��^፳�z�7啣8!�cڊ��ȴ>1'PX�~��X��H1<S$�Zis�K�5��By��h�;	�S�P�\�����N^$҂˝������Ǔ틇hƨ��L)��ĉE��x?����U���
\��.�/FJ�<R���U���V+���Z�*h,�Y`�B��Y3>0�W&!Hb�'t�Ԯ��7�1I���hF�m��t������%�i	0���������z�㨢�ї9D߲���g��<�}+za��,�C7�ˆƯ"n.�귺��g����-��A+���tz���C�!����촻uz�Dj$wA�6���"�Z�>L鶼jcj�n�0�%R���ub9el��;m�N�Ʈ��������ڢq��GG�]����y~y�=��������t���>��/��������u*�R���N�PPV�dOq�2�ޡ��V.�M����.�Է<��&��KDR�7�U�f���ܺ�hܡ8w,���	�T���@L�B�$�e�i������,�BV��%������W�`JA���D���'��B�c�=!�ZV�@uU-���_�;��[jƅw����I᯴�,�����?����(�
I5n/� 4��<�;�z�O�?����0�u�?�;+�1�����
�]L���&�L/p#@p�F��=7Sv��⨼!��;D��F���M���q��RY �̞@=���T�D�&~�Hyנc|�ӽ`�9��B����	�B��&o���
���#Y���\�EP��բZ�NVU��Ü��$�B�crK�F!q6�b� ll=cxۥ1��E-9�wdH�����S�}yr�׈�m�[j���@�i���ǳ���g�������Em���i�D=5��C��(��[9�5�Mm�59ѭ]����I�Gɡ�U�be=�%�-�H�C՟(\�����%���;��D}�N����V�p�V�&�6hq��#=�D�Ū|���Ԓ��h��[k��_IHA��a��������)�~Q���t�����u��.0<2'�6���J�|j��h>�V�U�UD2���c4��0�|:��f5*W��\ۻ�'[� p��I��]v{)s���:�sz���I���B�X8��k:	��[OMϩD*�u9�Q�D��x�OY�g#N���w�����K�T�m�Pq����u���-zJM�š�����H�nl��4�+e=>�<�	�b��[������T���l<����'�Aݬ�&�B?���t
�䖨�2����JEߊOm�Ec�F�C�}�h��Xe�7t�`�G�
�H&ic���E�E�:�x^������Y�d��>V`[6�߉h��j��&�D�8�^��������ϵ�R�*o��l��}�P �\���*�ܮ�3&�ԛ̿d'Q�CƷ���À?��nǢ़��j+23f�A�G{��{�}�ڰ'�36���^�I�	mpX�<�>�'��m�=^w�_ ��N�`,H���������@���Œ�"8ya��j�if��䤊�!4o}��;���� 
�_��@�&Hu��܊u`�A�"�+��q�3�U\��(-�WR9&�:�P����"Z��\f.�S�cO�M�g�>�6��E�i�o��1Ά���ď"b=)��������{�����e���Eo��q�?�Pp�H�9���?���R~{4�����y�{��\�s׷{���9�}x��}�.��|��Dj>�%p���%�~lz�q,��dkT?��p��T�����[�Ӭ�zfWDa б����rx/���
` Wu�pй�3T��}Qu�NnF5����N	(B�ը�/�{��9�v��$h9�	g,-�D���G*@J�`�P��w2�]��
>VHܻ��#SݡZ'kD&Q��A��~��2�����z���ۘ�W]�_E�;_j��T=��7��)׌8�����s�f��*S�O�7TMT���
����~�S�EQqI
u���)����]��f(�, �G��*�uV���Q5��uW!}��,d(��i:a��c��'���.	�U�O3�F��06��iW0=(t�,{w�H�^������@V�ZK�������1r����&HO�Ç9����=$�����et�� ���|�F�/AJʲ(��j)�ziΨ�τ vߤ|)pT�C���� Z���=jQU�:n�J�.d�/�C�1���w�_������=��{*�fƐ,Uʭ���>��zȥɅ�e~��ڗ�*�ԃ�Mr8 jǮi��ڇ{��ٵ<iޤZ�,X��F��Y�>�?2rk��]L\�~S����^,o Q��Dm_"9~Zͺ�ux�Bu|m,��*���:�"J�Qm���<��$_�w�˺��=gy#���,گ��r��-y�SS�<{ǧ�!���iG!�='��/��	���ו�}ի�c?�'��&8�F&�L��@�ʏ}S�	�j���Ա�{E�g]��±�\)=���m�����9H�=./񉅬�w��XB��$<c����ҷ���c�Ί��x����ԑ��2���q�M�OψF`ܮk.kd���3п��쩘@"��gDA�Rxr?�m���|�M=m$�t��H�5�J��+$>@��շ�Co�S�=�#��Ȃ&���]\F�S����e*�'����#鮘�i�(�)��Ū|{9ro��`\炢�%;cg��<R��"�$�M�^��=M�q\����	~G�Is�0�R��L�$&|��0j����3L�P3�h�_!�(*1ƿ�V�% QE�ԛ$T|���M�A��G����a'��Ǩ)t.�ڄ��3�t��R��[UΉ�@�$��N�O�0�b.�F�xx��:po��R�s��|���� I�9]B�d4�]l+M�6�5�B��^C�SQe�$��f��e#��J{Ί��3WQH�:�sϚ������.ӗa]nj�.�s�0a��,1<p�MEC�`�m��K��ˢ��({9�
Xc�.�-����������oc�k��+�J+��.�>cTEkT��&�`�=�@�
Ŝ�)z�#\f�5��@�'�e��9�I��`**�5�:�\|.�g�]p:Cg�pj'�_�� K8��g�)�H����x	�y��US_��t����AW�x��Z&b�2�;�v�i�`]�~�+$8����iP$���7zP�����5����6�yĵi��ӝ��]DDmn��"�B��x_1q�ae(�)��ÅU�(�yv`O��r��d�N��:gIFOjI��f�k�`�N��^����#X#[�B�r!�2��Y�����FZ�}A�*;D@����'��k�l(��]�N�! �ǿ@���7�g�BQ�k�$����!o%o���`�d�M���}���0|L3�8˳{�7z�ؐ�S6�'Ћ���<��z��*���/�3&l����궾�E�_jY���ܒ8.���ϊ�p�D}�$4 ��A!��:+��䡀q!h,4�#P��s�%=�������E^-j��[�>懧��v�9Oʫ����d{��
I��2�1���*����N��e���,=�K�ϵIr �� ?Tk����ƪ����?�&� x�����<�&�ƿ!��Qy}����8�T�ށ�����'�R���{W����eKJ$؁��1Z�g�k�"�>������[3�"�� ��$��%�v�\ϩi��l�_ ��"�����zR#�bC�z6�y �48���.;P֣lP~�sQ3���A�
p4i�����&BQ�xT��Φ�s�ǩk�'
m���rO�WK!$;;��2-����̮�M�ݭ�*9B�z�x�U��9�u�'z���f^��QY�IDW��O�Q������#R�-C_r�;����f�q}z�Pո�޳̫E�v���x]T��_��/���՜&������X�������?fֱM+]8醥�J9
r~�4�������)V5��U\?�����f%�Q�z�.���G��r1���7�k�a�E;{��U_�����F4�P���2�qM�ټOŵ��b�o:�D"br"���,[`����]\���z̋��D������L�cyQ;��/?+�{�!�I���#��?ߪ���U����d�W��y�Dу<���C���J��`�Ȥdƪ��P�M��r�R�~֛詪�����y<�R�Ie�|�eSlˉ���9��_�N�r��M��ka�'Y�[X�?��Ԙo=����ld}�j
�����-,|v�شSfF��΍�&�F�!]��Lk�Ш��C>}���ҞM��sZ��!�i3_X	�P5���["��D�4˵��W>B��Sb	W��<��xo"��v"�;G���%3����6�a��'�e�/������{j�ݟR��2���{������/@5h�C�
ch2���²�qO��8G�֏���8�(�M������ϭW�w&/�E����*W,d;����M�ۺ���׸�ɻ����a��m�ެ��DTvH�d~�տ��՝���|k�'�^H2UAS~9;:O�/�������m�������S����\��P��dܲ���2�Z��.�x�#���������,ڣx���p���>���O7�+;3�Ă�,T�w�%MEr@9tU�,nEَNQo�'�o�	a|���S�!m��M����;+�=*���~�i՟&����Gಋ�U,O�@�32B5�.J�����ǙIWC�Y,�TZ���,��Eo����V��	Ldn�S�D����x�N��'���K>��ѣq�(x�>O�'Yӌ�R��{�d�������'Ռt����L�0���|��4GH$����q/=�ϧ�,�5|#L3�9//�ppmj�Y0�PucYq�������fMSD��T'����pwA<����C6�
��2�졩�5fpI5��V�'��L.T/�R%SEW��Pn{���a�ڎ�k�8���b��.m�O���O<>��֌[�i���[Ɲh��NL�4_�(����冖�:_�ɫvY�H�x�.PI��.4��?ړVr�*����;�Y��~cӚ��eL�U o�6���Z9���qm�0�Q�QL"ݞW�|���76����!n�RO��Py�׭��Y�D}yƯy��_����X�Qs �e������{���r��!�+��f���s%8�:�a|`P�ISl��d8�0�����T��B�CiPb�mЌ��hbsrհ!ί��Z}��j|]��)� �Y���5��7֖ȡc��T�&F�zB-�x�e��3y����r8c	�0d֜/X���n=� �1��H�E�[�U��KJ��OҸK�4g�ڐ|����Z� ��]�Kwy�mre��1)��,{�mn�K�PX�����$���%�B&����h��:=��������4�ݏ:�_�\ �?�P\��` Ғ��K���6D1����ԭؤRA�Nt�i��-�?~�m�J�ǈ�����S\97����^�.��b�ߧ����V����|E�_O���9(��d��_�/2r��7A�a�� ȱONA(:j�����~�eV��H����Q���nc/�;��:����E��`�6(�j�p��	�N�ދ��f�#�%� ͂u�~rvP�_���#�C��j=�o���-�C0�W�����f�򴘗��qOI���q.b��SvE~�!z��"jc����Y0SsՖ�>���_�p�z�>#��D�j���-�za\!A"ck�-�u��?]�Vt�ө�6m�l�d~L�(�r�1\&�h��s%*]hD�4�֙!8E��J��c��SAr�<�au޺/�]����w/?l, RqH#S���Vjq>����ТK��_�<���Hhf�p� ���a�G���$u/X�'����6�<�y��5��f	Jp3% ��6k�?��FG 9��U|�"�TΎA��|:D��ڸ�����i����}ZZ�b�XbB�"�%�!�d��/rx�<���֛zR�0}�wH����2f�|����f�鶳� �h�c�:Eos�}j��1��6�M=��Ǡ��~�~�zײ��4��#���F&V��8�@��@�[i���A�uͼ��O��]��M���GA�*��6�У�"e�;
=N���r�����|e�7�I�6@a
�P�j�V[Em�@��0�T�E�����e� ��&��q������yw�uW�u+�
IK�JU.^oB���-�y�9�L�Rv�����K'3��<繝�<�|�5�#v�[���K~�&NƯ~-J�*3GUXP8Z��_��@�U6�+K�;2*y�0x�9���j��"��T��f�l��ϐG�'/6�ej���rz��z���`�ۧh�c�k�Zh�V���O�H~��ř�̹���aB��ﭧ�NViWSi��>��3+KmU{J�����D8�(�Ṩr�����9͡�m^�Udm�y؈�3��9�X��R3���{i������ÙUɬ���;�'ۊ�{ٰ�7�d34K��o�����Yc�S� R;�:L�[0�7B*s���B��p�H�X��lS�E��"�G�+;���w�ڦ���kܷ�HC�Ʀ*��0k��Dl�V�B��*���uap�"�8��{\���w���"�Mu3�w�(�}���!��u%#����c��M�D;�d<��ZL��.B�k�'.�.�}��O��pP9���kx~/�6�7�����x孁t��B�^_�����+mj�Z��J�D6���!B*su�|�4I�#v����?	�-\��D�0"�
����u%��'�rWbz�-�9.>�y��5>��4Au�K��"l�o`wXO^K)�Ri�^�J��Y�x�ZbW�*E	EN߫&j�.�4=�$��ʓ,���������^�V"�����L�����0g9��IZ�)���p�r=�T	"/тOHH�)¡.�(Q(�v��,�C��,^��e��V�d��?ՠ����r���ѰL�2ʄ��]Qv�@e����a(��4�݇^KA ى��z	!NMx6�q�kI��=��TJh����}��-�G�G����X�����%$ 8��]� S��tR�z�x����_P؏�$���,2��EFȥ��b���{E�o��8���Rt��.�(�;�ڪ�ؐ�z�f�d�P
� /�*r%�G�[����F*���s�8�;jj��2���2�%b`aX�vNO����9$�.�O/wRi(>��I�␏;Me�2*���N
[P��D N.�������g��5�t�]ןQX�p}�7}+�[�Nߦ��b?�~�yJ�!�=�cq��Dz�ꊅi�{�Z�:�H���V�<	�~���D��o����}Uz�z|?�q�ٱx���P�,C�ٿ��3�/#4�P��p��١H{_���������В��i��s�-)�4��9xAMQF
���@q7&^�ψ�zL�f�KAh�7�Q����^�њx�9�q�t
5S��8�[g,/M���0�x5�T��0��'��,�[�{J:h�i*uʽ�x�K U�<��F����(<]�F&�!��~�p�O|�۶D�?��m��a���:�%FB|�6H��3�����c?Fc ؏��0	�sS �e��G�������΋��-������W�����̞��_O�Ï�M�����ĭ���;�xw\T��\��ލ��Ee�5_�Lo���2}��z�Xbk�A�3���: 5λ���i��νQD���o��5}�����Ùo��Yf�PQn��'v�������\n�D�D��l�T�z\�[p�4�L�B��ۺ��L�IIՃw��������vsF�z*#h��y2&�%���=��_���3��y�,��9�G�r�G:���'ؠr�X����R|v.���:�"�Fum�p�jĻm%˲�t����s��Ic�m�4����\��<�	s�G�:-�h��t��DN������:ȤE]zJ��2�5�.'bZ����l�%k9�o�.2#��[�&�n%"��o�I�7.¿���% j�+A6���/�I|L��⧽� R�L}���K�'	��1s	������~��ڭ��%R���t݀H�<R&7�ɟ:��h�w�@�����Ǳ'3����*æ��/�_���ilUk6w6���~=9�J3�w2�E��y* 2'�b�:����xo�Sd�bgvԲ�Ȃ��f�8Q���` �ô26���aa)qw�.�,�T����_���߹u�i�0��}Ǳ����o��!_�~�E�>&R/z%�t��Quy�(��v{
�ѭL��͑�#E�ׯ\� 6`�B����ί����/���� M,��v�#��qi���^Ɲ�oar�	~n� �O��X�fk��2��jo�4��G�fK���\�M�`3щ��CK��O��rg�Vi�P��z9�h�Z�xF���g݀��x�|@��n4�����ƀƔ�K�My~I��S��{���sZ=�	;�1f�RD���j��E�^|���;��γ-eY����w�gQC'5�6��73��Ʋ=��TRҰ��[�>�R�d&]G�q��<ɂH��V�ސ�>P�>	��9���[�9�+�.�E�!vPT4xeR6|�0����/o�ӑQ�_�1�g~6�?_�,:�8��$_P���[���C��a��\m���3<W�����gx�>�s�G��LØD���i�j���w�1���2�}Ӌ&Jz���}�� ��r�,ɮ������n%�ذ-������^h೩C�u�WI�)Rz	�P`M3��N���.{ Eb�������~w󢼃��_�H,E׹���6����.d�����N����Jꢬmc�f������*��}�0Cʴ(���;��\!Q���j
�����3�m�d�$�J��m��"�W��;!�ǹJ~��J�������y�!3&7���h8ߛ�{G��C
�Ѕ.�|tQ��E�w]J�ANC��FrO�&��xG/�R,�R|�E����NԜu5
��r?dː���=v��l��?�nC��9�����8�����h���q��> �:��8���>�Ҩ��Ece~�Uܰ�뫢�u���7%��eJ��iN���"�#���1����?1�=ʙ����!�7�5E��#�5���9瑃%���-�`9��e&x}O�p�%).P���DfO����6`�����{.,��HM�4 �]ɈxN��������ԋ�x�5Jc���-	�7��jR�r�^��c�sZ�\b����utȟ����EG�F��a���O�������JKi��X��B����C�z�E�[6�v�g0yX78�Lk8
.S�	�� &�����"�ô���h,|�<������%F���!���+��J���407�m���%X�qݓ�w����u��pc���3[a���4�@�idLZ�'�{^���U��Kp�r�բ��&N��v��?"�?s�=#΅ۂ0�oi���^mL�(���~!ƪbjI�R�i��$�6f�Ǘ6���$�+�Ry�W�%��7�,�?m�;�=�p���nxc_�������O��=H<�O��M�Q�6E�Ρ�<�I{�Cf����^U�rB�3|p	���~C�!��:dD90� /B$2�w��3�'�O�Wp*F��=�w�2���0��_~
���=>��x��C���$���a��{��0.a�k�������9�6�Bw��ޝޛ$��n�B�Ó�~���[I;��䴦�Z��z�.6���w.�]�<��ݮ{^��ͶZ������� C6,p�k}��l���1�t!�Fh�@j�-)�:���zЊ�J��k��${j<�;Y��m�_( �E�|2��������X��p�v�*'|����d�����pt^���{�9�8��ǳ���M�\��`~ 2W��?��j&��7���_J~�d'�?>/r�5����f[�xjJ��"*�������r����^$r���qO:Xۃ�.0>�J�~�YU?z7n;y�m猤���X�z$n����h��=������{�����6ߗ�q�L>^&�Ǥ;�A+��벰�;,f��Ѧ^�'ح��Ș9�?ėd�C%eֿR�.A���Csw_��4�3� ������!+DT���W��%��|`�C���D_9�1���b��C_�)sBꍇ�� �ԴènmF�	�B��\i�(-��:�f�Ar��!9�O��?vp[p`_�N��;����I��ǤBTo	���=��3^_ۃz6�OO�t�S�vo�����#�]>�Q͔���(����<UÃ�e�E}��	k�I����~���YyV���7�87�����?��\�)�!ّS�	����\:��3B���L��3|X֮s�]�F9�(�)�8PoͦvM~F�J>fz������_���_��P\�|C��/��v�;��1��NW�򣔷���Wn�� "�_nP�e8�	5�!o+s����,ȕB6�-��)��&��+�}��Bd%A(b�^����;�	��,���ή̢b�
x����$�Q*�O8_t��	��"@ڮ��uȁ2���SN��	_�Ad]�u��HM�4|���L�IV��1r4,����J�LK,f�$�L5��d��h���h��Q��O�� _�t�/P��Z��v��c��0�ڪ�Xby���8]B!2:���T��1�<�?�$#�����R��M�[aJ�?��=U����P~3��o�g:i=��R}j!=���qE[���ի��i�M��t�k�+�3`�R
g���!�B�~�P��R��kD���4����Fx�o�׷G^L�?�d�����|��}	�[�v	ji}b��q<k�oT��9�"[S_��҅��&����ۤi��8^-�}/�8�ϭ"���;�@@{�C�-\�Q�;�}c�p��2y���ӿ W��
�N+*���O��/7�P�3ч7��N���I����t�A���rvC���cH�+�է�숞�Z-޿%���c�B�H�e�W����}B���~�f�t��OAPP���@%�CPO�%���@�A��x�|엝d����t#�`���q¡���hP�1��߸@�9V֨$�J�B[<�Y��x��?j��f�{5�H��ܹ��7�~'��Q������̃�H�1������2	oz���C��C0�C�#[������>dvzK}���WMA���i�����|H)o��3�@B��t�}9�9{]z9- ��?Sn�K�r#����ǰ����@���֝S����o�t��F8�8���� �@��pv4p���6��:��@���$���t�����7����=j�E!��/�G�_��ӓ��$z���	���8�iM��2�@P����9�n���.ӂ��mG�w��r6���7~��D_���ȹ��"Z�=0��\�U�j<f�>��̴j�e@Մuͩ(��.U �bT�o<������. }�u_�e]A�O�W��t/@����r�p�o�"��C?#QV�y�.���Xd�����6�Ts���}^dN�i7f�ϒ�	��6���_?�[| ��w���q�����S�����x�����/�j�*�%���I�:<*��� �uX�Ci-�A� 2�
���e��(��J�Yvw���i�;C�C�.�z���$y��G�ĕ���"�S�t���Փ��=��7�P�)�2W�ӦV�đ�Q�;�D%s|��}}�
���p}!r_��?�T�/H:�w�R���r�#�-|=�63�+�g��ϗ[PtF>����g3�a|}9�j}@Kqa��	 ��^= _3�]I̊|�V���hE� V,�������0bpñ	��E�� <}̞¯�����燳1R��>w�0��I��|��ϩ��~�҂�t�V�]��f�=�̈���>�)�6�?a�:;���F���ԉ�o)h�q�:�a�Lh�z��T��\�i�0p1��J�	z�}�:�C�p�[d�v��@(�������h��U�]� �tj��DS��h;��
��F�]{";�}�����3��0k��X<��,e�� u�C�q�U�������%D��,�9L�y|���}��U	�{�S)�0�ϣ���N9�S�v��_��5h��w��V�~�pD��%
��H�E�b`��%Рi4j��ۜ��`IDOu�7q�"��"s^-�D���4��D�|�{�����p-��� �!�!Ҕ�١�	̎]Ԓ}�~������p����3��0C��bP�|Wsl���&��?j
���ՀA�M�T>�[|���xZ����Re'�L��UŁ�l���m��qW�~�`�2n{|�qC�i�{iÏ� ���-�Ԯ�=��5�$<�oM�A���#�(y�P+��K @�>��["^��ת�����N���z����_~���]�(��od�X�ܥ����M��AM�Z��û$��
�UQS�ig�=�����Q��f�u�M��Z�������&.��o~եX`L>����Q1f}�C�2�:�y�5�v~�E??7�??�|��
9�F��]gv[�YܶuF�%lȻ��=�Q[g�ѝ�9��L̾odg6�V��Nf�>�k4F�	��+	��	�������עG'���r��
C��'�y�g�L�6N5���E����.���Y�5=v)����݌���_�T�	~��r�a��Œ ��l�/�D|L���W�7� Cʮ�ы�ϴA������YX%Vf!���?I�>d�u��@��RyK��=��F��${�[��uUm/���e�W�p�{	�E��䦬�;�*����C0��4��{�4��K�&�Լ�ME��{�C��ւ�������Ǔ@�_��Q}�*�X_gI
lX�Q��%k�G�Z4��TM��@��|��vc�P{)S��^\��8�������׳h�%��e>F��W��:�]U�!Ԝ�xo1���Z����M��5�_��d�����q
����p�� >##����[�6j]�����{с�S�p�F�|B-"��!��m����
7��������+7/����]ԥcP�����KI��B:|J�-�Lқb���e���'�IM���v�����57�͜ �|�b��Nk�'�
�Vm�%u�OA	�bwh�,N��oZ����*X1¿D�♉�
K��a����ۣ�as�zn�4���0�F�&'|(��;��_�ֿp���-ȿf�UB9���v̺�ϵC\ј2�	��1{�O��\�;�UT/(-h���G}���K5���}� ʚ=u���6pSqy��:�:�D��q��A��/Eyh�Ca��_���z�9o��ࣦX%��0��B�t��=[���\��T��Y.FTq�z���y�	�!��Å]	`����7�,/�+u�Iw&�x���<��7~4���x�w)U)Z��$\�m|�w8�7O-��Zx�$kL���42<=ܨv����$�.G�G��9"KC>�ҁ�[=L5�Fw�ۜ��a��k��C�T
��/����^������3��AF�������L�I�Ęg�ͨ�׌t]e���ד��0͎�֔�[#�LZ���ܑ�}�R��3���O��wYH>y�S�����we8��r��i���Lĸ���}�U�l���v~s�Y����o�����s���;<��2[��X��HwBB�!r(�^�N� 1c2~z;�<4�H
��5�ʠ��u������B�zX��X4��=����.o�l�?����SL��f^��2J���Zf�g�[�V��q��X&���`n0Ĳ�*cG����d���~c���yիP8�;��O���nH58��w_�M��Bc���m�K�a��w�����Z'R�F]����H�c���WŒJ'���[�� ��׫�>�}�}9<�!5	���cY� H�*I��������C��S�����l�>��(ѩ̷˻�Y>��WT<������ZlPs�� e� K�:Dޮ"�bqAk�`i�7 ���8��V.��d�4Ex�4�x��E�݇p�YC�D����O5��������>Dʧ�,"]L������-H�� ��h��:��꠫������QD���Fx�O�̲ب,�f��s�9�֧��+�D�4(�o9m2�-��e�ā �[x߳v;u���o=���ۡ�o���s@����h�G5���Jt1٤�[�G/��w����SF����=���Oo�
���Q�4^�O����'ب��R�Dr�A��C,���9y
#O!g���=��awf��IPs�%�dͧ � �9���`�K�)t|�����al�z��u/���/�L�9��W���#J��S�κb��b��fe,�s��1��un+��i𽥱��[�N_N�C���}#"�22mH&n̸��S��)w�+��d�IW@]��͕T�{rR=�-�zvD����X�k�S)�œ#�r�J����#�H
� ��
7ND�_�>\g9_�.�M�;D�c�(����.6�hPI���F5�����xX,��4J<>��Ya��=�et�03��]%9ȘlƘeO]]�P����)Ƴ��/�J���7K�~�0BI�<�q4NsU��ў��1凡���;X�D|�\�,�xN���^�⍩��o�F�W� :h3����s����tN#:-��W�睢Ń�#y}�s�YC�ՠH��6է������	"ju��h$��������X��VQQЉh1E���bY��$7H?i,}�������B�dh�A��ׇCzA{,�Z6 J�V$��]
����K����}5���2���bѣ�H�  zNL�g���3;�ߘA��3T�I\��0Lw�L2�Vm��I�b�g�x�[�߃��1���!�rpa,�O��ί����M�;0IA,�u��t��Y&����E叛EyQybvƲ xR��*H�5��~G�a*��N�;�'x�X�����3Z�s04t�3b+U��](���W��4�ke�����ߪ˿I�����r�d��.���6��̶�j|�+0S1[�&^@^�h*K󶗹~��������}���K
L���w�a��b����b`��_��?ܸ�#�1>#�)���-�-���L䆼��}&r{P�`wN���Վ.�!ZV�2��i.��9t���Ė���������Ŵ6���ӳP�)�-:�e��/���>�*d��,@���Ȩ1B}�D
����~��R�Za�aaM��B,��3[˺Ȏ��� �f�u�X�p�!�ֳ�A�.ǉF��>��>���-���n�h�]���uXĀ����6�;j��I}�x��\ݧ��^Q��Z,0&����~6M�ϑ��u�o,%�?�*.�is���>��`�:�M}����u�/�.����\����$�-Ԅ�5Z[p[?~L� �#�hǂ�M83��(t�����Ģ��]@��h����Zh���F�E;�zY�o�k�z^7Yt��UQL�9���ȳ:�uA)z��׫�t�i�ư3ؚ-��ȏeM�J��o�9��
%���FJ�6b�5}�V��$������|��~��_��e����H�A�'�͓R����p2�E�X����_�S��w�X������t-���(�v��Ꝣ�$��x<]�ŏ�b�m�rsz�����
���I�?z��|���c�K��tly����&��A▥QT����<��P�.\K��������SZ*�Qk�]Eؠ��L�<GlǤ�~S)gx6�c�_�o!+2�j&zxF1+�(Jm�=�DN`'�Gi�z�3��.�uڙ����:"�$�I�P�Ȑ�h=$�@�*�vZ�I��X�i`�:��4__2�?�<��&b�Ҭ�C@�<�Q�����r�}�UC���/���:!�����__2�&<M\�H�S9ǳ��Q1��FO�KG�p��o<c,��Ix~�K�%�^.�q=��q���(�T�D�`�*��h�&_\4%��׾~�~ގ�Z�	���L?Y�j��դ�X����ٯ��̾�8d_ӛ��*�^[:�����`��!�v���z���9m%����
�!��qD4�ˡ��ВϜ�Gv>q�NF�x�"�����OΈ^s��SE��w")�{�,�2tw����ۤ�EWH��h�q�\�:�F��Z���N�,�����נ���6�Ԇ��m;�����փ1v@83�7B��F�hܶ�JV�~��,d�it���J(���Ob
4�+Mv�8\���:M���{�Y�a��w"�5�2!�.�����'�^��Y��+7�O�+�WDT��j���!}4��U	�� �z��(T3 �����Ǐ���O�J5ˌ���D�1�r��t�\����7��f-�L�#g��]πH}�(	O�y��?��}��˲��ʙY'a��,룽5 �Es����%��nu�J��n6�a!L����	�OD	|+�#�G�̈́W������X�N��艭^�幈��p"Q��~T�G��~��&�W����9c9G��9sJ,��(������X=�ޮ9����cޮh݈�>����K�I�>�b햜>~o��;�b���f�b��DR@�9��B>9<6��[h	}��J����,斢�Z�Y�,8��O��j�d��_d:�Ʃf��j�ƸU|O��:^�ȯD�K2�u�k˸!���,����Ɇ+#����E���)�D���b�������_I�K\�N�����K(��k2̍�G�Qz��;
sÄ�}�"�f�dt%ȸz�4C�<v�3�����]��Ec�?�;�2�*��O��b��/B�1�>�Coau��O��������[:u,ϸ���6���`o��N`����Tf��2��pq,	�e�Γ߿�▜2e*S�~�����~�Aک�7T�'M�ۺ�|/�.D�[x��[� F>/r��zY�w1�����H�$z���$����i5^�?���	�v�O>q�J��`���{U�VWQ��Ǵ��O���K�u�Z u��E�	EvwR5���Ba�]���A�˽����w>�����dֆy:53IN��_���}ڟ�I�>��zH��7^����Z{�#t�g�]��'t��]�A�
z�qREO(d��V�f�ދ��9�/��΄�"y�M�� ]�1ߚ@��O����v~l��ŴiQ�����w%'U��TеL�/c,<��Ѭu�4L��ܿص���s���0Qtj��MX��d�?���1Gs ��2�a�c�=\��[�[����m�_h(����Qۀ�r�m�`�jy�ϩ��L�]h���_�*7>��ɥ�-'ٕ����t$Wv!;����@�64s������$�k�q����T�f���F �WK&�'i4�5P(T���JBp9��N�c�͠�������|?Ÿ���1G]w7)�M\�&�C�hX�)���ڙq<��6��W4��M���Y��Y� �j���@����:�]�u�24���ѵ�	FW�_���y�����{����O��[����wڴNZ4v�9�Z��wuJ+��'J?��)yX�������0�����Y�H�2,�~1$O�)�(�2ƀ����:"uPy�腫�r1���h�s:�t抮�1'�}�|<-�4R̐6z�?U�4�a�@@ǘxĦ/�D�T��X�>,a�e��*�z#��_jt�r'Pá�^�}g~��h{ɤ�|�d]�ㆣ�g1�32��G�,�x�5F�>���� ��y[�S��z��XN" Dc������ʄ�K���r8"7#���Mh����jʊ�������JQ�ژ4��d�z̞�<�K�͞f�7e�%~�P�5U��:�0���ա��!�x����J���]�����%�Z+�����/��v�GR<�y+� ����R����@���Fo���f(�9��_/���ߋު���C������Ys��d��g7�&���3b�V�2W�ԺtK��KE��ߢv�%
�-�b*<�z[ݻ.�4t��`||��r�iP�_�@��v.n���?�,���s����<6�P�_�%��=E����0��K��]�.<�l��5�c�"o����g��T�����6A��(��Jn7�z��h`g+X��5pО�?I�*�RF�J=������F��y��lKea��A�,���V�=Z��R�;��A-���ӝ���'����x��:�c̼��zc5�n��l.���	~(Yiku��5J��T&��j���U�j�lAn{�hLN��!��H�F����>�1����o��ja�ւ@i]���{��TZPU�i�5�D+Yʳxvo�TNN���V��E��W>Ѐ��x����ocf[���V�	`}��1N�b9��y���bI6k�Y����1@�D��XD�\���m���'�s�O�_.Y���9�Ξp9^+�ĵ�m�	��sp<!��l��ucM��-Ct�pra�>O�n�����E����_���u+Q�4-G(tΡ̉�ɍ��H�qSv��r@��H�ĝ�E`��As턵C�#�/S&Ɋ�M �N^Y�ߏ`z�N��'r��ܡ�cr��
�^�dW��2J���?�j�/�@�l2���~󏽺��p��/�g���%}]���jz5o��~�3E�U���k��@N�o�%�];�� ͸�D_��ۏ��+�Q�Z`$��*�h*��r:)����;і-]�h�'�*�M9�jW�1?�q��T��bY@lE$yt��^�����85T<��_���w��G��C◛4?
ZշA�!H�(ٚ�aaN�@|���t; �g�k��@��hlL��4���ϫD����#^��c��i��w��L.��~�+�pTI@�Z,:fc�Q<�=��ٰ��CpӠ��%_���[ �괎v�����k�sR�v�: ĩ�,������1W�s.�&�ǵ���V�IPXh���Ug�o�0,E�=
K!O�:�ؠ;2� kM�,����i�9�����]�Jv����5���R�Z�֎f�1�7  +R��P���(��> �P��"����o����[@)�ԜeC�fq�=�n�B�/�!�O�@�rs�y�/�[�Ď���*�!0@Ww6b{�8�6:WثS+M�#``�ڥ1P�+~�d����{��!�"�����-O��\���DC�?� ٟ�g.��?�wh�${~��7��4�
��	`|��S�]lb�RA�<h��C�r�\\
�>���N��GP�tDn���Y�b�.������[�hs�Ps
����H�T1��%�K{���T#���`ĿD��%ޭ����v'^��?���
(��]�1
q�C��?��T��\��v�_M����iu�G��ؕ�8O�����	^1�Ι��i��#ȇ�]=vyhH0s������\��S�����$���Kŀw V�����{I�6�ۥK@��7�Q<��m�X@��CcQ�5��X_A�������#�
Za	� ������� ���s��� Plp��H��	�������	�����+C��f�)W�������Lk<A7����'�t`�
^f���O�n�q u3m�#kX��1�ޡ�+Q�T�=��ǈ[^39 &���R�ԣ�ј�+T�J]`�Ep�
��m���:N#����U�5lu*L��ڧ����$��/��=]1Q[��ơ
`ٚӊP'��B��g/C��m��A��k/� �K[�( �	B��+�]n|ʭ��_Q#-�����ւ�zk�����J/�%��觙��;�Nx�ap��|��P���X|qo�!�_�7��F �oW@�£�����b*��҂���h�;7,F��6�02R�=���g�|�$}�՞1�-���~��� ,��٭�3m��x�z	*�e���/7���&�Q罷Й�%�~��~b02��~�E�<CD���q���(	��	.�_ڵj��5����0+O�z{{O�_���@�'���ࡌ��Xbx�VQ)7���`h={Mb�ޚ��� �� ��C���
l��/|F��j��P��'��˼ �� �\�]#��
��K?�?��Z�ׅ-c����3�f�Ee־� ��/ML�m��0��켽\���Z.�� I0�~7��%��.�t����#�bn*p�FSp��kC|�'?�%]޿��t�^�4&8��qp��W����#��[(��� ,�&5^�,M�ߟʩ��d�T� B^[Ύݗ-԰��RԨm�$sh��͛��Br�3~��~���?�1hl�[&W�|��\=p���ϛ;:������q�?�c54�g���t얶QpTu�L��V��#]�7,���(Ȥ��P���$�y��7� 9�-��"5������b�����R�2�M��6�˚4Z��n��3$�XV!�$��M��D���P�_$�j�{4:����cx6`K�ڇt�(� @�O�u�be�qΒ{��}��JΦ>~��oB(��>\!5wH�M2�����I���Wχ��|H�S1�� m�($}�M�}�Pz�����]j6�'�"O��S(��$hM�mV�����M����P�.�ˋ����l m��e
)�4�sC�1+�ȉ�ic��S�Cb�Q��E^��m��t"0r0-�V��|}+s!rZ�\�w��]|=z�ׅ(���R*�Vw\HTff���XȢ���?Xs�n���/�B��rfʩ���Ҹ�R�U�;�h���\��OSp�ͅ��1P�Y�A����c�\��pI_��蟙D�B|k .V`	cu��3sյ�`Ǹ��m��3
����W䫏������%�'��6�Q]g��1���a�U���{2����V��:�gb�«d�_�s�����p�\b�������%��{�a���-�@g}?2�ɖ1iJҵD_�Q�O���I��SQYʅ8���k�ܬ��7��ܔ>x!g����AO�A�"4��Ǝ��R2�g��֑�E~�+ M�tKAlâ�����|��T���s_^�/.rn��M)F�3�
3�0hj�`S�p�� ��e���K�=o?ű�C[S0¶]~���0��������N��p���thh��yZkD��o��Lt����̯�s���*�r�z* MC�aP8��k7�a�pN�nk��HwQ�f!QM�����J��������vY�M��u+�3�+��zh�e��Ӕ
c�Z�c���gk�unՙ��.UF��@������#�:��f�3�\�Vv�&��}:��t��%�_�@�^�D[q��_��F@*H�~���sk�`U�A=���k��J�r���i�>�YvއW�����O��Sᘋ�ZO�*��E�{�N(��_�:�\��Tc	�=��ȧj�~޻˃š��/#E�/P7���;��� �$�FLN��u�S�ʱn����@w�B�n NZ*�!�(`�� �g[:I��t",.iX�Hn�{�A��'���\N���[��)-N"qp�?���2�`����rx�z.\
���J�k�h�wdS��6ڛ�%]�`�������X����`�r�~?s}61�� Zݏ�`c��i|iQ�����L�(�v(Es�È�(��[Da��"=��NjN3��3����j�9��yt4�إ�spG
:�_Ҹ��öcqu�R��� ���Ȣ[���ț��h��"8�ܷ(CD/9!d�<��7�C��9G�=���F�9���HgT�n:O#�ٽ�BK��ǅ�M\XB�
�X�r.6���(�϶v$�O��է�f�x�F�%���U���ñX�5x�Z���.se��e�Y�8]g:]we�'h�TAL]�7j�osp!�e��(H�~�=Z����_�P���^�ĪZ\{$@T�4~D�N�x��Oȗ
�I��ɊX	�.-�{h�T��)h�5�N����VWM���1�x�d�k0H�1���I�1�a}4�G�c�U٭�)���i����Ʉ��dɿ	�A
��:��H_��~��<�a��/�)�+5���2Yu�(SO��;l��9��b5�7m�`|������c�u����X���ϮL���ůD0iO(��ѱM�sp."Z��е����eq>.kG>��;��>l�����&b�a��X�W9�J0����7gg�/?� ��"��2����.X<O��>�8�q��_��"ߗ)�Fd�2�H`����׌�-�oɗc�:z�J.��d�F��d�G��� 㤭^��9Ҋn�j|��тN���L8B��C���D������3��G|�h�v�v<>�Ƃr�6�.��m*��������V�&��u��|�� Xb柏 �kP"��'U�?�%�g4|2�����	��}�k�ڎ��_8�	rж�#)�N�<����
L�?2{���}��|��5��Ҹ�DYk8�S��zz.���@g@�i�y���R=?M�ŞP�PW�#���e���:5��`W�G�����?M�L��x��S��#d2��Lʪ��� ���G���L�pҴ&�5̳?ͣf����x9�J6��MP��ℽwX��qA{N�OO�.�D]�����r3���;la�c$��q�T)_I�����W�1�>E;� k����9��m4ҢU�9�/�!��#y����4\`�	'������W�O$^��P�ث>3�S*��c�(�ј�K����QQ`���$��/��:���� ҳ{v��yK�a���� �H]��Y;7�<^��s=��F5���j�昴��*��c���+�F�Q�j;4�oۮ1�>6����#�ۭ��ϓ9>"ri��b������ ������Q��b�����Wg�[M�wX}� �Y�^P}���5�@+�x�C�c.��������!�B-�}⽧�ܤe9掔�v8��e������ȯ���A���W��#؇�y������י�ֈO������2AQ��{.�ǁ�ϝ����0g������ֲ�Hx�5:�n�!;��M������8�a�����f�ܨ�:B�.�Z�S�Tt���{A��ׂ!�ω;��7�o~�>j��ۓ!���s�E���e��+2"�k[��ʿ,�n��+��uT����c�����њ�C-i4p,G����2��TY�a����=�Ԛ�,���J���y _�Y����Q�Xj;d���jd&cᯅ��}�}���*�]*rJ}U��;�+����,%o٬9BͩQ���.�\�1�`���k'�Y�w�\A��+2�}[�q�G ���A�)� k�Ӛ#W�-��@�#m���ŉ��S��	;���g�78�KAN��wd�H+È��wdڶ�ʻt����o2�\W��� ���y����Q��c�1� >/��A��p�|G����D�[W#픿�r(+�����l,�<VN���#�h��rUf�g�S�� ���Ī\~ke0����\uBF�M����a�>��у9N���5�_�<��9���6��z��d{�|m��4� �P�iRʳ���ik��a|eؕ����Q������_9�DZ̊��m��#��_�$FÇ��:� r�5��9��@��x��߇1lR�ǀcJ�w��af�P!��
9��)Ky�7,5�zW�p~E6[ӊ��H�o��F��{�1)�(~�T=�ݼw���Vuė$�����ӵ��6�$u�rj�>��EB{��y�c:~[ȸa�'��C��x���L[7�j*J6�=4xHq���?�/+�%5��r������i9�H�5B3i�߬�4M�O�f�46S�n�l���ϗ�5�/�6�_�"�w��\��:`�����W.��Wn"�`ֳg+�4��YwFo��2�K{y����h���\"!�ׇ)��԰�aB��%�˒|��d����:�c�dCr�ܤj}1t�ӻ�ˇ�P�����<���{ؠ[��ܰ�����@���B�cw�����M�=���u��f�mdLnc�~���m�'�Ӓ=͒�͒]�J{;���Z_�ǱjkX�%,��Zy%��[X��X��Ɠ���3��g	sYy����z�)aʸ��"oa���xoG��Ϧ�������aCh|1�J�W���n���z�_�ǯ��:T�aXN(�F������hU"J~zH��H#cw��b��?E*X�U,�K��(��3l?KRǒ��'Q�����������nDe��$?|NI.`I�O�� �7(K@�OX��)��x2w�J+���p7K8<�Щ����{�%;ɒ��l��,̆�4�l/K�E<Y�@���%��%�7KVO�GK�"K��%�3K�\<���F��Ǉ�,�4��$��6�<���}�%?@	��΍'Lc	e	9V�M�Wht���K9K�ŒM�'�h�>e��X��X��������X��f5K��z�O��jY�o�)��,�+�dk�d�c�>b��X2_<�CZ��X�5,ٕ,Ye<�8@���.�rS��}�t��3>���t�������,Ew��a�f�v���͗�ɜC[��9F�:?��~���Ey��Gmgy���1Ϻ.�*�H�}/���F������c��.j�[�%_�SK�߯����J�0���x�fw����m>����wB;���IP�\-�=kx�S��rR>^���T�&���I��%�a_��$+�!����D�X��.�	�И}��1<k�%���#M�=65?`�T�J�2œ=�ȳ��~������m�}p�^W�sL�C��p��$�<�������}z��i��;-�~2ޟ.���	\��W�����I�"�l���^*��ޤ%~*k�y4�R.M��� }�6{)�$4s������&f��2y'���Ԉ�Y#Z��z�Go�}Z����p�7J�r'�������NI�'���mc��*L��j�:�����Us��լU�B��,�D�lF<�7)�Y��40F�;�$��p0=�{7�L��fa�5qk�
�.�y�=��IQ�N�[�����5Es��w���65�A���+�?��l\��J�ma�21��8��o8�j0��t�������-X���Y2��Q�l
H�mI���J�~`��g�job�z|}���a6W�=������X��5X~ߌ�$�Z���q���1k�X�Bl
�z�z�JH��f�"��zQ�Ml����X��35��j���J�ڼ
z��ט�c`#��@��r2*P�J�,�/�a��K^���^"��)�5!�J9'϶���Ȃi�H�n�;�������w�Qv�2�?�%<���D�3^��\��~��::�/!��Y�ςW�%����S�%l��_2W���Ks�<�R<��Y�*����ٟ��ޖ�$�].^�Yv�A�r�g.�lA�aù�tuC
r��T#�@�:[�ƚS9m�hy�@�	�=�P�90�ʪ�y��ua!�<�r��FgE�VT����)����12{k{��Z}-��`��2������W�i��W�؏��B�[8Y��~Ω,�WWr�����[첫PX�Æ�J��-ϐ"C�+���#�N���D��d﻽�.�_����}3�/��Ds��!�����u� o�{����A7N����WT"�s|pExA����RA���[�>��ݚ�Fmv�l�m��V�J�$�&fg��M�3��!�����g�.��������J�<�zc� ��FQ)Y�%/�R��S�9��m'jc�ϭ������9}kGk0�`h=b��/Ü�Fv��������+l�5�� 6��w�]�S*��wA�1_a�7u3iƯ�����d(Øi,��!��b��f�7nj<��R��.�Dxk����ཿ4�ꥮu���fR��}`
�����Hk��7��,�%��6[�I��0���6�b��b^�\r��d>�Σ
j��[όw�'އ��NaZª��y�f�T�KP�a&��{���B�(��u���*<����Н�yo��7��z^�lĞA�1�[L%����tt����&�g?3�v�+���T~�	O��t�����f���!�Es���?��B���q)-ŗ�Z\��u���r�6r� K����F�F��~ 4���0J��$,!���o;�{?�Xٴ����~�� (�(�����(� �(�^�=h�{�n�(��B�)_��ԋ����f��w����G�UV��En5P�f�C�o4��X2���e;O��������k�Q�����ˢ~�V
�z\ԟ�F�����h��A�ɤ��g����[��Xl'�Nk��G����#�Į����5'
$G�x��Z�)c|�� �#$�e��ҭoRK}<�Y��� >}:�rFuZC�E�9��k.)�uauݙD�?O�g�Fp���l�B�D������2�II��M�V��D0t�A#���l�/�܁��t��rB�l����lux����v��Z���aPէa'��e6~�ް�|0q�?�tU?z#&XV�V�Z&�w������Qif:���$����(�Ix�h����z5�C�B����z��@��D�T��)BPM���i��k&�5)��<HT�	P�҈�t�9�jB�K�H(��ٯ'�]��L��f(�e��l��6O�7I(�Ȑ�\�`k�W��fa��e�+9���v0���B󖂎�Mq<����j��u`)�5�¸��S��2����)�-���r��8e�V�d4�꟔8���ku��{�皽Z�h%��S�r����:sZ�Vd��qW�3�#�&I&�I��t�ЈU�#2F��M�X���6�oud�l�@�0���g��F1ՠ޵������$�A�;�s�x�%�\�֗�\x���_1��;��l,H.�PPX�r�s|��y��wd��h�&hC1���UG�f,��s��W�b��A�]�D�&�G�B�h6һ�i��si(�4-�镭�X<�lt����A��;1����r�Vw����դǍE%�};��R-3��*�U�z���ȃ!���R�=�2���7-���]�\��aft�
	�'cQ�Nňy�N�+��}b�	J;W�{�G�9����ӡU�0(�ۃ`����7�hjD -(Tg��aٿ1��5��j��G��8'���x��o�h|>�n��d'���3)7.z��{����S��3dƒqז��)�+��)�}dXQ�j�pWH1��9s.U�"�����qWp��3���ȁ��WO��o0�2��MiL��@l���R�e�8�_�V�!2,�ߺ����@�:���h��u�_R�w=ެ�(���4��dD�_���'h6�yσ�T6�%�Y�MN�|L������r�w�vŰ�h�4����Fv�q���%����[.D��˵q!R����K���Pp�a$\3ֲ��H�;Yԏ��~G�v�o4k�K�&>����[&���6*k�p�����Q=��8�\F�%�,��]'\����{u�JIW���-����T��ç��R�k(��3�z.���&�"~�<�3A��a���t"vA`�_��[��"��A�g��ǩ�Xķ��G&���j�#N�ɰ�؝��8ۚ� H�G��4}�hr48==�T�-"Ǌ�Z�?����W��h�﫪�xqH*�.װ�I�D����9�`}�W���e�O0@�.J�Dc/�nSm~$_�ߏ�7*��.)Š���@��m��"5��:=M'��T��o�|8�m����	��l�����E믔��5*a�&ǥ�VW�E�?6�Jq��9񥺭DwO�I
v�41��K?x��y�#�B���fEj�öo�D5o�䷃n����{W�Ș3�lؾ)> ��?���W�e{G�>����D��0����>�:��S����1�l#:�=��?鋎4C�2�'{�@��b{J:���ǵ� 3`6̟g�7ES��EaZjeE��Ĳ���J�!gdᕜ��S�n����h�������������[��-�_!�k��}Ftˮ��s�~��)Y��8
Ӣ�����R1�����Sz!��٦�}������	�g����(ښ�'/Ʋ��^���#�c���}"G����'�9l!�/����p5kQ���P�	3�x�;$��,?�,����T�&d�!�?%3>=~FA$O]M��Џ��5�]��y�X�>����
����K�͉x���Q7%���x����ￇ����<<�*���t�f�ZH$(H��$5�8�%H�N��A��F7F�!$�ݍ��,���2���>3:.AP1	����� �XE�B���snu��}��=�o�gLS۽��{�=���0S�{e�4О�/\�����8AW�gL[�ë���� ���R����;>w��y�MI�x�g��rv��3包m�umO\��'=��L늷%W���4�s���O��->�?AR���l��nNro�(4���D���'��;�3�QO���?'}L*�=��Ms�M>���稍 lzý}Ԗ#}�ޖL�O���,����Ɵ�v��g�v����8}MOL��q$�Ia�3A�ہ��i��=�L��+�O~�䙉O s<)_&���g5���?5㷿z\>��ә���+�������=���@�c٢�pzfg�H��hG5�ۂ���;�����vQ��qfo�+v�X��Q����^��l$~��߂6��+9�lj��Q;�B5�ہ�{$�[�\TOZ�Fڍ������?M�=���d�-���H}گ���qZ�z���@��k~"rdRuԍ)ɲ�>8��t?pP��Ji�}�D���+BǸH[�.�֦q����TL�\�n]�
�t�}���Y~u�l�_�- 2���svy�3�o?G���F4��NlJ��ٿ����f=�Ϫ�Ҡ��6��XT_�G"�R�w]���#��S:��*bz��h�ͶIg���H�yW�A׌�4�;3��|?�5C����j�������Z����G��|4OP� O����y�6�Z��8�l��� ~���c,���#��A�\�\�ʙ�٘�@z=�"h>������hT���-�<u�	�Ѥo���Ri����nĸG��A\�/�=�G�p7�\`]:��������������?wJ�E�����V�2C�0%���%�7NI�D��'d:6�J���Tꨏٓ|� I)��)-^�G��6XR��D9&�3���Q���O9.q?�=k`��,qF`).q�W�:�Wk2|'a�'h��.b{"�XڧR��!9M�����,B����&�"y\I$&��P��4�b�qw,n�g�������=��ՇXT�I.�H���W�|�}���^-�&h��������x:0���r3F���}�����M��|���(�B��@q<�9Ү\�?^d�F:�J%��j�����_��d�����7��X�A�3!��?=�ߥ�h�KI[Muw�IC�����Ev�
��wz��^�s8?;��nf��R�����-Us�?jX�z]?���3���1q�g�JT�5�|�5�{Y�Wٌ~-����-���`�d�0^�զ�+�� ��ʽ$���t�-f$x;��Hq�|�(-���
�%��U��*�_�i�,>R� ��WX��R?��F�XA��i�UNU�����V4d!&��>ekI�V�C���C6�SЧsʂ0|���
ֽ�IN��	�����w3Y�������Xo$�]� ��V'�#���ʕ�]I�uU50%Rd���%��������ϱe�~_on~�����/'S�J&��E�~����0����pk����X�5�/����6����%X:�/:����pcj�7kLvQ	��_�ߢ��,LY�:�Dq��׏��5kY�R<��o���+,Ơ�y�٭;�<��A�>��˺/���)�a���T�!i��p��hR���%EF;�|�Mj �r�U�pG��^b�\DK�{<�F����tBȷ�O��bKq5buP+���M	�s�n�B�,L���E��߻Z��.���,Q�/&5�3E����+�p����2���d�C���;-�p�j���(��#4w��[F%�W9Mj�Q�|�w�q_�?��W $�3���,����aN钴��y|#`ݷ���̋�4��C��/u�`t��������×6��g�V�)}�=q��>�H��Tw쌇oÇ���TbQt�bƧ����i9@�/}��K�i�E���?d}����7هw�`��2C �.u
�0�ݹ�fL?.����������0���kK����0B�kJrv�Rڲ�k��%�S�mX�g�irD�:.�ݔ��]o.�F�V���3��B�F����'F�$�'iB^����#�j�u�ʢ�0����~�D�S�^�>Z��^ˆ�|�n�u�C�3��LY��R�J_�.�4
>���
W�bE쟡 *C_��b�m2I�j�B��ɐB1K�\ɽ4T��	k��S��H�T�TȦg0�ϊ���&���'|�A��m�$���;\ƂXR��.�p:�x�!(U�R����7D����W��$7�C8M�x�`�3K��:�|xF)�A�i�����#���>�Y��[��Wb,��X��!����������8�TRK2}�My8�|4WR�s�%t}��T/�Fi6ȼ���/��>����xE�9ف��`Ad�y6%��L�÷R�������������y�͇ۛ�E\q\_N^���c��D����b~5��D�p
8�^��IC�D�^�ǽ��BŇ���B.��̮nr��I;A?�U��2�'��撊f�@5�#�l}�U>��)%1#�U:V�-Ix�Яr����&���Y�o�!��O�!*�
|ʏZ!�*��R^T��p��Z��u�q|����#�V1�H*�cKIP���9�����&n�g?�ѩ?��f�ɇK����0��r��ίm������͊<���R�9?�v:�
�+�a�@l��/����>>�m2�4Km��;Ms���\��UK���0�O#���G���(ԟ�X����*�ë�ʭNW+֢�5~gŝ�{P�d�HyX2��G1O�͇�w�b\�^z�/�C�RTN&r���l�SjU� :�Ђ,�&q�)�)w/���C��x5��P��| `���u������"[�S��ü�v�:=���Ç��-���Z�a'�;��}���o;����W�����dl��ak��q����2k��f`��V����� �P�9�a�W~���T>a~gc�e @9��_%d'��Zm����e��bns�&���)pI҄��b�NP��pѿ:�eFzO��IO�?�^0�����ls7B;X7g��ɘin��"[�M�R[Ưܕ-*K��v%��y�壜ِq����pf�-�]��'�� 2� BŉL���qU��Z�j��8[١��o3�_ь����+�f�c�u�R�v����9:��d��Wa�| � 귁��5��^��z�(�k��:��>j���SJF����m�/��y?u1��:x��*����O�����I��7j��oIѷf�;�f�EThI+�p�5�6����K :`u�Z+�K���);/
|�l���?��X/j��Y�>�$���<FC��?�g�}+�����I�w�G�vǬO[��8�OՙH���/$4���gD:�Z�8}JnVB����u����|�����'z�?韋~��%�>��dj�Vp�_i��_�G9��>_b����v��uR���M��Xȼ��
\ �л�}(�'�;�y���Z<&l�=��>�U�T���H���K8�&��Ѹ���H��[$��3��r�ա�]P�D`�g��������kC�)ӗ�`�����[�ݜO7O�o��h%C�L �Bʿҥk�h�-p���&,,���_�5]�h~@9��Ǔ�Ԇ7����f��S�Z�h��s�G��9��~����?b��cIz�@(�xW���[��8^&�/��@��?��d���[�'21�jbe��� �_�B��+)	��<�;������ ���?\_�)��8�?/�j�������Cq;_���+���� >�`rW��Z��=���+�%Ζ�4ƕ3�6��.�b��>�� �2� ��hKK1�OM|�P>X�T�Oq�O�b@r��0����X�����A� ��?�M�M��>��I:��;�c�<���Z�~(�%�֥㌣��&yi���v.r8ĺ�"E|}�{g�8���<��@05�^�ǏM��pˊ��1�8�'a��3��]x�"��9xq�&}:u��֓����`��!M�.tj������~��3�_cD�w=jl�����ut�lfB��_�����>���}}���A�w�~!5۔@&�x�<`�#ٙsV<n8��{�,������$����xȦ�ǘi��L�9J@����ywL�d�ly�V��ٟ���;��ȐL��{;AÈ>��]���ίN�e8ү:�'��>%CR~���PI/s�7c��Y�6�e����b�SR�A������[$�L!݆߈�����^��>��I��+�?ts0�T�O�X����m�j�;�y�{�D�)��2�>���N���c!;�F��;N�xyV.�>KO��"�k����:�]�
�B�pSwwI�����󢳩�H/��Y
}�d�=&U�N�����%�I}���a��S"@���T�x+���b"������C�׶|���ա�cLM�`6��l�d��\"�D�+J��\��,��r�G�f�Es�O��<�I	����FQ:覓�I�� eE�Ͻ�����?� *],(��՘�F-����ц`��籲�=��絙�{m��^2���@�'��n2t'�,�k��@�bխk���D�L!�q���/śa�:�nI��V�2�A?�;K$et|�jsu�$P�H�6#�QI�Ds� �*2��}-ŴZ	���a�#79�Ӥ����my�p���W����V��o���{b��YP�d
��Uvġ"�Y1�nl��Xy�pu�
L5�;���&[��,��QR��X�9=��6u Jc�'O���䫲��M4�3��#��J���@]h4��i�0�T�������HR}��@uY	1K6��C]�Tb)���I��2�8�$ߊJ"&���f m�T�*���7��*���:JTO6��$����_�d%G�rVE�)���ڸ�p�����	��}B�K���v�]N��:;ky��_M*�h((:hb1e*����]�����s!���c#���yT��9A��쥜FV�帔B�V���I�n�>l����c4�JXԳQ�\�6�Pe_�s~�s	��!V�	_��"ry��;yqv�l��l���+�P��6?�1�o�38�W./ڌ���E�^:�����05}��D٢|��[��S$�b%@�f}Iy,걊Z9'O�
D���5���O[�clpz�쀸�	��dw_��,M8�Q�W��n��ti�|��v$�`��է����Κ��s������.w\�|���X>��G/è����>;���d�B��%���rL�t�@]�G� I8� �Ig���zK2t#(`f)�<�;�������qV���`L#��4��t6۲��!��YĦ��f�"z��f��L�3)<��Q=�{�&�{�~�Ϥ5�����|��o����[?Ic��"Ԙ��nK��W�+�$�5d�A��V�������ګ[
�د��*rrL�3k$���g���S}���44�'5L�XL���V@t����Yݐ��&�v��D�,zl�}'A������>�3~s����5��:@����&^�dg�����Q>�2Ag�{�ש����e�S7�>�,�E\��:\�EN8�M1�Щ�9��J���o�S���3��k����d�W���!�;���,�>��d/�%���+{b�g�)Bםa��*�&a�Tq�_k8�{�Le��x��V+��rG��{������G}�l�l�����T[�tM���RZE0Q R�P���+���l�wfu�t�����k��P�',����׫�#�((ήI��|����?����>�&�����#�+���W`���M�D�lTor|#�TiB<B����+z�)�1����%I�ʧ|H�l���vR��a��t5�b�:?�\0�Z�(z!��B�碣X��V�����\�s|J��>�UN�-����]�bN����9�?��h���J^0��� r��G���s7�;h���A�5M��綛v_��J/~��n�D����-	�@>��#��C�a�S��óV+�Z<�C���>��n�R�&�8�R���z��)��za����p����-���$OR�:��T��y��\��������2�r���������K*v�b�mC���>��VQ9�k�n���K"�ZG@�)��U����}��z{��X�K$iw3�9�&�j�Ţ�`Q����E�s�v�T�]J������-��N�t�R�_��S��jJ���t?�8�m�Tàp��3Y�}5|CT��v5��2���(
L�XN������!l8�ʶ��2Ē'?0���<��V��z������q�6�@̊����u��u�1�� �2����=#���.w�a�y^E31���?D�XۓdFW�lb�}h!��J��`!RƮ�?0��b�o�$2�.vc�y#5�ގ7B������;Q�?�j���~�A���f*�j��í��_ȭ�k�*�����N��)N��:K�RA�$$�>4e������i�@z��� ����t���O�I���d�e�p�>{Ȣ�U��o�-2�
 ���	4��q�X`*�d��U{㛔�b���;T��6)��+��r��#��0-���W�Z�`%����ֳ��?�}=.��VR٣=�'���W�����Vr�:Q���v�o�� ׽�6 ,
�z��<J%e�?D���Xz���q@\����r�΂��9���J]�yX"���'�z�B����Mf���6�B��]���u(a��]����D1�p.�����u��M}��Ś���Ա��/�`�3`��E*E�J�t�FG�+������;���u_�����;&K$�ovx|�-�h��p������rEedG,gu�n=ǉ�v���TOk<5��+5g���4,��^��U�*�����XX�6Z�q�&	-�%p�z�p3Z���ގ���;I?I��x�_��a;���|xmF�T��ڂ)��k�(Չ��n��Fo{�fSL�c�$��y���W���lh�.����-��u������ù�Z��p�RYneOI�^����+����wWp���m�6l��/:ű3�`�_�R~������)k�Mr0������.cf�5�;'ϗ*0 ޏx��B����n�[�f����z�����H���%#Q�N���o���6���\���W���z^�~��]~�ݩ����΃�/����ů`��&���xD%����3U�7��䴛R�Z�f�;�Uv��B��ƃ6�ދ��m^+��"��f���6���E�"��'=�*��7L��#`$�5�P }4hȇ�� z}_{�|��d ��KM�9|Tp�l+����-�L�!$ś\���n)�,� l�L�U\~a��%�2l_h?>nbc��;5�|d�R>��m�H�̏�1P�t|�����|�:Zpq࠱��ae����<\a��B�0�@ѳ�Z��7wǰ�4�O��r�I @��a�޹�tf�)�vG
����p!KAq��,v>��X�k"Ѯ>�B�56Z ����ٮy��F'쪞�y=����.�B=X��2��-RGѪ�Fv�N��[�Q��B������$��0�2��/�q<�3��� �S��*j<�Y-&l���I�AX��]�ܓm��=���iڼ\"B#�,v処���r��x�>��������ȋ���?��e��;�#�a��`f�T��Q��;Ez���&������L� Y�K��8t1hR�|�J�K샏�s�pu�r�Y p�;�4{)�7j��N���A^�.�ue��P�)i��#�ٜ-��L�>�؜���4�fBP><�-Q꟭�Q�F��W�DX\(�����uc\�q�t�����3�'mj#r=Z���M�"�6�JxM_x�w�'��W�i���\�G�1������n�#sC
Ҷ�x���)��#`]|������w���({�o/������$[{��|�S>�/9N'��zɟ^�����";�\k����A�*����-X���l���Īۂ���G�����/���c7��/y�U�M�b~n�W9=���Ef��p�&xX�RD�Gn;:E���K)�����p冩��P�Z���'r_cTm��Ў�v�l<�� �4���t��l��#F����/^���p>�By���l7��h����~a��`��3�_��,Cy���E�(�&���q �+ˈ�?���o�f�-ӫ;_�������q���������������῜�����!I��vIa)(�Si%�C���;K�&I�?<�}EZ�����k�>�C�<e�ƙ$?ǯKuuT*��z�6�Z�=�������+���>��=+��'��8�����NěZdfM�L����<4�+��Hg7�P�7+���A���ؙ�T�ت���ż��WД���y����>L���4%��]4�'��#%�q��ծ;�u���͢j[��N;���f�.Xo3��In���Xz�,��I�U���T�<j
�����	�)��5JSc׸�1e.��8��Q��Rv��Y!%thPIE��S�p�r��)�#^ԟ;��b���9�N�y]�T�+��ųf�vǌ��&���X)#����`��E;lT��Zc;�f���Ok��|c�hz�b�S���r?}���5��<P��î�S��p�Xғ����ϰ|�� �:�Je����>�^K-���7A!�?O6�L�DEƃ��c���r� 0�4�~<i|��/��Oz|��T�������#m�(s�����W?֍��xiD������)gg@��V�!��2�*��2�>X�0�B7�%�3i�؃8��i��������t_Ґx2�I�����fxYC�,/�#��/l�Ն����V��A���Ԇ0�.ܠ�u*��$���H[5���������-�Dc9WG�,ƃ�q��zy�9v ��$�l�r�gW`|�G��.x�N��(.�Tc7����.Qi�v�S�&�Iȡ	�[��Cø!p7"
����x��`2��T4��9�sj�hGN��ͪ�&�Ө�:���ȡP�T6�G�h)<�m���oAM��6���/�tEb����Ո�@5��8i��o��_b�9����~ܸO�'��ʾ�.d�[����-��B�9w����1<�^��O�z4���oQNPW-�O���qn�{��wE�s�1I��*8�<) �`PHh��a	���������(��f��V�yGc����m���5E:y�-�խ�eC��i��������6�|�u� �;6[z\�Ǟ}G*��0���Ĭ��V�����X�r����)�c����ߪx��VƿN5��ßij�]�g���;���~�/΁��xJ��z�7~���?��/�e@�U$�o��I�͙����Y�j·�����u��� ��$sU�{2��'m���\y|h�#:&9>z�I��Q|D%���V[�R��'�N'����'���v��P�2kLFm�Z�+���R�r8n.LK10=��*�P��ѯ:���!
=�x�w�ja�/�o��-�d�Z
�Y��5��RΞ��\��8D�%o:	�k)���S�ٟ\���q��&�����k�@� ���ӈP�Pd���d� �F�y��B{���veW�a�h����l�|%x����Ar��ԧX��$KL�PT�oH����ӡ�a�(*ց9-ˡ;�o;@+���[�����^	�F�|��+���B�MR�Ly�:3�]:�A^T�8=^Lis5lR�p��p�-�S=dI��خ���N?��h ^�S��z�K*���}5�r�zC�_�
O`Փ'����Kto����#-�{�^�ȍxb<%�r̿��طrZ��$���W#@�_�y�vW���^G��b-J3Wf�Ď���7���lc�pv��¯��z�5\=Q���i/HP� �,��d�&q�}��8?��ڄ�'��Q��¹�lì���������U��ᾬW|d�)2Jh"�8hڟ���^��ro
S�Pj(���
��gg3��"����50ժ���Z����R4�8D���Y|s�Y��؛ƺ�}"��e�EG��9/ԙ*�+��x�L9_-�C�ޣ�2���L�b��Ϣ�4��Y�>��.	 Q��Ŵ���?�&B�9�<�끿��k��j��������ݏL�H<ؽʇVRS*��~�$n.aއ��l
�0^�ܸ'D�ެ<Q}w�_���G�Zĕ�Ã���Q�-���RV@��~e�%��O"{���ߔ���</T��Q��|�j��r��~`̃��Y��"��;o'V�/Rc	J*�ܟ���}f��8u��!K��3X^Z2q.����`�P�F���$�x���Z�?5I�<��|t`�ߵD�#��q��F�v��_�(�r�/�n'G\v�I{O/�&J��9$�P��h73���=��k����7E�R�,][��l��\���%��%ڌ�Lm�]Q}�Z�x�<o����F>)�:c��X���R�N?�=�J+]�V�?"�i�1D7�w>J{�Y��4��5hj��w�w���u��Ry/+�7���q�.+�
���U��Jb>h�u-���,e�C6Qy ȿ7D�>��M�^r����gdX��d��&�XN��`^����5�G~���Nve����������$"jH��2��"8���e�arͭ��l�LG��L�?�/�Wǻ ��ܕ
�'��� �C�ZșsR�(F�,cgm�y��~u�Z��!�ɶ�X��S�1`�E�=1��D����ff���နh�����f�?
����ȴ�Y�{H���R�&g����*�Z�I<�h�ސ?���ԏ���˘���0Cf��r�+Ƈ{q��S��J�jq�Ͻ�9DuyV��°�SN̯a.\�����p(2��*�W���HX�p�SqyB�b$�oG��N>�:6��u����X�UJ)^�� �7~ ��"�^��!�i���S�aLW�#ӘR~�����=!��x�R<��A՜�k`~t��mZ�R"��o7�ow*M�icO/�?�	)�x��M�^�	2�;����a��)�y�Iݰ���H+{<$�+O{��`A���x։X��6:��&�̆�}!�*�~�ZA�n�Z�Y��Q��n�U���^i'I���̓f fŃ���y]1!67��d��!>����+F���3�od�n��õN��U�#�O�Iįq��X:?���1�<�'PX=���ir����B�����6K���{�Y*�J;H{�&Z(�Ճ�eG_3"q�,�zSV��_��Xm����uv�+&>��Ͷr̓�?���x-��`!`�������t�{#�)�`�Kz#���R/3J{��g���>b��S�Q�B�@�,�������f�m�`��\�ҵ|���Q7uz��lb��Ax�8c�ǭ���_��)����W�����%���=�眎�ܲ`1l�0$�����<�t�#��7��TRW� ���z�`KI�і�vlׯ��l���,ÊP!]�b��}�Y�7�3U�
�E.1��xj6�'�>��8ģ-r ��p������(�#����(�m�ג6w�kY j�&�k���Gn��(�g�"��������4K��>�"�	���ӹ����f�|ǁ8S�����X�!RG'�{(*E�_�	���-��f>�L�d�W�p���XA�?!�Py������������������]8��u��<�'PzE��clœ=o�Q4#e����Kg�)�lgiɳ���5��`3��#��sﰣ��Ex�����f$�0�j_�)�9�9����0S��LG�rD$9�XJ�>�V6ШzIm,�đf�K7�'P¥��8�J�Lƥ-�бb�B%�C"�^]bҏA��	o�Ho	V���s������Gu�b�QU����d_�P38m��C��|	7i)}�ɧz?_��� �^�@T��|�B�f����b����|���L
+l�\d�'t?��M�3Li6^˘GԃuSI9�G~��@%t`6�<Z����A�ɭ���l/�.�؝Qp�����gQl'զ��+/X�v'v�m�tǢ�a�J�Ŭy*k�%Vg���No��|���_*�Y�D�&n��Q�"ϙ.�!8|,��h���E�EiA��X7M=���,��fa�?�X#�1�v��O�
�����m��p��~��\����o�X��f��l�����I�7v�z���3��R���2��C��d�7�x8�������+�C]�@_�սM�.sX�����C��)N��e�ymFI�C�����tU��	����=���v���]��h��b�HŉN�K��e�ܒ+��Yi���{8>�vqr ��qK�)�L?����P�&�T�=�=�ݣ�4Vx/���0�j��MY7����|�ST�+-��\����1,��7��#�w璭 O�ȅָ�A�V�V�ӑP�|��m��'�*6��W�V����Ija�_�p�R�%O��Hw��
~��N�� ���	1��M;��	���Z	�m����J�KYVŇ���uF���Yw�p��t�8#nh��e�X����Y[x�i� "�L*~�VQί���v��q��)�q��~��1p[iD�L3�J)��I��|�j�A�e�\t5'MZ�ǂ#����P37IΒ�����L� P�����,�%�����?����X.�KƄm����O�T��̂t�Y�Ź|OG��W5�+Ź��P�?���p����uؽ��y68`L/�CIꖏu���EK�͇)f!_P�T֝��Vz4Эy��`��X��)2+9�1�HP3P� ��������ô2Ӝ��|�n��;��X+�D �f�Ǹ�Z����*���ۨ��q3jE����42�X���C���=�?�ǧ	q�_@�G#(���� �e��f�WJ]��?��v,U�5w��e�"�ßlE�C߽3��1j�gjq&�� �L��h6ƿ	L�������T�	���c5�.q�@��E���
КOF�0��~fm�|>��YM%������hO\1Σ^-+�JE1�}2a��cA �����J�����ju�,G�'�:}��z0+`Q��g�E´}8Չ�-����$���=�i�Z�$��I��S��0���%-�=z�������g����I���a��gӃ{���'Q@�:!|���p�3���ߤ��{S����-�"��3o�4�_E�R?�E�s��L�x��-������8G)�m.LK5O�P�p�=�}�?V�	�	�X�t^�O�7��#�W�\�E�M��[�o����������N��Z]\6�x��0�"l9��G!��܂T9��[�"�����{�h��~WY�Qc���� 
e�>�{�����t�t@ɷ�"�:MRgf�+h��^A�(,
!çr�M�����u�_~�����G|C���^���>�bA�u��� �|���g�9��g�:6*����309D�!i
6��=�D"�*CUWp�͸������\������bE��}z��!�L{P��<�<��8�(�g�/f��XCh1�9����Oݱ�ɨ����h��>�����z�Ǔ��V� ���Eì9-�z��U_@����*���\����ԻὒE���l�#�I��_K�R� �ݾ�&�ZeFЮȷ액;/}_-�g%E����EYq*|�j�%�,Y)�0k�����E	�pf��XBK +��#�^4����`ޗ�HBQ�6T~韥O��g1���͞a�V(5�X6H�U��;/��!�/K��|��p��
�8��_z���B��J�I�e@�kբ\h�jP���?�
?���sG�B>p���P�C&�B��� ���<��B���~�(k.���A�wYL�g4�ҷ�oP9�����GwG�aaWtAK�yى��O���A�.Z�ޠ-y��	cє<C��)5J"Os�|���Srw�܋q�8�`E3O�����$�&k��u XS"ú��SU���<��������+!�<�J#ˏ�TbY�oQ�Hwݟ����$J���T��>��3I/����m�NU� H�ƝO�vv�V��E�M�����'W;H�$�`���x��<>��|�<2�4����C\����߂��(�-��ɗ����X��b��o���O���W�	p|�U��(���W�������/6��	&
z8<9@1�:�K��E����<��sB�+�w�nD �)�>ŖŇ��>e~&_�x���H��%2ri	';�)z���A�G^&�������)�d�Y7��w�;�����B��X��	=�V\����^id C����q����P�֟D��y��ݾB�bU��*��C!L猵I���h�U��f�ky
x�&��Ie��d"+�M�B��;�pW�S��4��S��l
����#����ͻ��8�V*
U@e"x��b'�l�������dJKb}D��7�ϟ�޿����	�Xqw��W_<���	��/-��ڧS��4��An�w�ٓ��8GИ"�.��3W�O����f�	i�ԇà�ق�$�D���謦� @b�R�r�+^�ү�A+,X�c��_��:Q{���B_a	阚��M�F»����"'�*m�s�Y�E����q�w>�S��*i?o[�4x��c�w�$|����H����l�菬�I���4I��=9Q�͚c�D��4�˧�uKX�����||��|sS���\�f$�ޫ�^s�#�q�D�:>��a�Q�_��'�j����q�?M�<N�<R%�n�����-��)�N�W��3�P�l����C	�KĈ��M��ԕ�\�'���8�
Y��e�Zm��3u��ɽ�v{L�5��YT��xAm�Ĝ�Dw��W�Ɣ-^�V��i��]�V!�)��ˀ۲���ژ_��#H/L�~��������j�n�$#��+_����X��x���"��&�a�~zF��ie/t���Bg���A�p���`�~��U����?֓(XHo���M:S��L���B	�ҟP�ї�����3��&:�A�u�Ýz���E��G�L��"����M4:� ���מG���5-�z4��R���!)ׁ}�|F��9`�$�ey���B�de��u��;����Ns(W���+SK%�E�	\�&J��d�[koH��Qq!��!T��c��+�I���'W���ʬ��*�z 	ߩ��q~�t������I��: �.E����EQ�Mܰ��?��^Q�z�44����������*��˿�x�7y�VfB���$��^$Hb��#;��b�4o�\�@f:�f 2{��R�Ub� y�:�*�ߦ̡�}�8��PƢ  ے�����n��O�_��ho,qQ��7���뽫zc�]g��<�����!.�_?6�2վ1���ڭ��� �5�Wց0�j��\��Ν��N�
{�0D��'�Z�� ;�w�w�;D�&��=�ࡹR(�!E�c�ѭQ:d�7�ȹ��!���c���u��GŦ>��M� P�T=�� �A��g��Mz��~$�)���7+?y�N	ɋ���:h�$���g�	�[D$���a3�O�Xw/���@�Z
��=}�a���>}OI�`ZX�!��g`�SO~�|%��j�o��|}L�G�%��|����c���7���j�����t�, ������C��߲V@w���`\�-xO9��x}���b��\��=?���P�Q��i��$ef�۸kib$e������M���K�m����Z4���:�"��gݖ_j����c�*�hR/�`Q��O��t[<�@?]K�6����`3�2�v��B]	AT�Q���#jJ���'����� xWNm}UtN��[�k�F��E, �SZ�ŽJ������ך#�=��C�S���&����Ӡ����`�����/M���R~�g���v:*qZL1�M/!.&�&�>=��>�lR{���݉�<�:��*h���8'�.4��x�1x[�ťi�1��׵�iN�E���5ח.�������6>�"-}���V�ie*Z�|tI�X��"�V&���x�������w~K�n���� bS��-�Pb�B�P��_���%_���<���HoL�U
���Հ���M��y'*[
�,lqU��U��X�hx��~�P�.%�S���`�����o%���I@B��\XNݪ�u�-��O@r>rJ�o��������x���v���L��*�����sE	�f�_4�#дOA����a�e�AImIe�h2˹:�y٬���,?������	N�父%�]*杌n���(
t�!({D3�Q4S���X�CƐ������I�'{{�^B�\����1�.�^Ow$��CO�[k��|/&�/uā�SE�.[�j<����҉�)�6^���e�3Pp�k�-�=��=�Zfg����rG#d4+������ɦ��NI�(VYC�����C�C�Pk��`��u�i�y�.���D���e|P}H���� yk���&� e��G�L�%�`��_�X{q�L�s��>�uǎP4A�+`s�Sl�z$;&��]r�B����_6.>����}������Q�:���|��5���������O�(�x�
�nc,���-��xWG���V2�Ǳ �|�g���̓Z�Y[-s^fc��̉�c��G�%.��p�f��Y��[�i��4�8�_c���u�!W���Aǘ,`�V�ʯ'`���W�~e��T>+[��+�2+̆	*�8��(�X^��}�YF��*���~���R�^��pV6���A�U�B5����vڋA.p����4v����I�6��c1*Om&-�;6a�.�*v<�	!��2_�tro�MW3����k���P9P����!��q�V�����͎��5s��?fg�*��ë.��f=F눕��RD����R����V~���)�f�E�3�ӇF�L���X��M����,�p+n�icЌ���E�M�,���^�j�6unv���5w�"� �&�������,@��#�{ǯS�;w�-f��#����+Xe��q���"6㼱'1rR�V/��0���6�yi�cYo"Y��޺�i&�N���Ӹ��l=y�_�6#��j��Y�E>l������U��W���}�S&��(�1A�����>RA���X��J��I0�J�9�Z�)%}�A;W�b��UE1�I����-���t`+�~��='@�Ojf�� W�=�]Σ��C28�l�k�,p�5�]�B�j�5s�3OK�~I=����e�\�i��&�j�ϋ5u�^pJw���(�3l��~s����:n�H�U5pe�T��=!j�z/���Ye�(:�߯�#z�-�+�s�|�'�s���`�.��v�%��}cm��1x����b�U����d�٣b�_;w雯��Oؔ8���=����am<���� �]�I�(�X�����ѷ��ƃ��Mz|��
�1�ޭiœ��RW�<ן&�e[%��m�S�kkA���
"\��SR���6擦c':FT�@�ܻ�z����f�U2&�.�DP>�$Ni�k�'�u�6l��:�깢�mI��!��U�+�B�&4�N�{� 7�Tm�����W�	9+z�hS�O{5�7G��R"O��9��n�G�")��	iPe���/*\Nή8�}������=�������F�ˏђe�l��E��������v:2��C�ݧ�_L���0������>�o��6�o�̞�u�2TCY���zl`;˧�� �ΏS(N�`/-vL�I�>eD|�?tcD����~U�zg����������&���l7`��uY6��T=�lOKn�(����U�=#�h��n}�3��q1���I�Y�S��,��(�
�Wr~Do��ʃ�.}�n���+��d믳b�2~O�޹�=~�2��>�����Sn���P��=�c�<��@U��U,e�
�*2W�

I�E�R�x��4�T�|�u'}avV��L(-�(E�����Y�|Ò�͢��ɚƞN�^|@Xy����f��<����%���� �Z�"I��T��VS1��aIx�ޟ5��|gf����w��y�e���I")i�2Ԣ�F�Q[���]�\8�k.����/+���{ͅ����2�Ge���C�[o���!���;�rBWz70�0C��zA�)_�~��p"��"�ၞ�Q�os�8�,���_Y���Ł������-���\��|��קQ�c?l�_�\�*��	�VTZ�'-TTX9&(������wK��H�*O-* ��_�S�z����
pk(��y��~�Qt�C�c��X}F�l9;�4�#�u���'j�IQ<_T�Ӊ���uxp��F�	!��OwuD/��s5�	��a�w�|'����t���u悇�$߁e��k�5�Z`�W�@4����ї����8��â��$�u�p)����d���c���%����8���eU���|�kW�U8�"D���M�Ň�'����ތ����і�5����8�\q �R�a����"�V����c�]J���/��/z�����1�zB<��"Er��5�"1�)���/�7s�G�>9�j"�>�&���R�V��Iг+��K�B[�C�V��v�� :�s�uű�V�t�)z,�8?�pnr����g(n���H�Ξ�#��lE�<������3�����m�Z��Fj���.�s�e�Z�����Z�
�0�Jvs�BV�3���-���ނ�����W�~	�ÁU�3�:��Nr�s|�(-�����vc�,P�\~L�����^�<R��t���p��(�Y�ᜥ��v��u�`-M�-���)�t�E~W��nܓo�|�"GD� 4�ǳ��*�������*I�F�Bk�+�zª�\��S
4��t��;Z�H����Y"f� ����ZJ��4���p��~��/��E����U�݇���1�zu�>n;����^�S
�p"Pz����+C#�����R�p4��%c�(��\��9�|ZI�����I����H��{� u�ӫ)�TK��T3�߯��7�0���`a�@���v<8�=����x|?��|x&5[�{�c{Bh�/�:�K[9"��sQ3t
 ;�t+n����#���2�*/����?��U.��7MT:ŜqR5|�O�'�utL���00�� \��%��H�J�DA�N$��[a<^4.x�����(l���qQ�!*�-�c,��x0U8���M�ve��/����ƃ�Jez6��*W�
Z`+\���mL3�6�]b��Z���u�~�B�t������
::Kn?D	j5S�����b�Bs���i3$�m�7�:�F�<T�`c�fo����-'�xA��f��3�i��$�_9E�����9>�^`uQXH�+ͧ�8 "儶�0���$�z̱�(������w���c���v�+�`�����~l�����aѥ��ю���A��1[���1��N>򜙺*Q����������f̵���Y��]K�a0\�h��S�]{�=޵�Tu�r�|��C��߉q�j��J��F{7�w�|�p^����O�u��n\���s�o���mU�����)����5�OC�:V�~m��P��)H��<��[����3���B�_]�A�%�ݯ�I���+�H\7��D��})E���mgH�F��:���]��X�1g�Y������2�9��^���B�[�]� ���A�P"f������Q8�F�ʇ����6����䏮vAi,V��zA9G�"=��T[_��p"L�C>��ZjH�h��BQQ���R]K1ۆ�}ϑ����d9_é�,� /�4��z���_� DPUl�	���봴kA���|N'r^����)?_��� *�[��y��8#�Eͬ�W�9+������I���gįk���c�KBN�_�O���D��hG���7`G���[��]:U\~���(��.ڪ�<��j�E�J�����0џ.D/aste|ď����g����1�+f��g/R�0�d����� 5�p6�5k�&�gZ��b�V��5��<�=�����j��_����PT;����xDj��ԙ�*q{�:IE��y'A�5���"�@�֊X�dvV�+�/���x���G[
g��(c��lm����X��l���>��nR��H4��YI������ϺCI߉Wgg�M����_)N��5�r����S��Uw��;^�z��<4K//��W�%��xOp�|+z�(3�eS�|vBw,��6�>(��<rapY������_H��x�NO�UY����r��t�Tn.,G�V��!X1ﴩ�o�G����y1؜�0�X��ͧ�0C��ٮ����y������
�9�v�_8A���,� �� ��b�9�J�qP�[%�i�{X��c>�rs��z]Gp\��
��*7���͜~��X��9����\����x���C>���0�����f|I�U�w7ʃ#m�E�f��c������y_��Gx�k��D|p��/*���_�;����"��.t"F�|����v_�w�ds���+`'Jڳ��Ԟ<ޡBh��X������XRt�+R��H{�D�>��&��h��b�������2ϯw�MYQ�Ժ�a!Q|��%?#��	���;�^)��1C:6O������r7
��f�=N����.~��%�/��<�N��`/S��15�H�y���O�`�qv���ihv&���hI�OQJ�AZL[�R\�;wQ0����_}1�T =/:މ�<k}�LI�O�� ? ޗՀ����w�:
s��9��;����[ԇ�]푎�B���E�����_�|2��.uZ��.*�^�V_�ɸ���Pv����b#�$��K���`�]�٧��J�++0G�Wj	eВ�8�Pf�'|��Ljp�K`���h���'xj!�I��5ȣ���Z4���Q>6\��'F�B�~T�g6��י��#���1tb~���A@Fs�a����A�:)�_W��I��O��B]� /�f��ԛ�A7H07���J9j5���6���h��[�N��|��h�����o5#��)����%�������IB+���'_���Q�Dq9_O�P��>ӂ{�_wψP;�|����A)�����F\u��rᆪQ�C5|}C�A\#WC����#�0���z�����%��:��W��`���SQ������=r��`Q�!�6�oJ<j��9�1{�T�b��+����<ȜX��W|+lk��w{�ϳ]�p�k�_JO���9����_����Yi CJ)���V�~H~���r�CM4�-����+���9�h�+�e��y �iQ1@N!�?����0+q�(���V����p�v`�eA4��DE'�� V--m�[@L#��ˋ"2��waLQq>I����z�WP���o�:��y/Z�������TR7ff��M|�mL�"/ǋ���k�z�+��m&��6��c��-X�x�0ɸ�ǌQ�4��?�b�F2$�=,'�L���n�!�ٞ���VQ�c�ȯ��%�rV|.�V�K�O5V^<�UJ��0�,�"���9,unX�V�4�����w|�����4�� ��K7�/�M���XI©��WB]H��$&�����8��X/��T4�+�E&@�D��pA�R(��pu\N"�M�B�N��7Ӄُ��Î�Xb���<�To���턶_�I*'�3�Y�q\�� 
ߍ�-�/�5��������H���?AE�qn�TS�-�k��Uʖ�F��~��@��,pD�v�BƔt"�y���t´��?u�*�4<�S��qX ��8��w1�m딜��C9�D���2�MZ�{?�~7��/�!�0�*9�'����0Bu޼�X�������]�(����&,�.�R�=�R���f�N2���.,�����Fj���J�v3���V[{��ڞj�V�&�7�J���Y"
�!�$���;�Y�s>�?���̼�^��y������ u�'!C�����!9h�{��P�-r�	��4Q˧��,菜5�	Y������9Ѯ�e7H��$ʺ��!b��^����p4�S��S܋H%�1�l�+z
�:�XX~%b���#�x��s9$��N��R�G��/�8��\��+\Вc�#hL�y�9��b��na�? ���M�g5��Ф՜J;p��x�w�+����B��X���z�-n�/"5��N��팿��x<%����E���M�W)�O.��d������?�{'���]*�
������x�4�y�Y���4E��Z��Y�Z6����Y�q���v	�F�������6$?�:�ظ�
�[�+�U^�A��:}��M-X|m�R ;?n7�FW�Z#b�<1��I)�W}ꬆE��޳�&'y�+S�:�X��t5��&�ҷ��e�L���� �������K^?)m���S��W��B7�mV��\�?���u*������~�P`��r�j1�mZ��ѤѨg+ހY)ի���P
(�Kh��du��Tu���MD���7�e�4��hs���&�^H��b@����z�Pz���>��ޝ�ә�o���u���ݢ~,�����c�%6���ةU����_���Q��z��������%7ϼA��܋'4�Il�^�h�6�A��{��<�o>n�~5oZ�5fEPb���{��4��s%.��E�J��W.� ?�3Z�_q�qĎ�	ސ芍t����{��Z��x���|d���)��[Nb18&?r�����I�����5����U�jR5^���J"�T��FJgo~�RE?$�5��QI�8_?��9\9߼Z�G4�����r�;OfquwZ��1�l�O��g���E���Zyӵ����]Ӎ������J^W|{U�f�bN�W}{�����{��U�?*(����֡�`Hק�v��d{��,$�{�:�1sJP	��C��@�h�I-�"h"P��E����;"�]�k۴MZY$*�[ԉ���k.��փI۠n!�ø*���t/(�zOX�\�߃S��|`��?#1��W+H��4���+浒��u�Ҳ�S��f�\�G0OD���8Bf�u�E \nl��v���1�h����V���o���oH"=]��	�^��F��|"ɽr�4�H�L��b_���v�W~U-�Bn�5�?N�_��>;��8�e��3|�+s�΀މ�~%�գ�����d�1<ny�Zb-y�2��ޣ{�_�W#�I�8��Bk���u�XA�fG���A�:b�B�5(�6������i�_��pVw� ����~��v�yє^΅��[j=�������ɟz�e��**�>�#F͓˹�rE������N����l4_8|�="~Ն�ɗ��@�(��?D"fUڜ�Bi����+=N3�����x�(k]���E�����%�Dw���П�;��D(�J�u�.���hw��f�
t�R��?x��԰��)�榈�E]
�/9��[�N���¸��LHWl��
��<��(�ީ�KyG��}�9J�S��9�;����Q�}�~��s��3�))v>=-�c�p�4Mx;��O�~�� `v֜�YU��+̀�r�%��Ҫ�W��z��ˢه�{�S�KKvgDGJ�*N�׾"�HU�$�����������f���ʉ�	WGX����.D��9��y�y�|�sM^���Gg %,@}����*fPRP1 �a��x�ax|����R�yo�����c��1;��t�2��K�d���.d���1�S�&�]΀`��#�6љ`Xp�����Nw�s�~ȹ���fveS~��e��[3H��HM�IZ�l���C��E$o�@�;(u6����6&"��%j"�Ꮩ�M��L>uN_�<H7vy��X�m��x�9��lRe�N�|��
a�u�>��T�I�zÖo���t��Z>�x?����<��1;~����0U��7�ޣ{�Nw5��L�����}��3�f2HI���UgǗu��ﳁ3��v�୩O��3��T��A������}�9Vp�l/��a5���#'�>fAX��!LM&é�I�`�ov/�B�ZT�޴?<(X8-�%}����sK�hͺcl��~����-u��K;�Ite��7>���[�ڮ�N��jCRM�%�����x�tB�i���:.���0�ڡ��!;���x���s����R�9�w��o�ۡX�ۋP��9�,��[\���y%�ECJ��-�j�C^o���{BDO�N���j�gI��|�b������tM�����G�^N|jC�#h�:4hgI�^�-x9��Y��I��SޤUד�XD��j"�s�f��sʿ-/*$�i��I�����?N�w�&7����4h]V�)r����Y�X���e7B��(Q�)d.(pw���'Z�os�}�E��
Z�ܼ�\�w�=�we����y���M�PβTİ~(��A�F�96 �(��9�Ԫ;�V����#�>��7�p��o���F�x�9+��TI[wR�-h����{~���c����=#��%e�<��o�`�hè��bH�#1�{�r�����������RJZ�fh�K����yh�F#f�`�:ߥ�c�Wmz���}��0�5�������E��q�9�ة�/�} �hi���K:�tDƋ�e/S���������쐥��u*�I�]\t���r��%���1T�@=��ȥ�X��D��+ï���%���5��#ٶ]���cl�b\Sҏ�!B Q����15?�?����d�$������i�3���.��9P:q����ʉu�%��/�.��E�ƌ���V��U��@4%�Q�svb�!,�	KЀqSq�K>��YU9��RE��j$�4��u�y��3�F���PQW(��d�_��8����s��-Jaj~&g��������V�ٰ�w�@��~/�ԏ��0"���]|��S�t��A�U�H��e�N�C�g�d�Er�i�B�ЀH�Y�9ĠM�r@�#�H�f����[�坊�-9�B#�;��ĕK�3�[D�x����[4V�ԣ�,�лsb4�G07�J��.�;�.�ǀ ���cE� o�&|/�"t����o��u�t�!w)�Wb�p�t�# �&.���4�gn�&�ȭOq�#>cN����	��w�n:_ �Z��fI=: �!�}'L'�逐��]v`��O&��)'��n�����HL�c�m�	&�>�����3�X�>I��|R��YÍ�#����ߧ�ZP��R�����[=����Wu�H��rw�Ms����J6`���1��}N�?Z�hAK���E�E�g�O�'�}#~Y��KA�Λ��U�_��oL�$���ޫʥU!��R��l���������K��� Z�=��"'�T��)bP�Aΐؠv�G,��q���gE�&���dQ��-���b��@O9��a�
k��b7%��y6в%���D=�����k�+��I'}1SŨ�d�q��i�2�T|��S�
��rwTb�6��y�!�-�����EWG�y�~Ô���'6��l�ƍb*�|Vi砀u� ���H�z���;G�u��9���tP<נc���Dɰ&��JʫL��wP��A���N�7�=%=a�#]����\H�v+�`�5��BFm�r�c���7=�,�.s >8Lީݫ�c=Q���=�%E���o�����'绐zp��0�f<���c��$'J�ت\�0��q��R��%����h��9�˚�:m�Q�l�o�?�WG����� ��T]���H>�G^�����kb�9v6��Fei�n�J��j\Fzor���Ƀ��C�<崳s�ӎ�A���b[�za������T�BV(�Ou�ɦ�	V��Bz��D��g����.X@*GeĘ�1�&�Yn�6�K�k���by}���z��ԅ����<(�U����D$&��m���y]��l��a�B�\A�!� y�:c�-�б������Ȥ�Q5ǘ6%�y9��U�(��"�H]2���M�?ѳ��v��5�$�����WGD:\��ɯ�����[Z��<�O�t��:e�а_��k��(�S�%���Yw�"s��Yxo-G�ߵW�/;�Z ����c~ߟN�E�mu��s�Uӫ���V!6��N����[�A�ַC�F��!���^��K��bN�
���V-gVD3Cy9��5�NX?����y�^!L��<�*�Kv���q.Gs\�T;pzy������)����t�̖�������M
ÙХG���%�C"Q(��oo�wx����P�dOl������lw�@��ðǬ�s�ԯ�������s~Q�yk��N������l����$�;q�\���jgZ�%�M�W[�����~V�����B�8C#�>�7F�Q�Tc���	��t8�Fv�F<�F��>�0+�S/"��C5.B�j��)�U4.�\��p�`�T��um���u|����\@�dF��F���˫�7͒���I�W̙��}�߅�
~ن�_�Euwr�FU^�X!r�J����������r��ܼ�js�Ҁ�|�"7�Q�>&e�̀�y=
�N%�J[�t2ge���e��"��غnʠ�ژN�pH##����;H�f���F���jɎz�*�J �>��^�]��EW@��}ʩ�-镠W�Q����h� *�Mˋ$��S���ǫ
� ��#7�!.%Z�ܱ��4�y9�%��+�R��d���o��6�=���!*��������h��uٖ�Vc.�����3%/CRԿh��*M�&��El�W�Ą� �>��Ժ&h���4���m�R9	�����cX�FRy������@�sU��7��Z3r?���:�%_۝���Yj� ��s��$��P�ʉ�4J�0S�
c7����6���E�n����R�cG�h�[��C\	wy��z�"ɛ� B.���/d_�h��3��us��B4#1�-�����9�r�ՒVR�}m�F+��al'��Z!�����v��]����r�h�S�L1N%�}c�z+C��V��B"U��ϢAW(��y�Ӷ�S�u�CN��Ќ�6?�WD
�f�d�nI���i��`��"ZO�S��&�h\F�+���� $Rޠ2��zJ��DR�v/��LĖ2|[�z^lN�/��M��
��i�Љ��Χg5(=5x��*�ǞFZF�
U��i�+j&�w?/b]����W��'2�n�}��
]T	�<̿;�S�-:
���,	��փp&\)ig��w��e�9�o3�P���nZ��\�;�(yU�KO<�nr�<լ� �߶/G����UB������c��#�fK��d��,�i�\��n���������p:�{U7���h�`�e{��B�;wӝ��_�bi��۰;N���SӾvl��ЙA���:bP�ք+@�X�}�Z]��i4G����֡vb��'r⇨gB	�����
#��S4�16���W�r4]X�����h��e�-((�#�����!�tW�֌t�����
����J��AB���A�A�
���I}"n�
�iB�9Sg�l������"$J{σ��Pq��?�%��Dj��yS`t@����ڃR_�����ut����;�����|@��Z�*!3�&q4��������դ�i�G
�J���}�whG_�jz�h�Ysn��yE���n��}=�׊y0����$xΧ�}�Q0�Mb�/�/�+���������O��D2����n{���C`��!��	"a���l�*��4GͰR{a!�W�Bq/L޷����ާ S�"گS�,4���������P��s�2�qr��s��ft�ԸB"m�K9sz�����ؗy}�$��]zj��ɪ͉�!�s*���F}�¡�۱j����N�.f�rb�r���F��%�?Ǆ���rD`J�no}��n���#�EoE*�^�E�n�{ǃC���p�m�hu�'��GE�	"I�$��L����n\��_�K__�K�IE�Y|Yf���i�'n��DTWm���]As��ha� ���%T��Jn�
�b���,�cod��g��g��S�P���t�%��w�ǔԈ���������ÒاM,Xn�{e�����E3���߁��!&;�'G����xx���9��Յ��"���
��Bs�ǍU��ŝ�=�ަ�����}M��=9��ҞY�I��>����J[D���%f�TR;�|�Dp�I�����rW�&��0�����:�n��"I*����&� KcH]қN�<Lڧ�N� )��qv�oH�~��~��ϖe��1Ύ��νs:�8' �c>Y/��qwi��aD��b�����R�1��Z�k��+��>Yu�O��A�n��:���U�q�1�qi�bސ�ߵ���x�� ��.' o����Z+�X��y@?b}/s7G���|b���yX�ZP4N�}�y�]������F~�hDj2ߺmX��R qP��IN ��n}݅��z�7��-
n���C��7T4O^?�EǍ6���:/TGǉӛx7m��!@PU�q�(������������Ei����dS��\�iRQ��S���>B�ʅ�~Tv��sXoӕ�&υ���s����+�\��p2�;�b�Pn*Ƙ;33�gu~u�N��i��bf'�[���J�t��u��iouߓ5�+�rV��f� E?�{]^wà@>:y^Sq䧖���>�8C�)�w�29��."���sZ@�
<d�޲VR�Vz��~�ل������,�.�wH^�7pbW�*9�9cȾ���u^X�'J��H�K���[������5	̱�W6Q�+N�)������!;gr ���jrs��� S���4���¥�a��:���%5scQ1�Q��:�j}��	R;K\���@�iGY�QW��=*�6�kL��}�*8�Y���A�[��&��'DRE����E�E�v�Ŧ̼���-L���k�:�]F�}�6bbc�>��Hn|��!�3ޯp�<!X$�A^t,}�TϋȆ;c�8^���/�fۛYh}�>�~��FZD�R���O�t\,/��ۨ[!}.Ձ��?|.�sޤ�Ls��A��,�[QqQ?QW��?��UT��<l�OD�u��X#�t):E��]B�]�i
�<�tP��h��6Gg����^�9�6O0�y�X��x�f>-��,v�V��q��\��.��oT���5![��nD?v���jum��-B!3&�+�j���;���J�J�8�ͨ��5��t�8�=��^O��d~��+<*��H��c��a�J$2�O�����
�~@�Ĥ�s�`Qz�|7 @488푡ȇK-��jnZ_�2�\䙠c�9	B���i�h�;�lWɮP�Uٸe��Qo�m��.�?�V�L_vp�q�g<��+Ts�e$_�� oZT�YV+T2��s�dEڪ�>^ySȖ���|Z�V�d�pf�"�zn�A�����GXT�sI���{DY�o0-�����W=�rE��9G�H�W��W�����'P�K�wg��o�rPҡ��*���ܰ��σÄ�T�|MD͇�c1�#%h�yR���0�N�e��uˇ����x���G0�Q�蟄�կ����)Bյ�v���8������aU�A"6�F��[�ֆݪ9	��JI+c���6 ѧVKB@$h��D�V�+��8"HC��>��bV@��o��
�z���&�����&� ��0�4�g�M�3��c�mW���{�/��@Y�RߟVM͓�'��aV��̓#E�U��Ҟv/Qs�<��7nW��r�������|��� c���½���T�Q��K|����*}��
�L��r�:�u��Qr�ON,��Ψ�u���iǙ��(��dq������E�X��)�{\��I~���*�D"������RX.w����R�椷M5ƞ��4�+z���M�#�_�/+�o���f#��Ǽ�i���f�����$���z�M���,!I�ReS�w2#�<��	�6�8��ʺ��>��#ǅ.�`�з!����o�S_V���G4�;ۀ+j�e	��o�����l:���S5Ė��f��ek(2eDh�61;�ҫ�QY��f�W��B�?tZ�M/��®�ֱ����,}��U�>��Ψ�G��� ���f�̜r��cN�V������ z��Q��u���kR?��iq���Ř1�r��7U��WK�����BI�nޭ�uI�e�Ҷl�)�*�/���(�%��V<fق�+���hɉG$��P�{l��	�r}�+/��:��	�����ñӵ��Eo/�X�̱�}[o_>�lc4ۄ�v��\�1�J!��-$���"��8u<]_Q=�"H��v�Br��4s^w�_���rKR�{� 8�T���y�_�
i��bVH;��h��<a��Z�[R#�CI�x)�(!I	���3����cڧ�t��#�9�g�wvқ�1�^I^9Iѽ�:�#~h�"�ʒ�uܘ���$D]���-��/'����}��zHuvw����Ok"�?��Ab��>:>���鵲�8k7�+m��S��d¥���e�J�_R�c�m4h���U����o��\:���6��<��اZ�!շö�w&���ޢ��(�5S�����_�3����Ne��{PV����` �$��C�{��L�>��q��La�+��'F,ߍ�~F�g��T����9ߔ2�N�:�>f@֐�a�ʱ�s�|�L��?��B|A[n��FR���/dK%����FyF'���Y������9J��:=�0���geℳ���8f ��!c���Ǖ�4?��$�7�0�7���I�Ʃ�����;�9���ZA���g���ld�۷n#+7�4�J�`�@|s�V��o�oZ���c�KG��Jˣ��_�Blv��tPխ�(����W�*���ډ�w�)͚S8i��Tɑ_�=��\ˬɘ�0æ�e�U����G�Sqj�j�k�b�4+�dC|�C��D�E����{E�k����'EGښ��Z���Nt�}��J��k� ��zPdK�Q�_ �_�U�c��Z�m|Xj�����|�J!])�	���68<gI���E��Y��������L�<�8���^�/ҽ���wT�J���6�}\*f2v
���o�l�/gV�!<m�'I/
���c��N7���\x<��w�*I����J��3k9o�T���e]a}MY�O"�)�}���?�l��{B�ǖ�;�,���䷂��W����)��tu�����h&�k �C�Ӄ�?��8�c��?�q��w���*����A�@'~���3
T�a9Y��2�u�����G�
��A���i�AN�L5ZB��$������غ�t�J�@����Eh�J�:_��=���L;�pS�'�_D�0m�q~Q��z�2�N��ڇ�_gl������"���*DR(�fdxw���͗��t.H�s���;L�r�wC�"T�EO���\U�Nbw�~D�4ț�)�_���F�w�3#�?����or�5$e��P'�Z��ԸAa�7�s���Ҩ�e��y�?;�'������d8�T)��Fs����lN���+��i�ٍ���ED��"�fe�o�(9��A�l�D��r�v_�U�*��WT��*�P���?7��#�>P�X�z�+;��Z�/y�>}�4��+'�<B.�S=��B99*�-�d>qBkVm	�+?\�uI�,�;Ɔ,��h�7!a\�7��ڡ����9��P#�4X�;��*��V�0���+MS��"mg�
x�`�ݟ��lx�-<H��/ 	��Ukv�y���c��t�f��CA#B/�T;J�U���e�Ւ}J��(G��~�k��_e��̈��Uu�hd:I���g�£ĵ+j3�H�8����s`(d*�S�Z#��	.�[ʳ��шԝ�wLi:�};��P1��o��-���k�� ��3[�-:��B;�����[mcL9y�����{|���T��V��^�Bb�5�Ea�I�l�̽��1Ү$BmOY+�|au�I�ДN��r���DB����!�IP�韑|�~���B�'���}�Y5�{HK_+%��tˉap
IGi�^g�j�/�l�[.�f/��$�]S ozWN,b�,Z�\^�U�c��ݐ8����8�Vc-x�Y�r��V�b����؀��w��[�@2�K8"]����r�m<5�߂��D<��}n������m��:]Cj�m�������Xh%p��%��YZ�}�޵\N^���6>2�8PiTm=�ǕJ�D;3[!Ϩ1=��ѓ�	DO�i[b�xE��/�B�I���uԌq�C�[G�����G�I��_������C����j�I� �����4�%Ӂ���6">/a}|I��w�ڈ����n=�N��<�rb�sGGkf ���B9�#���|�4�	ǿ��V�?�3�SC�9 ���n�Wսm�@
oM�����G[h�?4�oٱ�s̱gªgh�C@-��L��U�E1����kȉ��]��m �o���������1zS�K���$�Y@�J�Lj�@�}���s��|�5��3k���]�q�)��aT���S8\1u=�k���ݕ���sR|c�����*�6~�%�Q��e�M�D3��Wײ�.o�1'$'W��x��[`�=U8�N�*ԍK��Q��n�'i^�L-���Dl���ܛ��-7����S������y`� �n����	IG��o8-�x�籿@��S} ր��<��1���i@��1 �Y#A2N4#\U��P�M�Su�8���3exG}�²z��[�Ƀ���5�fK��#���j��J���� ��4##�^�D2/������fu��c���"�HAX��F�T�E���n:���t���:�̎�\�~�Y�����S�{Q*�Xǃn�Uku�ʺ�|��xx0���nѫ�d[���H��i���B���P~4�VhC��=V�cC7�$�|9�~��9�,h��=�d���P<�79���<� �����3��WK�a��/O%�q����l�n5:_����K�]B-%� s ]���t���ࢥ�K�����v(�%"���D�vYOY��,���l{�p���+�I�
���� �R���֟w-1��Zε�xb�c�r�=%��i�+!���\�ߵ�_s�D����ڷ"}Jc8�<r�Ƶ(߆��P�Z���V��N�G�<E���p�e:p��v&P:+1���ܼ��;���!����(^�������	
*�f�&6��mf$Xס�L��k#)E����D�����糱=��$�[?��1�E��Y���SC�J$iVy�tTљ��9/O��˪1�ȩA�P�� i1�۰%b�#�&��ˉ���kƵ^���o�4�פW���e�����˾�z�6�,�Ö� �ι[O�T�)�p��E�
�o� �|�H��X�ݯ<�oφ�d�U���m�9���τ2	M�8�+�X��U G;� ��4��ڡ�������_�r�"�M˘�"ا],������x�L½��T8�֗���[N�������X���9�8߿�T����K�`��y`���/ ���D�&��@�ͥ�퍝�<4߿��>�Zd)= ^�4/��3�>������!$�9�\�;&%�2����%y���a�"Q��2 u�aFhf�����ݩ,��=eiff��d���:4��Z'k�����+��x	.��o	a���;4���>/l(���Y[�TuA|��>�^�� �
��[?�-'�<v͸9�/_Q=ϮLs�ϗ�����.�"S����cbow����)m������M+
�1'>�9/�;��Q���ˮ�=��7ޒ�?�G
��)4�%�=r�F�=�qu����j�]��/pgr/jͅKaT�2�9�EU-6�ن���`�۵��+��ǐ�K���#^y���e��4^�����^z��-"�Rq�uʓ�{����e�\ѳ�v�<.v�M�Й-s�hB`EL#�a�|�Q�;
E]/����?�Gϓ��dܸA��յ�Mr�mux;�`H�M��=*6�/�����sc���x�İ����hF%QEe~G�X�B�P2_f=k�lwsf6x/�������^63�%`�ZR9��YU�]׊tT��˃���i��Lv����˚M'Tx�o�M�9�
xvp�� m��AO�T_C��a����Q�?��ݱO��;IX|�+�I>��*��`���($<����������F+�2��X�lQ���>����qk���e{1�p;�"�G��������^ �G�E��rYV��z�j�:�O�7i�S��V^��|h���907"C&w��-D��С�#�}G�u	���8�$���C��V��9��\�- ���FU1ו3��`_���Ni�PZ�f~lpDT�C4�!�#��� &�2�,�C��]t��pug����(��~L?b)�E�f�2A����Ց��Ȍj:�H"�^_<��/��u����z����xMDR�Us1�Mg�����Α��;0�_���A!�L'^Ϲ)�8���\k�\�|���Aj�H�aSݏV孡�Q�w�O`��`�	!Ao����gC����R�|6+q%���G�mE$�sC��z��g����*�BGM��<�#Tߥ_S�-q
LEq�M��'w���3�X���E���2�ݶhȫTڗϳ�<#�Nt{|��\^�� :oja6~��W}K5��D5��S0����G�����x)*栰��%�>*�5Wh\d��:l۱����S���=�}�@��׸*�� Jq��J�+�$�<z&�p�w�{Ϧk��T���i����z�� 	Q!_+V�v�*�:�_O�� � �;��!�Y��ʉ�������E��v��%Q���z���f��f �#S�g|��-|4�-�z.l
���H�*W�QSN�6\����*�]�Μz6���A�͜����S��ݤ��p^i��6������'�9��+66����b����pVevb|���G�`YPS���Uo�n鷍Fߤ�Yg)kX����Yv��bԛ+'`j�.C��ʑ���7�b;D�����4.�@E�މ��
׊���3�<х�1�q�=�?ɉ?�5"�U��d_2V���k����4$>���☇����ێ�l�11)�|�-���A�ZҨ�m�f&t�!X#WA�?�!]�o��Cl����7��Nfٗ��w�F����a`6�X��X�@�$�-�s�"AU��R��1x�V����o�;qmE�&7���� ���p����gJ��������}��-�L�\���`7�k�ǒH �n�rd�2�Z�ێ;D�A	��hL�ơ���S��f؃�D�G��M��2�F����e�j�I���o1cYOA�0�^��3;�U��RT.�{�!�+1�����"�=�P�r��Ho�N�K��{��QqG�+���Ʈ�*��c�ĊiE��C��� ��؝�X�F<�N�/*:��u�mB(Ո�y��?�6+���YL�a�Ҽ��jQ�n)T��IBo�h/Sh�C$���զ���J��X�{��ю��a�3��8�CG�xɊPR@�U�w��բt��0��~����AO6��;8��&�B�nI��0(��������Z����Є~[8	O+P�FQ�6��U�M@+c�����O#N vy��\���!�ƒI�d:�׸d�{�x�wO�U��FqCYW&v�k�Ҵ��U�aZ��~�Z��W�DN�4�:�{��uJY��w\j�d������70e����Y�-�2/�cv�A,f<�����a�_��7�)��ݲ���xڷ�qװ`
�ȵ�R�����.���0�����4�2ˊ}DZ#02�"@�5(�	Q%&t�0�tB���.&�S�L�=?(Y�~f�6����{�x�'�������]�)���ŏ��3�/����O0�S��N��Q(D��	�kQ�W=2���<o��:3cϲ�a�E�}WZl���N*���~�}�]"��'P����k��қ(�n����CH��Vl���� ��@3�����q���1tڔ*t@F�s�ʕ,\N�jR��C��B���Q�6:Ri\R�H�1f����((���f�P�y���m�Ռ}w76�e4�V�4n5�$�!`܆��PTV|o	�*'^�M���g'6�nh� d�i8UN�+��@��uf�Uހ~��Բb�?�@���!��7��M���cK"�͏~"��k�j�(�������5�@���CfD*k�����Pia��#0��/`���_d�e�:�7a��T�t��� =�o"�8m�o ����ݷ�z9$2E�\�1��U뭼*��*О�ו���q����&�w��%6�Ե�X�385"5}�_��,��"���1'X��1������j��W��6Nwh#�������^*�o֓w���
���L�{͹U�[�-��,/���C�Z���$A� r 18$���P����Vh��[1X܄�9tv}�1�-��K�R����������wl�8GZ��u>А�i�5�A���<g$�k�OO?$�[i��C�$�<$�Gev�U#7��q��PQ��m���J��>�̱��H@WAlZ)͓r�0љo����I��q�D�vxy�!�4yͧ�럆�yE��Bb,�D/e���izx���Nq���?���~|-���4��.q������y����!Mq�Ko.�rF�a���v�35�I�*]����?�5�)T���S��
�����Ӎ���c@���E!E~|������}h@���Jc�X�|��%)V&:Z,:��z&�d+_5�F8��i�{�yC�a�R�|_�WK�5.Ѹ�k��P�fi��������ENM�k�۩��a��f���'D��r���D�B��-��ԽܝiސY��Y5��5a/o�T��F*IX��]�:s���h�ZV��b�bk���kl5̛�v�.�-'b��ӿ�t$Ѫ���qA��0��4�s�B��A�c�� 		;d�����`�gM��9���qQ��A�S���>Ќ+�$
=��_���؆�<�N�H�&'a�s\�qD�{� 3#:��e�|��6�0$���iki�/�w�N��*<.�W��T�F�����0��9G�����oB{��Gq�����j�w��nną��x�	X5fN� !/�����3'$vǔL�n[^z{��"�yW�o� ֫&��'�s����sb�=Փ�ѧ�?���Ǜ3�w��XsFZ�£��i���b��+��7�|�V����AD3�����EAZё�ecsb���g��w����3�|jډ�����HT�F5�uN��I$z����رi�W�q��Rj��!��1&F-1�5p!��G#�P8Cg��!^�,����B�s��ҽ�-|���v��pTS��`,	�rc#wFX���p~�s�>�5c߳ˑ�ݘmP���l�zhi��U�����m��NB�e������Ά���-ӟ��������h��i�H�r
p8i� U�8{�*����Y�O ����A-���SO��AկX�)��9qF���D��7�����0���(8����/���I;r�(�9�HA+�	�&��*�����8�)q�V|��=���ÉA�@�����۾ps��hZ���_#�G��c��|���*^q��T;�P�?�^�TjJѹ�K$ZJS�P짝	m��=�;@�5�-�p������3��+y�ٞ�r�@z�KYm���t�H�A0_�c�8��xj¢���:Id]PD��z*�������/c�k�9M�S��
��9tv}�d4AH��c4����mq95�^t����?�����kY�5���<�J� X=}faHW��	�U��ťG任"l�^.�f-�D �2���5Gy!I���U���@���}�������kZ\��̅�v:mn���A�`�x�� kE,�:���9�Im�ަ�F|f�i��Eb�����qI�*�=�%� 7ᐟ�ak�Y��6Z�P44a/Է�ҋ���ҩk{�j���f�������6���s�<Z�lw�U��}��>>/�a@V|8h[47�`��e�'��lo꥾ocu9�o�ĺ�|ȉأ=��#X�L눐NָE��|�=�OZ��5�r��˗v�q��0��ˡ�������7�z��9ٝ�����X���x��O�:�8ۙ����4�^p�̃� �e����>�`��������:v@��*����EY��9����%o���$+d��$�H�Q|m+Ac�7T�/lD�+�M�ꦚs����c�/}G�8���n$�̕�n?����ۡ�؇a_wH�=7���;�Ȓ7Sr&�e��{b�+�AB����Ȥ��$W+�/��V,'�v�d�D��<yͅvf�żFD���~�&�1dN-�JX�-nv���3*)�R��x�^��!#fgh�N��:���cQ��!��̧�Oޞe{U��ڡÑ*�ϐ��ED�J:��촱�~��:qY���O~o�:�^ЁbD��3v8}ktxro��c�����dO�3��7h�������o��Tr/��g�.j��ַ��WCv���u��a͉x��K�������*E���*` 5�� ��~?�uWY4_�X�x�[���n�I�CU5�.�"o�����K������e��i��$�q���ٵ�~��q�l�����r�b5e~W�.�����D��}�͙��v��!��K1��L��0R��p`���O��I3�`��YW��f� �Ÿ�$����y�h'��/��R��aj1�F��y�d:��E����A>��'sp;>��n��pMF�?�$�Z#�U~WGU�+u-Ǔ-�6�����D-@�䎭�=�����Z�R9=�:9bW���c��Krb<'�\��9�U�xv91��N��;��/r��t��Ր��PAL��?���w��n<�Z�n�E���{��~�j~Y�����rt%f�u@a`�H	�;�Kmh��o�Q��0�S�N� ���s�f�N}4�)2�9P�Y$w㦫���N+���I7�_�ug�J��vˮp�<UWHBa��P=.G�RJ�S��#:��m��r�/���6W�r���)�iI���Esi%Qu8P��_V蒛����u�#���z��@�Q�N�GRH#��42�I��bf�Î%�b^֧�ؽd���w�ݗ�}Aw
���f�aՈoa�𺬙ࣝ�	��A��r�(� 'f2����8\�}\�P�KI����+1����'k֗f��1^?Ac�2��/ �j^��WI�ǭ{��=�פ~Q�����l����*;>
���9q�;���$}��l�	�	�n�����!��+r��0���x)��e�C����ܧ�PL��G�����0�� �h~\H�n�����vH��	 Ԙ�����&e�˰n� ����:ZܟQ|^�%��>��$���N?�^�m�LWE]���v1�N91�+���+=��1�0O��t�)������^�r�;(&]N���� rb�H���?����Il�)C���s��њ��u��iؑx���^�^.K���՘l�O�A��9�m���=�v91s��04��s���B��5���J:�=Z]h�iM��+�@ג�P�\��*#A�.�O�%�2�&���QLu�����A-�����ig�% ?����S�|#p�ߵ�e�l|x��/u��oӈ��n��K���ps��/o�c��^�x�Ź�0���u�/��MR/Z���"�9��{��.���x��m�%���blmf��_��GDG������X���tT��?�<�ϩ$�/(Rm�=����k�3��j�xխ����0'�!QHn�0��.�$��{�A@�ŶBC����.�J��=JO+q:k�8��dZ|�����	gWt���$�ᙳ���heԃa=B�kS:�,;�_����/q��9�����D��p@{�_�5������epy'� Ѭ�ҹRM�������7��D��#�G%"��r�Ҵt��teAl,��(̰�F�K��⮧f �lp;���i�Egf�K��^<	��Q9ܭ�r�<�(5�&� 	��3D��|�h�Dʲ��E����oCo��#��`���+L	��H��t"�< h�Fol�8��V��TS��w�c��JD��",�kpe��mF�ѐ�����Wwְ9�qi�+�W��g\ �-�`iKDu�|��H���)]��Q�s%�,3�N���E<p?�vq3n��@��Unފ�u��9ǖ����AC�הZ���������Tn�[���5�q婶��d��=�_��5��9��G�h7\�������U �8�Vё������D��p�]�5�nר|aV�wA?W�)���9�ކS����
@�����p!���>��r�u<�lqլ��%^�S��K�N��c�˛�Q}*I~�q(�\:v`u�χ(��(�˽�fі��3u#'�+��aag���v��J�}]�̟�\�y��}��5�=��kA�
HI�o��$b|�n��
YN��l��O��vi:�L5�����n���E�$k���)��i�Z��'�V^OI!#PH�BX�>�j�ԙ��p�+v+B�4��ا,��K���gIN��ϱ0�j7r}&Z��_�R�6����+"ī��%�F��zy�g�_N,bE��C�$�D�}�}��V�y���Y-�>�j�K�S�;�V1�+�M�5<Y�'�����t�/,LUf�7���w1a���r��� ���w�vzf�n�e��ӏߣ�x�
T:O����oP�ϩc�Y�O����dֺ�\�<7\��;��H�y�r��{�m�r�q����l��숐o�WN�_]�Zc�5(q�`�7�V���������1}\�`���U~
$7��w��FN,c3�/�ϩ[�-�w��x�c�+︾]\q�?�+��Qv�!���m�?�l�"��Qs�9jZ���z�]G�*�3l���.��sg�`�wy3g�^k��ѭ�si1�C�`�����&+Z*!<�D�g�RF�]�-�"`���D*�,��rb�4$@�MN;��9mrQK��
}t<-�&�Z~|�W3���܆
���������0�c��#�밡�4����!�Zl�'%���e�~1P��8G�b��^d̦�oh����%�3��^~	Ƣ��`�*���Nq��3(N2���L�!�����α�� �PELK�}/��f�ޅZ���?�+�j���b�V��I���r�(�6���z���e��Q���I]�ko��y�K8�c,� D�����C_���ky��gG�6��C�����~3 	�$�	v����|%<��
��֓����Nct�	%2Ko�.�ޒ�]�x��|���8u���7���Rޯ0��Ԥ���d4H��_N����������_+��Z֕�y��5������1=�؋8+r�} �ߡ{���N���.�:���l�a�hπ-ph`�"�qb$'���#KU|�Nwf����1��C$��<�H�;.��
9.�7laԤ���:{�+�/a����v���ju�D�ʕ�P�R���g^�����o��4�L����ȿ3�
�xC�+:��\b���s��D��Y�B/H�"v5���C슽��%�q��-@ӵbk������a��;�fJ|v�G��e�.;���I�N�0��s�zBjq��|T�X�VV�C.�m�k���U^�2�����w�z#;���I��s=gja�����cx����`��%��6.�H�}��$�_GM�]K�Ћ[+�:����P����kY�'�S��s4�T\I�\�+�.�^	1��� CY��9Lf�"2!6&���bv���T���V��b�[����>�%��T3��B��0H�&z(��QM�0Z2Ͽ�0�řK��
y�~,dx�5w�h�gee�<���b���԰�o��Q�&,���u�-;�Ʈ2�=ڬ�{`�:fu��	t���r�̭��m���k�7#OѷA{0gI���+�q�Ur]��#@�q�>�"Z�;4�f�ٍ͗��F�7�В�g�*�B��%p�'�/�U����Ñ U3�gj���b�m}�P�g��Ԍ���9m0�T�me{����{.d4�֛~�q՛FMq�u��e=e{Q?���S�=�u��'Fe� �u�2�c#D�"�1�"��wc�Y���W����O#�ܿM�7��b$]�X�DŰrU���<�O�����z�ͨ)4���ȉ�#�g�r	�>v9\%��ߐد�k߰mx��R�ܴ��+���z�xIl�fܘ��8�EP�4��|�V�����x�������jTϦ��1���:}׉p9�8u#����|K)�Ȉ���r�
PO����,>RO�%,&D��Jrr"���3ơ��8�D�*=5��"�$�x9�~�?#�pBc�o��{|�� V��ʛ����>�Fh��>z~dio��C����5X�M�tO��`���D�!�mW�{!JU��Y�Q|��<h���<�*e ]�C�-,]� <s�;���s���4���PȸA��+�p���-��Z�H���)�.;#���/0�/�_p�V��^��ROG)9�y����O#��^�	��ݵ>��j)�l��\��s�i���CE�� ,)�����Z�T	Jep��2ҕ����	�9 ��b��"���J;]v䆡LA��۶�;�5OWwzE��%%�ҥR�r���aR�g�%5��]^8����`%��D_N���N�Ń�)d�ԗ�_c�w����w �xX�
n�qX��E�B�r
��|[y5s��ٝzV�m�_)7tU�y��H�EL+u�P��I��\3.E�6���7C�֐��|�yؔ����^3e���C��cИ��J<r"��}������q8�=Ò�L@�JƪI��{O�M������o��_Y.��BAT�l��]c�_�B�1:D4H:��z��>+��"RS��U��Ӓfξr@3'o�/�}v����߃L�����?�֫=N���!q��֣��yM�^k�: 'G$,j-]�0��K��d�|;t�+����u]��S�D\H�
(^W�*�hu�#2����=�Sߪ�i��!��	 ���BU�H�d��uv{t�5���x\����<_����ʃN�9�zg��R�����8ϰ��"r9���%-d�4����c��c�m9�itvS{���!�1��"������Y��Y�����s�%��s]��>�H��㝪����B+=J��(ЅEO���}~��2*m�L�����3�*��7�ҁ�½9��s�����"H��ϭ�Kf���G���Z�]�[c�QMJy����"?~|u'ZG@�yMm�Ý~�;�!�h��)j58�jϧ!&0�/�c�g4}����6U��F�4d>
�ߚ9e W@[����zU������?�<|���o������-<�z���5Z}g�$Ό.�qu��Ƣ�r͌���j���wx��wB�:�2� ��x��ߘč�6ոr,��#�h�^����oq�^�s4��T�pƨR��f>��Ƣ�ըR��|�&:_ƖZ�I1�<<�C��ǵ�S�[:vՃ�}cH�dWl"��#��j�Q#7��\7rh-T��:��q�lRB�s�Uߓ��6�Z���B�GJ�j̉�һ�>k6�g�mzXh=�M_ )9)��?����ժS#'Y0�Y)�����;��XN��^��ڇ��AVؾaZ�~�V�+h^���r��Q�z���Jha��P<~���%�W����{C^[#	L)������2V�ر����e���J��.`�=�ie���BHC�j��?P+���<)E/���uuO��x�'P1�_N�b�m��-��J�t�"7��Q��pK���ˋ��($h%�� !�>�c&����S��?��:���S�+'���(OH��Bf5^{*�+�QTh���#����+HS��qV�I:4p������~���5�F�1��T�lLDd��f]�z��~c®;�H���C��G߾2�ְ��r9����k��O���D����e��Xf�R�� 	��n��}p��y���<�k�'P�"v��������A�=J�����}9��J�`"=b�x����&bp=����7�wT]"I��.�y��/���4����)�֑]�|ȟ�e�=�k��F���8�I"�`w���-[�P���96�y��N�&j.p{��-H������NY�bh��_$�Z��<���!����#�����'\U4�i=�n998nY1���b9�8i�=��r@U=�jҖF�k�����L�+?��K�?��<����M�@deѨA�&�5�Tw��0B�T�`�^i�ET.�ݵL����֯ն��Zm���Z�H%	�������6CD	j d����{��nP���y~>�dwv��9�y�{��t�3M�y�����P�W!���!��S�^U�|9�!�;~0�ײl���3��̼�Dp���Jx�9���s{�.qF�ٌŽ��ΟS��S�WnN�g��� G�}�����PS�T��!g4Q�@�^U!�%0X��R�WY��`�G;2l$�0�0�y��������"�P��?@���VG�Wk�M�p�pb&�u�Ź�ߴ�����c�x��AT3D)�BZ������%����	�������W6��)]ḫ(B������v]?l�x�&p�}���Ђ:B����ZG�P���0�EL�7��D�HKT�0�P�}�"�J�A�^�t�Ǵs$՞@�/�=�^]��k���N�r���M�핌%�œ ���	��t�i�D��M�(zua�|U��q~��|�4���^�5u~}��Zy?J�����������p�
xr�G՘S��6���=�04(�FЩhw��z�)���z(>7�f���Ğ<w�1�ѩ,�
�e�1N�1��.�i8lFU��n�@��Հ����Xq�&��F�d_��;I3�O��� ����HH�zڼZV���K/-�݊���]��u���4|1���Jw����u��)�]�AdiV~J�-�5�^��q��!��.Z���(�?��(�K���-X!"2�������h_r����@��H_�Hc����d���e�؜���E��������i�Q�&��n�o!N����ͷ�'s�|��Ϭ��tZe�z�JI��\)��jG�ib��)�N@�|�����s��B���;��Fm����x*���׵���0z��m���v��v�(1���Q��+�-e�e��H��|��i��߹O�n��B'�����"�џW����rDQ6�`;�`� $6�'���S6����^@�o����Uc�@:$��:���t1o%�������p����=��}�
U���ͭ����'}���o�z��=G�괨 �p݉�^������Y�	$�#0e�ǩe�N�끩�Xw�gvP��f��᳔ �����mJ��i1�I��Td��X����/�~�_Vʱ�r=�*-���o���YOZ��ɔ�8�@�2�u+;�Ն9.������F�4��v�#��%����,{MZjN<�V���T_�e1:�w��Ƹ�����e2�Ϊyc9�H�78��C�#Ze��{
��q�1��t��`�Wx�"i�y�	���1�Moet�sV��ˉ�߂������>�F!��!_Ao�nZd�h�+-���Vr���9.���-��q�^�ptw��|�J�������_H��s]cO����#j W��a�`��/9O�n�0)����Uݴ��hґ�.8��v~���/D3��5�^ҟ�65�jF
��&�C��~����M��[���`߼�hj�s9��Ut��;�bi�,�fs���,$b�^}�p�z��x�}:�"tr���0�&q[Q�T����`��5�Ϻ<�U�Ӻ�k�O�sI*S��1�����Av���k#{��Y5FA�B�!jO��~	�a�II��kmm����K8�(T4���N�oG�IA������1����ls��&����I"[��]$�-$�ZH#��BP�^N��'Űr!�+?��V����7���/��d�5���4�.C�kzE��x�S���$���
�*�3�MƧ�'�mA�1f�^5����Fr�u� �p��8I��|��C{|cI79��`8�����,"��4mƚg���O貟�^"1�9aպ��;��p
s��nv�ĳ��?���u���ƹc�G>��SJ"�lh�ii(�O��ؘ1օj�]�5�uz?��da�Kál�!�O��F�eE�Fpz���h۷�kM�B3���[���9\����܍>f���uE�2o��#%�������TS�C�?y�����n��&��L$�/�<\���C��;$���k�҉�����>��4�u���S]������NDW3�^�h�I*(*��8��8e�6�7�^������D==�z0 ��"���0Ҏ{��GA�M��u��/��v����-<�Ü����.�Ϭ� a�T$$��X��DZ.��5{sN=��y���v{���=!�}U�B#�}��q5ʖ�������>w��b"���^u}yG�����@��Y��c �Vuo�>��v�'Î��֪	<qV�[ץ=��$'�=�*��Όm�v��3r�9\�-��T(���#�ܳ����
ِ��l�a]�B��C%L��ݑC#�Kk�Df����y�_�+�oJ��a�߮�����6���
������]J�}�}���#�� �4��`�u�Q�.�����.���V��W�j�.�=!)����Q�o,�G�g?4j��m5*rP��S��R��'�S8��y��p�&��L�8��/�z�"��dTn�!k
rlt���@�§�*��y�Xy ���h�� :�
���i���3e�JϨ���% /�K��F"DT(:��'.ʛbmna��K��4#'�LH�f)�M����\�ԣ����4cF����|��鞙�Ȉ�ʥ�������F}Q�/��}>fͣ��#ƉxߐR��/!�H�CH��?��F�nA�y]��/q��[P�q�j�}��"���Rs�j�9SE�����A�kDݴ`�"�y��/�@r����2
�<�M~Y����a�^�A��9��ɤ;r�>,$��
��q���2���������̋���I�����=7���ҹ�~��#�L�dd\�H�/ξ�/�72{���A0vt�AG���g�L0���ey
��3�'a�/+*�L�*Q{�g��0L�a��\|4��%݀��׋�a���-� ]�-౶*� �o�H�
{|�^%��H����[��8�g��&�A�Ԯ�$��1#T�6 
3]�R�Ǩ��U�d�6�J�,�|�:����+�,�����5Hsv��R��*�ж>��5 A<�J�D=i��C##1ı��7%V5����e]b@j�u9+��ү�>*^Ur^�����@ �g�,��*��5������yH;i�π��x��E4DO`�G��r���E���8Q�W�/Q��F'E�C�j����ڌ�Ԓ�Z��T6�41X���@�_���ۘ>���&Q�z�Q�� ia���U���+bW	����z/i�I,�;������g��@yrŷ`��j�a���d�c=�c���Q>$����;���!t#Ph۶���Ӛ¾l��y�N�ڴ|��oS\_��&���9�La���h�壉v�����:V�!٦�����[~[��V�)ee)�2�'��+�?��@ИS�C`�r��®��MrE�ڮVڦ����Z@& &�D��X���})��s���~�|����`�Y?�$��U�׺��T��#�#O!�ϭ�.��a�Ahl����������2&$>Gx�Cy����6�d���}5z2�wp���C�ArG`��xfr�Ax�����U�w>�:�h�B32�l�3p�];�Ruf-��z7[D�'A�G{�e'M����,��K��@����+���_�ۼ��y����¡�|#P�����N��#�2z����Ӯ"����T�*q���rH��)�?��w_�����7�Aڲ�oG���$^���"%v}7���:`�B%�;���uf-� J~
)�1vVR�1�(��稻���S�lxpA��?7c��muF�m�,%��54�4�YV�)�p���8�Dݏ�E躺�"�]������ܴYH:��p�8�C�K�TbcP>vW�h�%s��4H'�n:6�yT��Z�8� ��ًcΡ{�8�����X������l_?� �o� h��m_?���3}���ѳ	�$1X�r�������r��`���Кa��K\���)�C�47���
�*4���F�P���W��C���.m�j���N�_>�&&��ntP���~��F������K�
�F�7�p���Ӏ�C�4g�F
��Z\+	���r��Gs0�����:�O
�1�y�Ջ˕�$����q���1��,ߥ��}��m@�%k�AL8�h��tZ�F���B�nG�.�+8>!:����9��/#:�CU=������;ta��VK�O:�`:o֟џ�m�>P�q���q�Ő��C�c�@Yf��S���(A��r��S����PN7��/�Ig�@�@BK�!i���~QUi��)Q�����>�,�]X69V.��S��U��G�z�t� �s�;��q����<���	}�rp(}(Ƈb�P�&�P�e���A�hA��9�j�C>4Їy�0�>,ć��a�\,?Q{"��u��D���.�w��	m5��(�����4ޫ��t�!gg���!c�;�k�롿�}M-�����K��������[B��/q��>��q&�F���Z�K�����@��_R�f�L\���yQ��$>6=U���b���Ŭ�	�g��kB��X���:�>B4[BE���ev�7�:r���5�?�S�S�,����~v�d):4�J�Dِ��e3쵏8D�~$��+�
7����\�fx�~X#W����D���ƤƅKҘ(b�5���t�2�ZPo1��$"�	�E۝$�M�;f���f���j������2����ѹ��U�W �����eQ���3��>���!|P����\ii���L�GF5��*��r+��ɋ�a�;å���hXx8S�Ȑ=��M馀�����~<�&��
Yl���I�F�{�P�n��!�$���a|k z��:��O��g���㻄�_MNf����nT-�VBVT���Y����+Ug͸1���;�y2R6�q14��9.�Z����,��%����7���G�����G��ߑ�?�(λ�w�gj�[�-�M��+[\��7�0�D���d��Gջ�a6|�h��sPe~�<T��!�C�~�y�S��:���X��ҼC���P��_āX��z�����|��+��ߧ�a;Q�&,��I��$̣�,y��8�4@����d��I���)�����u������fxz�4�"��TQ�k6
����h����!��^N��g�_B��t,kIF�]&��>�S5���a�U���p�R=q�VSo����.����aV ��e��c�L�b.:�-+�\�kQ�½W����L�>G3�RM�6���Kgo+n!�l��v�GFi����S�3Y&�Q'�
�5S�����4����&W��s�����PyD��n����uiw=�0w�����L��^��}�%���/�`�в^���t:��i�R�N-=M3�a�,��a퟿ӯ�~ḽ���{˝K<y��V�+�
��v�?%���l����ɔ����=��>8����곩'��;��	tj/lA��x��D��߸�k
�S�-=����sK�� ��Y�u^�Z�+iʡ��E��M|=V!�
�eI����ʦ���V7��.;��[�2hy��S��b���!���Ee���PR��~4������x䗌��Mɓt��������VB��b�=���y�a�}*����,�ؖ^���`j�SY��= ���>�B�˝�FV�tO�}�^�#���̸����eH����.Bd�5U�8YP��-�K�_���PVl}�.�tS�m��� 7G�9��o�3�o�P�
���I\�JX%a��m��Z$���X��� �H����iP��/_!��K���A�*��^ ���b�9��2�F�����Utw�[=�)�M��Tt��>Ll�6��*�bc���T�G���V*��O�{�lf�}1qW���1��,B���!���U�aя��~qs�������W^��d?}D��s?���#��G0���9Z3�\u����
Mo%Ra.�K��B��	\ؽOӑ)C��~nU]��A����I=՗���7`+sZ������{I���^_���\�%���G!����֥���G�T�k)i�k�˽�5��k��MǑI�~Ӫ�h�t�@i�E�[�g/�Q���M{q�D�4�����*��q=-^�&�jy��?�?J|���T�0�����������z��#��M�Ih�m�E;�V(Q�8��o&\��4P��{�;���^�2�F9��Ú<S��	�wF��tzlW(�Vd�R��-����������8�a|φ�5;=G�UGߞ��8�m�ם�����*�+�[��</�A/j�Q�=d��W�2�&ީ�a[9�b�!���#�	�"�p�Ñ�T{n='<v o\n�[
'�_�-,m�\��ڴ��V�_�#c�r��w �4�٫�8?d'd}~P~ˋٽ�%V��[)���9�� �Ú��^s�����H[�������w+�i��\i{/�S9$P�	� UZ4�-?I�B}�]�w�@���5g]�(c��ʩ�����?�ς�~>Nv/����i�k��/�[�j�8e����?�Kk���=a��C�����&�����j���BNN5���&�cDKR�bV6�4V�&~�4"+�jN�Br��b�Ÿ��9�o%��@Ք�����u��[l˃b;���3��"��i�S���+D�c�)��2 �O�Ч�ފ|�X�7�bj4n@����WNp�x46�����=˅hq+�Ĩ��A\fl����:������╞��C},ҕ����:�E�9.lM�u8��1z���M�e&v=��_��[����������׊M�}�`hJD��T�v�9�'%2rc0�������w|�ZT�O�t�ENEBs�RA���h�;2���B�v�|W䠺�D>�#$�)�^cc$$7b=���_�_� ��֦~�#)M�g�v���&�ׂ��A�S4X�	]c��T�ɿ��56��"K0#��X6��5�bd��J2*�E�Gr�K���~��ǜ�/I�`V,$�7�I�����jth��<��3՞�9hp�Q5N��S���oLK� #�C��A��d�:�өi	9��]E�pu�+�f3�oY���/���vX�s��Oʏt QhȈ���mf�ި�L�c)�V3꽍ze% |6�*،���r�&T6�I��oTOj�V�͇�i֓o��,Λ�����^5��Q�ٶY���8�������!�vc_��g���?Z��M�T�+�H��������0��>N�FD���kN������o�5:e�e���	�Y��SҀB|/N1=͈�"���i4�z��: �i���>�jQؕ���v�:�RbJ��A(1�i�)j�x���kN@��b�'�|�w� �
�c~��p���1&׭�F�l.Ǒ�fsǫ�l�}���rG�[�y��$Z�y� "/�)��J�&1A�C��Az��.G�t>���	0I%r��t�u�[�� J�[[
��Jw��&�`��	%�}�0v=�2�D�΋�x	�63�Y�#D493�~�'�J�u���-�mm@�1�؞J�S�}��28�ny��ĥ��|��^uY�%<d���6�J�}�*�WO*�хp��n�^�R�cX����8�~�x�;S R��r�Pn�����nB2e��kW�S��lD?�<�I��x�Oo�8�!���Q�G����AS��jzu?Ha}g�X�	�N"dF�_Z����s�]����·M��N&,�5.و������@/��x���a"
M�)녍#�:�/���Y�8�m� �,�VM��n����(���U��t�@7J��N?�9���E�(�=��aB�]#�Ȼ�2#*�?�ٌBɼ�r�Y�l�nO�:C��_j8l��s$�K���d]�{�o�G���9�)}��L�Me;Jz�>,4�G���o<,� <L��xk�cq9|�*�O/Q���i���o��5 mb|����M"6h�;@R�������ě�'b\2����<�V BoPbi��m�"i����F�i�Q}�_fW�`!���^$�~9�n�Io��ϖ�u�D������%lTLA�[��dxhl�C|D�\�j����R��q�'h�R��G�g���\
91���ă�#�����6`p�'��&h�Jo��zu���� p�[��Ǝʳ��ȧ�p�0A��I�����W�'yл`��dI�G�~��\a�-��1�Vַ��	�F$qe
5]D^�<��`��&��Bz��>���f���k��a��KZ�su���J���<�$`�6'}+)�$���qt�3����(��i���_.������Iq�Mdw�Z��@!�4Ǎ�ٺ�������>��ޡ���H���t�
��E��^�p��~�fh�~z�=�|wt�����W>�.E(y֟�dB:��#:(�\"ţ`U��D�[����F bU�\K�ͺ��.� )�h�RtZd��ؼ~`��B3|��A/Z	�і\�'%�	ta�!5m���?���Krw����g�&M��Wq,rv� 斨u�,+c�s��:t�!�Uu��Ag���⯹OPG<�;X�˾�m�7A��O�lB(a~���ʹ~IEs��Bޙ��h�n����s�R�A�<���������,������oR�`%�O�'`©#.�! �#����3����o�����7W\L����,vf�!ur�ór0���9�9��9#ʦ�\Tʵ�m���7�>]����ʊ���9��ڋق׉�v*�HuQ:6P�7��g!M��F��B��]0ZE;��������y�H��qZ�g��v�����ESA�߫�伽$!��{/=�QB"�I�p/J'q�'���$��)�yB<(&OXAjqs����WOJ!5�?�K��Hҗ�U�N��h�F���K��%R�̱��n��+���{�x�<�5M���y������e��DR���´}1�o�,��#�u�,m�:D�%-Mh>		U�i"�-M$�Sқ�AS�#�Rls������@�0-ɇWTI�]��;Gh�}����vN�[
�V=M��-��dZ����0U41�#����S�O�&k�o�J�)Ԕ}Z���Np���M8r��n����0�ջ�2�=�X�_=p���j=���Y���������p�`\�W�{W�1�v4e{�p�/J�k����j�"W3@N�M��L���Dn�`Ns����l�2�d�I��ux��"��cf��dJ����4ö^����$�^���@>���n��[���^ϻ?�$z8�t�f���"�,C=H��}���.��c�=r��I����zK���+��oD��՝�e�	�A�_�
]���h�T}�I+����f����~c(���W۝���8&N{ﺁ��#a:���y�ɬ͔�=�^��Ud�S��z���/�7֖���l������ia
��ia꒞�w�Ti���="��I#+�-����	��:"�����Uo��: ����$Sv���#��e�.V�;A�v�D�(�)[$�����tC0�����a��{�g�}�_&@"M���������v*+���c��Pq���rd�20��~���4�4;&|eZ�b�2geM�{rZ;��ukzZ����#"��b�9��/%�V�/a^��+Rn'$DF�~������rp�h d��M5���5&�n�᫐�%f�ܾ�=^��4��hO.{4�v���ϾH�d��18�ꌷ��~e����U��1���Ꟗ�j�w���.��.B���+0.K%۝��6o����(�H��څ�ũrU��F��|�a�!�w�b�����I��u:�,,����lNt����/%���.ĺ����OLq�/�\�9�xxz,���*2/���"_�Ӓ%@��n�����c�\բ���dQ��\�$����Yӧ��cŭ�����*��I��1@4�ʮ4ێ&S����r����^Wz����[r4����⺣r�L�5�-A�,?�^����]���Dee~�3���"����}1VlTJ�c��"lb:B�̭=�L��o��o��I�Z����E.��K��#v�c�r��a���0�C�VT"�v'縻�7Dr�Yr�=��K	ig B��v�
	
�pe���B����-v��FoЌʒ��-����+���#���&�H1�g��:�ȉ.G���9���-w*�7�K��+m��Q��y��-���՞�j��-����#��c��ǅ��=�\�[�bF�ˣ��ʅ�i�B����%�h5�Zqi*�sř�]9(�kDV��g�+���XIB�*s�Cpը����t�S�	�>?�;��^���!�ـ�x�c��=]J��b9�4�I�gD�FZ�~�Щ�P!��w�+rH�X[רN��_~� �9"{��#:�����4%t�kG�`G��CLP~l��z��iU���X�3�CϘ�΢m�cf_ʺ���S�G��յ?�uf=�}�WZ&�`uz���2]�Y���%��Y�(�r	f��X̒� ��L�������&����)�֏EU��#_b�\J��<<�#��7�O�w�~�e)��`�Ŷ`h�yH|"�0�������<λ���Ҁ�=��|�'��CH�y��� .�Ġ��(O��[�g
��W6�_=��t<	��C�S>8�V�B�Ĩ��eV�2S���$
t���| �K}Eq�٧��ѩLj�W��A��/�#6F[	��l"��?×v�J�v1UAa@�ѽ>eC��_�rdl(�"3��Q̒�l�KxV�0�o�M+&9V�&��7�� bǾ���QL�Ǔg�h�u��T
m3�Se�IAW��{��`��2W9�5r4�=.���v��	��#�J7��+�]�[ـi^8)�l�T�����J���~J��4���,B��_�|w��!�w'D�B���3ߓ�4�pTpG	����j���ʱ
�8�ص/|��&�p�1����������4g%�޻)&����ʡ��)�q����H��{�a%�̗fG� ��)|�ۺ^�����T�w�8�K`��: ��1�t�#���.bê=Y1:� �Ď0r���c~}	j]��F�R�p|ktq2fԆP��6�3;c5��n-vAFO�_q~q�\*��n�5���<qm���Y���-��9��ܝ��	�xK{��ˋ3S�5��̣�5����-<A����ڰKӫ4}!��U����ML���ֺ���wk�>b�^z�M7��t�m�1�?Kd򣳨5��/6�q��/�Uwf��/�Jt=QL�|R|.�����jo�����]�D���,�(�1��F�I���=N�ܛ�Y�^��jn�Y��i$�9i�^b���;Z�z �1��m+�Ur�#���|�Qm՘V4�,V�Z���R��tr�_}����o#Ks�(�e/;\�S�,��0kI��S�]�?G��֠�A�7��6�e��`m�%	��b���1��ޚZ�9?ӌ��Z��m�pW_j�X�[�����d	޺m��X�t�AgxPi��w�	���CJ[�s�,ڜ����|��0}oB?�Җ?����E�mP������b�������Z]w�?h\U~��ɚ�%� 5+��
j�G/�;�ÿ"�5�o3?>���^H_PL��;�ZC�0�_��[y���ےiz�$h�%F7�~�o3W݆�4s}']~�V��O3���N{^��*���#���zi��������I���F'۱S�Bx��2pXҦ˚�Q%N�1���k8'�X�w�Ko�.+Z��%6�b������~W�y�{��}��3�>^SP����uf��.yG�~�A�R�l���lT����Ѯ�ѓ*�'5t�5��Z�������k��\&W:�y�(�ﰛ%������#�0�bʺ�-���u��s\�8+����L@
*��4�ǋ8�I#y�>|�*��q6��7���Ր Ԇ+��T%֠Ɯ���uى�<z�-0����z�>�\Rz��=�D��>�D_6��A��%JF�9��XP����Y(���)���&>�4�No����ta�W�.�t�]�WДs��ĺ�y��Ll�y$u��	Yȃ��]v,)��I=�[ڟj\u��T?���#2>�#�o�R2�y�s�+�ۊH���9����,�P�@�T�^��!m�����pr]�3<���>Z�/Z�I��1�}e}��2���>N�?���>1JlH�h� �)q�H�xIRY�"��Te�QhN�i�{��Ͱ�Tzqa��l�`.m�)���p�r����\�Ʒ��i���Bz)e�I.��\�L��H�>�>�����E��i#s�}A֟2
G�� l�����)��E�-%���A���K��-���b��(�����QsUw���/�֛�lA>��d:�g�H���a�i���4q�Y���\H`���QI|��M���\����؁Z4&���}�/�A��_�Q�k�m���Y�����ʐ�oS�-Ha��"0��IF┾7X�%��'��%��ߔ�N����l�| ���Z���W�^�	*\�>��go(��Bs0�к'���S&���N>�����:����Fy������~��g!j����Y�k��DV��aY��͚?���k�w����;�Ȝ�����?��2����tg�vH��o�y�L�%�к�T�s��Wo���G������I�R$����h��nn��M�k��>�O3��!{C�_ٰ/j�Z�F���y�3��Ҕ��$����X/���w�i��`�5��N�f]K���C�Ͳ즿h2Fc8����s�]>LT�"}�y!�J���QwPF,Q��.u�����ZPN�N*s�q<�,�M��#���&+.�d���O�m$��;u�q?��u|(�Q�O,a,�I�@a��v�6�Huv�Yw~��EA&����n�ڊ*6�w@�?vU_*�e
���oyDִ����?��h;:��hn��pQWR�'X��ϥ���S�g���o���+��W�;��u�R�=}3�� t����"��h�]�iζ��1c"t���<N�B;�)���3���Q��z"�]���f,VuK8	�����}֍Lfo�X�iՋ~�<��h��&��F��,j�I����}I._U�iθ����W���\,��w�v�.$�Ǽ�ʾ����BG7�yMdtB>W���T�����0�7�\J�3�Gw@y����!vhD��5�l]�^2��O�_�~b!�f��&�|��t������8��L�X��;��e� 4��1޲�YS��؍|���"w��	����gЁ������'�:&��� ^��3Sgr��#��1�^�w�G���q!���z���ztk] ������g�rC?��~9s���-�6"3�|Iz"�cAʖ�����R�KH:��P�2KС��c����4=N[�H=�\nt�j{c�Q����ͬ�X2�5^�pN��B\�GCo77���S
Q����c�8�b�e�7�؟~�/�i�M��׎u���;�h2(�b	�~I5��w}�B�]$���T�O�3d�s��"��jQj��a�͚�J��}��2���rZ��r>�K��y��4���Rg�b�kż022�X�ۘ/\�"�� .-86�}ꦙ.��U��\k�(���i��,�~3�����8�,QM�����>�����$ �6�~��B"I��>��4���<��g0rpWu�	���V�΢�C�V����R��k�g��*%��@��g���gU
BO�Q�r��'��4>�3� ����c����6Ɩ72�9�+�$0��f�|b>�V��^p�����(o�v�ብ��A7ӆ���=�<Vf���%٩�c�;��c��YoX��IUL!�ϔ@.ޛdsC�R'Q�ǑM�l�[�Q�\���Z�:Ʃ��W2d}L�>'"ѧ�4D�4�jb�ShM^�|�Ƥ���ҍ����ޗ���(�@T7��=:)���Ф(UѦ��Ď�B��X4@������u�J���	b��A�.�u߆�i{5������V�Bz{H��5�	�:�bc��@�QRs��hj��}2�4���ܙ�L	c�/�M*������3�)� sTW+�MW8H�`?ɼⳟr�ι�*bJ�1�yE\�����ः�����~����|�J�gċ�O�����(+^�l�b��2?�j��N-)�KQ�,=�ԣ����!��}n�( ж����IC�j�������UbBͧϜ�O'��xIK3�,�.�`Sw~�p�ӕ8\Y};'��U�}7əBvX�Uͨj!b�+sY���:�Y������=x��?�,������H�V����&&�;�2�������i�g�"�����E��.��ȕQ�K�~�a��NU6V�<�>��4c��aD��Ã��?�ײZ�6�@��=(̈́ L/�g��H�	�>�VHBf�e}��qƲ=�T�ޛ���I�?�)�F	t�:�a��c�o�,�ä�T�xÓ�_M��l>[���
�������v'���~�~�m>Ǒ�.��vbM�0~���Z�R��׋����]�Mˊh�&���Aj�%�1|���e}ٲO���<�G8܏�d�s�6y�V_%�l����7�ɂ���c�fI�,��$���/$W���!�Xr���OL8N8W�$�8��F��[?��Z/�/�H����ABp�S.��jr̂2D�3�0�{B�E�Q�G��)����e(��"��l��+�'��Lx:\뺨0#�,�wM��z�sy�3��=@6-�\�����g,��ğ򩵪_V7ؓ��K\³�SE�n��()�24�U��)��U�����2oh>�y��}`.DM����?��d�(|����I����:���~��ձ�˱�˯o�Sx�o�W����ä��G��Ì��=i�'�����$P�?n��[5#�!b3�y���f�������}ݕ������#�;���R���{�9���;QA#�ݩ�Y�ߚo���>�y�I���D����
1{�_�	�(�N����\�.��.�9{!cOF�)x�?1����{9$��7ԙ/q���X�x�}"��;3���-���O���
�\�|5��0���$O��TCj,{��2���86��-�T@�%�ɝ�W�"z�>[Ys�Zy�W�����U^�@����lB����~S���'K��s�G�0B��i���}[��JH?��?��B�Y������*�J&��.�(�R�~V~��6���h�K�����\�6��,�M�����!�6]u�3���A��M��-��-�@8�����
����堐8���ZB��M�X^;,�����O���@Ue��(�����nf'0;z�	���Īv�/9%h�ա]����#�&�!�����Սha�υ>�Qͭtx�_� ]�������^�-<�F/u�P�_�%wC�������B�wt_?��ަ��!Ŀ�F��&�C3=D��Ҟ ���h"�AWc�:�C���>�E�fk�ZmJ��� rQ�p�� -n����i�LG�T5j9k�(���;�(x��qỈ�N��\�@bkt�3T�i��M����a�cz�������x��ۼ�C���F^���a�'wt��o���S]g+;o�w(��i�;}�E�ȹF*�<+����n��ᖱ\}��q#� :vJ�F�e�����D ����Y����#W���PV#SSA�6����܄�:�4�U�e���z�qX��_[�aA�{)G�)	��Y�iw�L�Lk{R���8�߸Θ�N�:�;�i5}
&�W��:�y�<���\�Y���Qg}?����q�;@�
Q.j	[�O%F�t�L��B�׺C�ߌD�n��P��jq�"������}RdE跸��-��5���e��sA��fAS����ڗR6�AL�_{������K�����~&ev�.=�+=ƭ�D@F���������}@\L��@�3��0?s�K�� �T��.U��I���l��e
�C����3�P1�r��f�+�)߾8O�u
�	�
��c� ��'*�i��$�)'����Xd���M|F�T,�Ԕ�t�;�� ����.g�ܺs�����澘�� 5;ãN&����D�-��<�Ϭ���S��%��c&_Hd���)�����}1���r|�����ԑX�4�O	%��uW!��Z��u�q�'"�[ND{����2�˰�ZW�����Q�'����"����L���t�F�%&�F�4�]�I�#�_���D7z 3����>��븏�9�t�W9H\L�D��Y�e�SF�ρR�t�AV��0),��L݇6�Ѻ������:Rٜ��� 98P������j�2�Zq~�^�	�d�����ZId�O��m�TyW�� ס�~ʆJg��u4Ԣ{�%b�j��aL��.��8�ﯤ_�^Dk�Į�yÕ��N����E
v�:͹+�O�A�&ZHPC����MY��:M^ ���"�ɢ� ���R�T:&��({E�83qt�u�y�)����]趁�����8�JYL��E8z�����'��]]@��CA9�������hOmM�Vb���s� ����#l*��Y"ҒS=�De>Zomb�a�m����l���a�6�耳�\��+�1X )n���#wѡ9�y�D��G�d�k�]�!Q��?�-���ze����1��[��LHc���MC��Z�S��mT��ڜO~͒�%4��<�<�ۨu���4?׏F6�:!X���둵�F��I��P�]]]�RA:��o�]`f6�'c�9
w/���(����];��y0�5 ~z
+LN��>A�*�.��җ��-N%���ŭ�4P<���6P[�Q�p?$�FD��h.��:���D��/�Ώ颾�2�T��`�Q�mN��n%���̮s��y�%���S ޳���C�4��'�/*b�A�?®�����7�:��2�o')�t�.Y{^"�T	�Ƕ����$�e�	���e��an�e��	P"4g�:T� R���^f]�V��#�B�M���xA�=�J����E���0������:c�[M��H�"q���~E���wnL
�=�pQ���M�j�h)�(��V=01�C��������!��Q��]s�Z���Q�"�����L9 �������p�wMc��:�5O��Զ�C�	;R��6�~��k�Q��٤q5�wVTj�-���������ʯ����U	�``�J/�3�Kw?�Lu���2`���Ї���`;�f���#���>.B�Y���1ߧ�z{�]gC��'��C:;<�4:v�S��uC����[Y�𨗶|�qq�n>җ���v./�2gnMf����aT����Y� @�x�����G� �"L�5R�&}��Q�+��7��c�{ ;�6Z�Gl�z��ɔY�]QAk੢]��,L��v�����H�K�)o��e�-��JC��e%'�O����G�k��XÓH�ΔQ�5�|�S�m'��c�y����`�WI�7� u�9֯l*�M��rx�VsL�g����&v�� (��s�n������ؘ��m��kX�:X
����K{���
wk�bK���΃�"�rl�嶿������9�\����ݯw�������=B��6oƞ�ꮢ׌{��<^�P�����v�A�y��_շ�r�o�̈T8�	$� ag����gj�.��\�v<�v��,�j{���_��KE��V���;ͦ����b�'��'H��Rbq&S3<�mc�wI�\�_�}�+�n�H�Ŷ��;�4k�Dn�+\��){�!b��gvmI�($�����D���V�����yc��zȄ���2�f�ﺢ�� y	�4oϜ�=�w��L�e�,��4kI��>}�����5.cߴ����]���CR�iS���o�W!����o��J����gY�i��L���b��x�C}����9[���PE��֙F�r���c�������&����a$H�@{/Ґ���!�����p4ln�r+BEw�}J�?;c��t���K���v~E��O �na���A���S�^���6�
Ů�|��{��_b6�.r�"T1$B$@�T}���B�����Z'�ag��R��R�7\����Dwz�+��������$F��"�Q�u���҅�fW�������	�2�%�Ȋ�K�W���_��w������/6U�u��XT���8������ T����s�n���,�g��x�l[�f��a��F@�N�-����m��$���'����f�Kg�4%���w�+4%vy�ޫr��Ί�C}ي�J�i�*��1�3hq��"q���'��������+��S��,�H3��g���B���
�鲇�e�f��������{����t�����M[3�_�^tE���c�0����=�$�L��t�[J[P_�L��s��&��zi*c_�85|gŔ�o�����3̦=�AhQ����xiv5��lo�����)'��Ͱ���f�w��&�s��,��L��mu�+�g��2�āU�����X;����\��_ٌw��+�Φ+����H�&GV$�7�0�N7�~�����N�7����3�%�3��=�t,d��%P�1�f��\�UnƝ���$��gfT���w+s {�wAy����C���1��\�8�Ƌ�^F��l?��X�uY���J�;Ӡ��CW��3�����*r+9t�L|��U��̡����CZ#���+bE�N�~i��&b��ٲ bzj����,�%#[gjz�z��j�R��Mt��e�^CT1Z�(�C���n��=oY���Z�x#�M}섽N����c�j�<2*�)s��kO�����+�O�*���d)�ŠVՠV�N.�,��Ы���^��^q�v?��I�j� z��_9"���Ы@�^ W7��_�'mz����z���L�DA�n��}A�����W���/�+(Weѫw��UzU"���;O�|NI3����?8��iEJ���
����lz���)ai���rH*+�0�ެ��+���s�7���2Pַ�M�u�Mx�6�wDoM�"���k�.$���eh�uI�	ʦ+�f��I��#	�
y�����MrcH�pſCl޸����`Ӝ�?��o^'�؋��{�b����g��Ë��0�c>�7�p��)��Ϗq��n�M�y���Ѐ�k�J�_��~��|���iG鯑�_��~�}��G���qOa��Z��4��sSSb�O�`��v�>���o�ӯ/��S�\�ra߅�{<�/�[���	@��ұ����@*4�튰29&�1�ہ��$���0��.�(݋
x��9/G�����0D�4����9�o�-;a�E#��!T�����i��AB�]��鲪��GH�e�ȳ_���<�d[P�^��>v��h���`�����;a�##��Y>IJ���I�/r��C$�jl���5Y��=�u�������>d�#:Qh�4��H4Dn�Ԅ�K�����5��������P��Jt(B�2�-�4�v��:K�/+��� z6D����S�ǆ�E�(�#=Ucs"�{��H�\?H�3��O���r�U�yc�G�o|�Ѥ���JS��Eֈ��;�Ĩ�p�r7�_�i���Jw��2���+P�&��o�	���?Q����`>31Ү9�S��.�VF����4m���������O	C��m��I���.-oG�J�-�'n�J�Q�ZIW���Ȼ�1z�*e����N�mW|+$����ҝ����ۂ���N5z�}7mu��;W~����K�ð��'ZB�ZM-ʖN���[���Pb��?��Q�v�I�uLi�'�Q[��k������Y��#"F�S��-��lh���NzC�����B���4#7����5������=�잤�8�S|�b������h�sQ��f��9�>��;�Ď�0n�S���o���\�4�sEH�i[^V~ߺx�=��_%F�G��ȴ���t��U�j��`޲rw֘ZtE�CY�����p�G
(������$�r�����I�=+cz��"3�W�u���q����������-��t����U9Ue�59t�m��}��r����&�{���R�w�d?Koa�Q��t����o���y��e!�KiL-1����ϳ_�Nw���%B0��8қ����T�M�1�%���>pz�wvُ�	53{S��E��;�|�f�S"쓦X)L�����zPX�qՍ�Tc�͏�]�,ɕZ1Q^n�1�L4�ep�qJ<O*ͻ�;�L�����G�#g6r��r��,�|_eŀH�jC���Y�W.Џ���}��7w䉒7b Ϊ�%�نy�93�M�.��/��,���䜬�5�JADy]�v��MQ�c�Blqz��4��{���9����IFU	J�2��`<��JK�0<̖l��$��d�/ ����8�Lb�O�q>��mP��ꃼ�D�Q��s�U��"�s���^ń�U�H:��줣��ՙ��aAu�hk�p�	��;�9%�[g�/�'�v�Yb�!k(�4֝$_y��6d�R�U�C����Ý�So�O�R΁���FY[Ȅ\#�[�74Y-=���|����(�I�^t+��"���ia�4�5��3��e*�����H�F��2�l
;/: ���ݿ�.����`gڇ[e6�6)��	5����{W-�	O��j�>�6�R�C�v��	��4;ec��ɸ���}L�P��-�4 U��G~�-K`�ns�<1NT��-xS9��:;{�x�$�2�`}HQ1R4J����9��:����x+�k�^�[���q��,�g���8H;vڵ�`���_��!?���B�i��ܑ)��P����A|��O�-;���p8�@��8w;׷*�ә<������MY�}�wB>Հ"H��&2�J�H
̝�L�~�M6����{�O`�6�y�3�#�X�}2Ж�n=��|=��W�|V����=L�9�H�lK���
�kG����N<�U��}4�mnZ~	��r/�e�إk�h[n@�8���1�_���4/p�r� ��mҏ�.�N�I!pF��mt�q�J�{��j̩�7��ג">/�]rqW=�L�7��1��ϧ��d�t/����72�\�w���r8��Cא6tkC�>���{}!c�;P��G�UъF�4#���tv�5o�(F)�@��+�m���h��Y!��/!�:X}�.�w	(Xi�W��*{���f���r{y*KQ;"�P6�ی6@g};Zm>�L�_�Ŀ�2�� �3k���Nk}3`�)�1n��+*JAf'ѱ�[��ӌ*OT��+�$|�����e�UH��ۋW�g��k���>y�I�б��S�����闛d���ih9w2s%|���t0QSG�V?@l�x0��k�:B�>R��	�|{MA����#�v��D�FOLSb��r�GH����qn����8ӧ�r� ]ȗ!A�_H�^�� f7��S�9u�-�"S&�Ul 2@<�%09А����pI0��tg���t�'��J�l�[��F��Ô��Z��S��J��Q�ϕg��܃𘫱�j�ñdT ��Н��P^X�/����W��|(�Tf�*y�ޅ�Wp��A�9gZ���t���PG�L��:�jTW}�:����p7]�ӆ0�J��!���5������qH�
��ĢH��n�p�5hyU��yLH�U,�2���2���|�TQN�bJ��e5���ȇE2�('�yA��~��hYP2���e템b�U�+=J����6u�'���=Z���ou� 49�g��B.�.��j	_qP��|�����.�!EK��������u�`��U�k�pU��I��=!�:,E%.a!:�}^��Z��azڮ��u�~�hg��q(�@鸤�E?s�H�< o�=�h:*��p���ic՞Vw�C]p�Ƶ��&�A%�+�87�� �[`r��φ|k�tq|����m�4���_f�l�?84ag07D�K����+&�s��5��:<m������F�Y��#4~{�@�G8 -G?Nⵍ�(��NId`ٔU�U�n>�^QI�\�&|΄9K��.ݯ4Q�Bxj���@~��t��PH79a����(����}�����B���y�ho�d���T6�?5Y��0溢�y�.e��I�z�$;����c�z'�D�ʱ
G��{�8`~�4��K�]��k^Ԝ���]!K-6��"�ڟ��v+k�مJ�2F��t<���Y��7$���I{+��^���a:vg{�r�ؘ⍖�^,J�������t�CJ��GƯ���_��Y������=?L<$ɦ�
��7�?�yD
�/��g����#�2,��	,�w3���x���P�0�ګk�ʖ%!}Qqc�o�ϡk͘�՜/���M�YHApk��{	���F�V�P��贱nM�-���e���BF���}�v| �_\P�N7���J��uHh���*5�?.���09�Ǘ�R�+�L����,�=�fxL�U���Jl� ��ic�h���L�	�G��r:�@rd"�C8^L+�jƩ�Z��HJ{�a��6�� ��Z��)���:������j���D�˂}���j��*�#�#��Y�r���x�ǧ��E�Ã��C�2�w��u�@X8��ig��`b���u��?�&>�3G^�|Jz|ޮP�Z��ĕ�[ʺ~)��,�󁮷5�64GC������P�q:�"�--\�~���{���p:c�13}>gN"��m� L�]ge��8�Df�gs�VC�&� {YH�u�@�}��;��9w�uљ��JzI!�UB[�'��{I(�>8&�/����u���c�}m�Deˬb���|�C��D����=\N�	c�OQ��Ƣ��$y���ic�˦���mDk�v�eJk=כu�F�&����U:��#���*�?�M!@�D-Z�huU���yi���M�H \t���R�%���`ώA��s���6���9����RQ�"��CD������y�I҂�����=9�9�y.��s��`գt��b�/�zr�%���	P�l���#/�Rtr�X?�v#|�pڇ�>%[糾��y����z7\Ԛ'ɤh��8��9�Sܰb��X҆�̕�~��l =>uR�O��P�6��zPk=��6�ɛR�i�l9>ez�O�䨘�0?�#�s"mAwkO.+�����Rj�v�Uj����eFf ����Ě�PB���
��:1/��z��pd|�?_���vz���ޫ,88��G���뾷w�?��W�O�JDI�W{A���)"��ON� m���bs�<�0Zd�c(E�<��CY5��k��J�ʛ~�c��ta����G��"w�k�G�-�>Rw�k绡���	'�U��=�9`t�ctd��;��H�J�����8I�_ᑛs�M�3���/��2�����缱�����u�4�:�����!�wj�8B'"������W�����!��@BX�+~;��oi]�ۙ�yc��F@�+�� :`�!���o��C�S�'�3��6�����Ef�^�Cl����ys����rI6M���8ΤO�H��g�5�>��}(�&P)Im�ڿB\z������#�����q>7:���I�gw�ȏ) �����P�O١�Bb�1��ͩOT���>�1\u���\0S$�����9����Ur�O�0@2u����(�,��ݲ�í��!��[h:�sx��*�R��1�t��X��˗IUzc=���Q٨̈��X�A�٠*�3��`�j�s���C��L�_�t�O9��m(�!���j���l���������\�Lzq�iD	N���a�w����q�x�+���G��:��얢���<��D�8K.� �+�B=���Rt4}C?���%�d�q5�}!��A"A#Q���zzN�C��L�t�bV���Ն"�K$��s�}��C�Z5�>�,�I�������vH�ә,Vr�ɍĿ2�H�-W�oI������qN`��qZ�+E/�18"����8����I�"��`�%B'O�h]{�n��;3xV$h9��RZi��q�����؏H�����+u��\����~~71�;6���i!��϶|�i�{D}���+��)zOPp`.�'�@�f6�ᰪ=�R�i������M)�;�O����� �ؿ�
K�K|��r�'���*�/�~ǈxe��
���*���{�w�S�\��P�/Y�Z؈�/��bƕ�	��w���;ҟC����f
F����N�s{��V� V�p�P�J��˶]����������|���L[�Q��0v�1i��m�:��MR���J!�{�U��K�>,�<��/���p��4(����V9ۉi��$��n���V�U�����^$P�靪���h�����ԘRt��#�9S���u�"�Q'�Q�앝��rq�����G���~"�=�4��q�0�����p�r��H�o�>؟����i�Z8���YH[���W;�ݡ�"qjY�?>��	��}��fI��?��N$��-U�jۨ�΢C]guA��nE�G�O�T�Z�@4�����pB0��J�z=��h�>���/?*�=�)(V;Bg����t/y�#�Vwfyt�&d<,8����!j�p��+bȭ�	�I�w'Wg�v�J����t-qm*��mkEƴ�l��z��H��4>t�P$Ģݙ�W+���ٟ�gu|v���>�����|v�vho��d�>��⧗K��ºm-Ug�H��%
o!���(��3
!\�����C�������l�2�ސ�I�z��9�9� K�M�pKC�4��[���o�[Nd����g��2�Q�t<�CZ�4�I��2��9"P/���z��o:.�������x�y9��	ˏyGV	#�����!����W��F�I�p�U��$�k�*�\�=Sm�6s��ȁ�O0��V۵�c¨Z��m1C������D5F�A�����yfKEN��6 2k5�!d�j���ew8��ܥ��"ie�%b���~�{�[��$$ 2�m�g�����ol��T�����8�k*����cazgׂ|T�Jx���׃��k��u�s��~f-y]���w�G<��r'�c����u D������^W�V�m����d�C�	����Q����^#4h��*gM?!ğE~e�_-3s�b�rd�l1]o��
�d\��9bc�y���f��άXH?��#TP�˟����p'{��������X
��~�#����"@S��Hy�T�k#G ���˭��ht���dcc�G1���(lb�~�E��Q,�Q�H������Mb��>8U��V=�gCN�NY�3�~���ؾ�]���Y�HG2��#Ѭ����a��(�%G��[���1���e5(�f)���ν��,+�`h�~+�u���gC��*�H3��#}�:��W���j��,~���h���"���?P��
��f9���M�1k��%R��|Dn��"���0��@H�J�#�\�#�l�+�E�إ�?�ǲO��z��c�h?p�~��	N�����wx��Fz��f$�؈[N�X��6��c�.����<nd$Lx�OB�|uHP5�F���Y��Zalv��P*���~��a�d���r��I�f��'�
��B��>$�i�<�M��{��c0��e}Ozqf�鄧�J�g�"���i�№��*4&j}~�Y�|��ه���Qφ!�R-�p�6�A�Z�����]Vw�3܊|�Fi���#ie��~�O���4�SFr�ж��A�"���hj����ȧV2k-���ղ����Rk��d������.��i�c�NE#S�?
���|�w���D��h1�I��G����Q�҅&Z#m9F�k�ԥA�� �l)A�둼m�v��NN��9���7�g��Zs1�}6�ѐ��D5SN�z�\��AI7wF9e��q�®<	Q��".��ؓx��v$�o̡]7�
��	Vc��y'�.��oY���۫h����A�N7.Q������F\˰#�~K�p��#t�sTa<FU�C�lZ|A*�%��"f�(�6e��L��[Q�t�ŕ��vX�QƔ2z�=%x3�������Q����)��4�n�!4y������Y�<NQ�Z�'eM����k�أP�,��0�Iĸ��(Vv��*t!�<�rRn�"�5	J�+����U�_h�l2�G�_163�w	^ 7i��cD֮s���M\8P+�[n"��օs{�XDA1l1g��M�	����b��+c���k�f`M����Ŏ0wQ�Xa�.�aY(Ů�vf�,���Em�R]��z��/���՚�Q vm]�H:���Ň���z6�
��	܎�!C�)��� PdO�����-�8+jT�v��/��_�x�tųUT����,�a��7�����"��,�e���rls(��>�u���3�H�I�U"U��׎�Ǔ)NmY$\^~�r�Ev���p9OY��$]P�v3x�#F�V:$_|�M�!k�6�����Xc����N��͜Mb����T�oӜp��\Z&�`�M�F��i<�m�_������	̟��Q f��S�D ���n����V"������X{��[��*�rS��g���W�Kd�.�j�H�	fU 4��G7��"�y��M�����M0El��!��S=�!EG�za��^t�;�)D{]6��F)�wj���Gr<XD5��h��(������kr$r�8o/�m>�Ν&w]�
V���MoC�5\%�M�L@�£Rwe�(~X�nt�'̮ o���l����"����Z�"��@|X���� F69���_�ՅAԿ||��[�S��9�0�"��N��Ӯ�� Uc:������)��1z�#ݪ�!)f!�V�.&\Q�@��C��ADy�b�N�"��Qj��? ��A�� �+6o>ϭ>2i$���f�A�&A̢�`�h˿1�����YΓ� �FU�K����Z12(�xt�b�i-@�յ"t���@��4�al��5h!�o��M�o2��oO�%�n%(&��Π�����7�7�r:O��g�T��p��� E����Rm�"l��Re�v�"��!@���Mx��"n���Z�2�qz�3�������y~F/�T�6k�s��h�%�ك�1���Y�F�_�L��n������ckv��8V�Gt��ԯ��}>�2>N yl��W����fj�c���Vr��0��/� �� �;L�/.�������n�ϱ��%�A C�0��u�e�I����۰��˿N�����\j�lB*���{�fJDg������^z]-��/=>i���M���O�q�D�l�� 
|�^.m��q�L����@���B>��:̼���8̳PO�x��,Q�o�3tU-��C�	{���_�|�j+�O��s��7O,kC���:G����6��Ͳ������Į���[�A��.�������n��Q�9!��f������I��hu�L�)�>t5ܣ<ɸ�D[p�?>�Q�I��eT�ז-�S�rX{e�A3��b�W�{��&C08�?�r}�1]�^Tyg=Rh�	�f?��K���#SF:����[�)��
�.Q)�W��h�x�)z	[�g�,a��j���7]� ���7�$� 7�A��`� �TVE� l��'J�xI�Fco-�h�� ��(�?n���M�2����X�8}ԛUOM$Op�Q��jGh,�'�z����J��KCꡱ��@l������&��
�.�w�$^� ���#��߈~�N���M�|$$6Yl�=��w5D���|��h�|[w��9��2�"/�^J��a�bu��c �Z�rjn�r����,ؤu7h����޴L��4e}�@�=��II�B8�`�v;�j�D��#�*eW��������zs���_Z�4�w�vs�Mj��[X�b�Q�A�$c����
+� �ψ��!E}y�=�4��ߓMb�'?y����#�i�gu�i_��Aa�S�Jc!�K��������X�O�\����ψ�.`��	���L���K6x˺����E�9�gSV�?�
��gDg���{ ��3�i�y�!����y\���������Fj^�mĻ0��~5j�	��tĺ"iu��0蔑�R��vS+B�m��V���E���l5A��j�·�bh�ӈ	�*����_��9� �G�����64e�nt���e��U�19�#!�M���3��Ej�������E����^_�ˠ��w1��%c��#9���
!��-�9�I;l2i�c���/���	4�b HF�����y�������eG}�(vJ���ǭ��֖�(���b��������M�[���ɼlF;#E��7�m��A��q>�Wj�*���fH&a��~�,^E�x��=\�J��&�5�T��$`䮙��b��X�5k�ư��ʜ�ט�vڝ&#��4&_0r q(=����1uq���{�����a�q�8;�~zǰ�W>C�s̞�r����}Op|����J���h�0�����S�	���*)��nө��*�'O�� ס��V���X����S�՟2�##Ⅸ���ց���E%�r����<��+�S�D�)(�x@VOҚ��E�KR�P4tr8���;�w3�й+�li� �9������i3��e���T뿞〸>�C򴭯_��sRޓ����Z���v���"�V�$�8I2��Q�:�.��fl�����+����ml��rXO��͵x�s�Ej���H����,��[�?���:��N�>�ڸ�-����x�O����+���=~�e�p���6=�jƯ��݂ ��Ә��*�\��Բ�;��Se��w�J"���ݰ�����%6cJ�� ?QN
��5�Vms���(�]���ðdO��p�����K�2<����&�YYR��b�|���b��44wq���f@W�:�Tk�c����#�[K�����J"�Bk�[�����?��Oe{V�F�Lo���4����4����;�/���s:��<���?9�x������xR�	��͍�V��V�Ò'��;OE�")��%��x�����~1�~$�l,'XB�=긋�����pb��$��#�8�F����M�Ih���0���;�
X5d5,>���֒xnd�z_��7i �����;�)$�pШ:��,!�Y������+�ƴ�U��^M�o]�}o�@J?7]_�Rc?ܛk1�DL�W�/5vݦ��g���:��W�����2��������"�ڀ'%@�t����E�Q�m�ԭ�g�PW�"
lHn2T�ϩ�����*Y�h�#o�L�Fݫ�����e/�Ȋ操��rd��ު�KH���cTw��������3-H�����v������\��~.v����)u}��(���*�W�#��W�pm���!1ڀUN�p�mo��Pl[U�~n,����i����x%OK���/���qZ񿭢	i�L���g<�2O^ZO�yHV�-���|��l�9�"�_�Ȫ�[���XO���h�;������r�ߞ��;e�ʯF|Ih����v�D%r$���(�8t�����0MO����?+:��z��$���a�c�n�Xnʼ��W�xM P�_��*r�i���ھ�H,�\V�*��ؓٽ�mt��S��#u$aOk'<�W�>4���k�kUr�U�-]t��˵��6LhVj�C��\HM~pQ���ٵ'�����j���TJ�&��W���zE��V��4[F_�WiR�1��F�l|�L��l��a<�;�k�D��`��&�yO.�dw�I���D߲}���*��z�x���j��EΪY�#,I��<�Dϑ'��#=]I�m���	r}%�|{eu"@�݈��p[I���o�8|����H3���M���rd�7�y�ndZ�0���o\����<q�CsRc�y�eJs��dUցL����B�P?a��ݴ����_�C��?�ԣ��u���(1OJ��Q����vzc͝G���o�(�h�i�^���[֭;��Q�ͤ���)j�1)ʢgO|��U�����_��j�^�DG��#�@
�jU��:z�δF�R�RYŹ�"�[$O/^��>M�ݎ�vrt}g�2���i{_)0~;=N'@^���*n�tl+i;����i��]��E7�_Sc�29��Y�s����`� 6Įm��deuX �ϯ�/��y]��D�W�/��l&v���z��>��+{��r�5\�r}�ǹ'�9>i���ףz���D�%j�S��L�yƦ*��C��>e�DR��k�-�S-��Z�2\�r�k�c�|��B��y2�m�k����6�e>}`��N>/�3S�N�Gz��.��*�Pm��t�H�u�������}�e�Ȳ��=���v�s}[�6�
��<����g�N�h9��}=�P���(�B�A��"�1�,�UB��H���y+E��J�Ou�"�V�*u��$���(K%m�U
q��A"� �L�x�b���fײ�3xC�����u�� ���A����Z5GY!�t"<�ڮVd� ޯv�U3��r$�&W���]�W��ꌛ�GX�?�A	�3�QJ�;��"_������Cz]_�������G�[��%|S�#n����Q��>y�F9�V�;r�zjۡ�s8h��2n�:��'	κ�$�Z�>�حwͥ�A�&�
sU-�*r��Y�����})vu��I�H����lR��I�����=��必��t�+"���&�=OͧS�mm,�w+�It5��~��Z[��-�.��'�ҐȡNB/'w�'߰Qס?&?���$rr�R��Z1�O)�b���C�sz�`��R�T�]�"J���7d�����BO��<���(�7������md��9ힻ�b����ݫ�<�|�F��փ���A]�p�ԁ�����{��i�c���NTp{7��	��� �H�H~o痥�6����`An<�;��r�Yp��ˆ�p�vV���QZ�W[�,4ܯ�����x<%��<w�UB��ڷ���H3G{���y�Ѐ���%&z���H�)�O�:��H���:EtK(��0�O���y�c�ф���u0�ND���:.��h(x�k�b�u�4���)z�QR�F�:��U��ZCFNS��N�id�����qL"��b�����(v��)�o����lw'�L7�]�@Ӕ;қ��Xj�p�Q�q�*�;J�r�t��ƾ�a.���r�G��ڑX���Z�S�kF8�?2������S� 8(�v��� zO�]As�����䄳�ǵ����J��(NG�5HI�����ߓ���A�	&DU�v�:���X�R��V��2�QO�q��|�]I�W�j���g�e4�Iu��Z�����/�upw6���t�u]�W����Fv�D��y�C�@��A��
�����񫎤�pt��p�q��y>H`L��5lv�\:�>�ȕ�h����[&��!� >2%��	�����[P���i����r�a��G64�_"&&n�J��*۹���,���s	$��h��~;�D�b5��}����q!�|u�H{�v���?�2h\'y���*�vh�,�H���2�E��o�[��*]R���t��b&��Z���k�>�~!���G0��د�B(�rՠ1Ě���e�8B��te��]�a,_���胯232��*�(��<�8ŗQ��")@��~�񈈆5�ɺ:�a�q a���0���!�Vх}x�w�ù�|Rĵ4ݯ␆k��Xx�oj��1f����8����D�t=J S���a��@���S�U�Y�`V<)̦#�ȺM�g0�YX���x\4D犧ydM@�}"[�G��O�3�bF���~wa9�N�������C�
����-T�͑��İ����fb�2=�o��ʪ���/Z�wwcq�'񆴚;{�y��;ѶƳH�ITy�l��C%��y���ә�ɍ<7kV�������h�GK���Cvh����*��}=�.�)�;l(5�/ƾ�ƀʼ����!҉��_4�Y��ё��"`A|@�p�?�wPtU��j��dƤ�et�+� ɥ���|(��I��˽�\lᓼn/c�;ϋ4�EG3_�EJ[��䬔���a��o�R���v��]�cI�mRl"��O�,`hhHev� )�+~H��}
Q��#�y�-^,�b��g ��# ^��+6�������>�s�h_�{/���I8l�?ׯ��qT ^�p+������s5����̮��H߲�<����Mv��V��b�����lǇ{�^�"s���~e��/`PoD���Z�9r�ې�V҇۬�_�ꊢYv9��U�R��6���Rϼ���I4����x�-t���#E�K ��B�vo��F�;�f1�~��+������>���veR$��B/Մ[��K�sg��'�P6�Hÿv�ȇ�Sk^��e��&�^Z�S?C��X$VCZ�:���_�}�lY䰄>���E[��I1��7�Oe�Կ1Ȃ��Ah>�7��vM	
��2��Sא���F:��o.�=��(��O�)�ǐ�/.�W�4$i$����ԁ� -E�K��Q'����dm���I"��� e�,2.��_HC�"�(V��1>=�z����sl��+�)����އR��`�z��K���H:�N�~��=%^Q��}�n_� ��%lW����;��[3��98���My�G�Bqč�U�N)�9����W���ܼ�t�i��]�{՞��x���۟u����ه��M+����A��[��n�5'��V ݾ����ȃu�V�8eʗ�Y�ާd2zS#�'+G��D�����.'� R<�;����'w[K#��.�?�P�bW΢�*c�fk���a�@�K��&VF��;�P��"x`O�b�A�4i���J�Ge+�T���7�++_��}^��P�`I>Ik{6�BKh�&:i�8�03lw=~�s
|���v��[A=���v���s���Y��2">"N�o���[p�A+�s���	��R������4�&�s�%!ꓩN��]]��#����dz=��Ν_q�L߭lӞ0������bXz)��۷���=?bX9��J}�@�8�ţ�M��M'� ���Y�-��1�W��D�
�as��ɞ#L���J���8�r-{��do�۠�>j�V�����X	��n3�1��ʹ����j�H�j��졫��dY��M)�	'�$��U�pfh�\���e�z(�և͐���~S�Wu{h�W�	�+빚��L��=�)S�11� yJ�L�<N��3��P��w��8��o[��7���'�K
۵3�m�JHi�3;0���(=}������z�ի�2��Sv֯�(������N_�{Fh��C����Ύe���~��5kӈ���@�3��#��e=־Ի�F�����l�x�?c7�e�oM��V��q����b	<�i\�"T?�5*��U��s")���o��j�/�?�~�~nfE��~3t�h�v�~�e`�}��u�Vo>Y�?��<+vZ�wAHhϿ6exm��ߩ��i*���}�'�8�p�Ͳj������|�� �k_a��1�β4\�g4@A���uy?TFa�X`
m\6~%�Nװ�iy|=%�9�/�h_�YV�� W��̌Ey�Py]���x+������ߞ��I{��k��VD_�I�]X�ݮ�(ng���j����ܠM�5��h�*��Q�V*�9�X\s�X��f��|q��-B��_���D�ǩI1����7o�^[��_���b������ ���FoQ��e���a��#�\�n���3Ѝ/��:�y��n���������ov��z"��C�%�*�m�t@�I9��P���;"^�n�E8��h_<c�9�4 e�z�[�6�>������ho��u����zD�qY����ʑN�6�zq�h_�!.�e\?�j���.�Z�n�YZ���-�����P�2�X�x������3�ɂ"aPꑢ�cd�����W�ݟr�tZ���c1u��-�N.[�V4�J����*���๝Éϻ!HBt�U�-]3��W�m�W<�rM�Zƒ�i4�,�L�3V�6<p���z�7�/䐝�;B��J����j�'ٮ�JV�/D��߽>��8	�fk�0�sW�|�\Y&=��9<���7<4�;${:;���1\�=|�X��)�����&�M�=_�9jI�͒�iv)Ʉ�����?��OHPf�$�R���n���H���.(�nĺ�fX�����@x1�1^;�����h��>�� k��{q.I��9#��<�|��V?���nK+q��t����R�PȔ����R�	��v�����;��J�X��G�Q��a�V������^N Bm��Rt"�������p�_<�|��O��5�SnGʐE8�o�)�1ܿ���������V�6޳(����V6.�)�u�T�|U�=#�+=u.�t�(_@ˬ�K�|lgz�M�[u_�_U����^�����z����'pB��r,�%���g]xA�١����<�~��:h��+��[z�O��}��A��N����)}Û�}��jۭ�\%5�h�_�`�z)�N�Yl�: ��SE@�y3�#��0ҟz���wB�A}��sZ��n�r"� Z�*�hwh��X���$�o�:����	+~d�����$���xp(�L�2�����+�������㿅l���C��X�^\E+�2��ӳH�-R���%-D������C�cr/�1��(�}�Hy��AlaE"��oB&5��,�8+�����Z�H�~�]��ŏ�@�:*��>�8TdkT� ��*Wz��A��P�n�IpV�[#�Vc7�+'����i*��_�$`W_��s�p�4�П\������amY���	Ϲ�����C�֗����m����7#v�y�{f ���YH��[�M^��B+W	�Mү��"�ZЮ_̹�o.��/}�f�p�wEԈ�)v �qW��k�DZ��~��9�w�,�߽.O�4!Dl��+Һn@z�?���0�?�.:#�DY'��ˉ�x��?da7��,�_BD���L�a���Aq�Π��a7��̈́���%��H��{K8��<e=�9�'�]��
�����Vc����5+�.}�vY	!��6�zD��t����YzH����C�Y�v�Y҉��(�΅�h��ڈ)gM0kA��	k�E�DAamV^V��j,��E��U��JA.�{Ee�×��2X�M�)�ml 3�~�𪖢�s����\c[���~ p�Y)�&��'}��F��s�f��,_����[����H�\�0���ur-F!��J����es�,���D?�H��.ks�T�x>!>�*�Z<ĐN��I�-�NL��M +ک���0G�Sb��D��F+t��D&I��	βB+֘��7�G�ƫR�s�Ra>ˍ��p`%�v��/�zr_�WuK�lh�ń�4�H��8)?m@U��5�_����C݀2��e����ݲ��~I�滴�r�<Ɓ�M�}J�ȝ�Zp��iE^�U���a�x�o�xhۜP����%?he��{��0�y�<jc�l�_+Wsʯ�e�S���|(V�w��yr�!$X"[��;;�{	����H���281M�F���}�B~��߈,��R�s02@}y;Ϲ��Ѵ~p#+!im<_\��q��ml����@O\Χ<`$H�kD���4�ݹq�/9{��-f�l��.�y��?��� �:B�Mc	�b���&V��K�ҹ-�'gX�$ܜ�+�y�y���42�2�#	,75�U��X�'�#3�f=�?��)�%��� ~#�į�����G
�Cr�У�lnk��Q�?.���TH��ש��`�������i�YΗb=�I��$\7��X*�}���H�s@$�'�2]�ڗy�w�Fq(�����z%�Ċ�j\Ƨ���?��N�}����G�1��do�ye�"�o-)Ki��R��,�S�R�7Ⳏ��E����0J h���@�%��u���ĵ�w�:^$��:�G˪��t�z���'�$�Y�槱a �[@Ќ��s>�>�uIڤ���v`�}�CZ������q�6'�P���@��_������B`�r_�k`^v�@�/��u�9@ce� �e~�����ď��/<P��mV��R��c�1�Rc�>u�]V&��/uu��Ls�;iP��6S���x|�F���K�Kv��U�'��52�3���L�>5��6�h�Q����e{�}������������G%Zrt��cw���m�qS�/������D�?L�M�ǧ,-�o�����t����H��W�2�ԧ����vs�c_���5�s�'�bᕷ���AL3�tH����I}��ז�dq���g�뾺����S��]Ν��r��]K&��$B#3��.Sn�QO�7�Ȣ�Iu��V�:�/��O)�� �k��g������m���Ȣr��K䒕���K����ze�aٹu���YRn	�	��Ԡ�2��';;�O���t胴dU�-����?N�N�,vYBsQ�l�����@��JFq�]��k���f��Ʋ�e=�Ԝy�9a��|����	��,�\�/������&Y`2�}��i/���G��*�^U����[��*6*RmDX7B�b*wө����Z�HH߭X1A٣V5`4�"\��n��؉���/��-Ÿz8�J	@ ��/��z�e���J����R�M��@9����u��X �"�)�/��fn��&�>�IO'�&�?8h�c�X�:�LY	X|̏�4���@]O�������$�O��r����&��1e	��wj����������CI*� �W7C�S�܌=Q�qfQt��ռs֍���r�|����V^M����]�S�Џxޯ��T�6������>��9��䝃(#�K?b)�QD���kV��_�/EW�LSnD��p+�����
��¶��IX��Q��cV���V6q�Yv#�{-��W��;�J1��=L�����¹q�|(*e'7����Zo��\��x�[��/�Q���'�B(�їB��XOs)r�G	�υfcB���ť��օ~h>��j�E�b�TU�Vű͍��	��c{��Nt�m�,�aԓ��a�Z��`/�l{��/��t+�iү��=41��=)�Rj�(+'��{�	�U�DZ/%��-�G^J��b2Ϋ�n��V-�NŽwRC�LJ=��
�!�����Cs�g$�����_��|qw�?^e�}q��7��a	}���|�NX�b�|�s�5�3k=���|�~��K��@l�C�)U�
9������x���K�Y�0}��|s�"D-;euK1�Vs�շ�;+ˬ��)�&�A���vU�X3~U������Snua�_� {�-6��M��|��i+-����j;��L;�s~�G��G8�-�U���'0*%�(�rl���� ����J�'���&ŮO� o�9j�Om��̑�{
e���bGKs)JV	�R"��H�=~�,��KZ]S
�ծO�n�1�BK��`(a��/;Ɉ�zr@䆯�aq�+J����,+�����a�5ujIke)���f	FD�A��8���7��/��yԕfZb�"�BY�MLU���L�gĳ)#��B�Xt1���~9B�V��Q)[՝�
}p?t�~n����@���bx��F������Z�YYe�|��^\ZC,���AcQi�zU���#U�q�
[�/���x��)� ڄ���+�[bؼ�30�p���õ*fa��!c��c����<�������8U���e�&e��Ъ��y���$�@�:�%ػ�`� |���ӟYp�	]����뼄�%e��ֺܡ[6�X#�RG"$��i��6�Fw "�����,�M8����K��x�lL�ׯ7pި#঍�/Ϧ/��*�k��C�Z
?�PW+���++�]=�2c����?�}�Z��2�����Z�����Ĳ�॔VW3D�z��[W�ݑ{q�`C���m?��A��I1�^M����.ħ���$��}KH�E�Kxd2�|4xK�v�sm��������Z��]�&�������؉x���)K�ՠ�:%�>T�*#@��L��-ۡ$���z�������^�:(�~�;��'[��M��]��-=�!D����-Rt-��n'�L�΀~� ���(��Y�Ň�}gxI�y�v����V����S����#�r�o ���Q���s6rl����|E8:Hl�L��l�{-��N�ćɢv�᥺��O���<��ɯ�/��DV�/������6���5��즑��J��[kr�4��4�F(16)�;��h����~,�G�i�e6����r��y2Ę��^����yl�}b���J�s=az���w�u��չ�F�x_{���;���V�_�
@P7'�o�/��H7�rS��*�x0��ٿ�n*��W�~z}C0�q�닜ۖ6��|�θP5�?�⏆M�b��+rIE��Q�>��M>	_n�P�f�*e|j|/RR`��y綦Vm�؜ۤ�{�[������(���uGRi����p�O?�<J@J�+�ꬠ�ڙ䯈�_	=�a\i�#���Ů[8��BP����t�$h��=�f_
Y;3�}�%�Z�
MI#xE��a�,su��$��76�Y%�D5{�Y��4����o�Cˢ<����?�)G�����_��*���b׏���~�#���>7�̈G)���ȅ��u�
n�`��vm���(R��$�ڨ���2���=�א���_#�9�7vpw�Z��]P�p�1�s��1졥6;�'��ڣ�K�?�7]�D���Z�'l�wg�������e�Z��v�_��r�A��A)"����ө����s�T���+,�q�݈����.�9JG��;QI���h���&��&�R�|�p.c_e���S�Tbx�|� ��J�_(v��W��y�Q>�h,��d�oЌ��4�_�ۡ*➰bx��7L�q~uVil������� 
��Cz�ȫu E�� ��'kK_zyW�2�7��ZzYi4��:U]	Z�AD*�>t`�VŰ5��Z�5���I��=4��irV�Io�>���������)saC��ꥒ_�����Ya���ML�$x��[��oa��B��t��/�W�������[�+X%[�R;#1���f�d�m]~u��*�@l>� E_��л%sh/��dI9�Q��8�_y��+��"��e)��g��Rt�-b�� �[�*�{`]7��̗��GiN�1X�����󨞆YE���� ��so������yγY:��YA�Y�?�i$7�3��^��<�͢�>�v����ȵ��Z�N4ȫ�4><�o-<�o��tV���w.��:���H��E{oRj�T"�T�JL@-1 u� �Z|~��'�P�v���(����O.cP�� h0A@n�3��f�ń_\�����"�!>v��\�٭k�=�����Wt��z�G��{�5%R�T�ݞ{Ē���:L���uv3������ X������F):�fz�*�$�7�0�*kE�}��]É�V��oNAд�F��-�ݑJ;՟QK>��QjK<ʮN�9V��@F6�5�|�%�ge��e������<���]9���#�Z���\Y=%�3���Fe�亪|9^�UP������??��._�~k[�'���ա�ƺ+�{1�=n��I�_�o�=�w���L�e��p{*Yb����?&pOT���p�]T�|���t��j؁Í���ϵ�w�m���^ݟ�O��9#eu���
N	����Z�#[���V�]�R5��8��>�J�ԍc��K��9���+�V�_Pe�,�Y���v��Ի�o�Zcm�^e�]Z���`�i̬�O鑕�J����9����ۡ�t�^!�������'F��q�G�yXW�S?�K����#y9�^h��lr�����3����|�7�R�3,`�F��[q���SȔ����Z���0�W����� ������[��u�n3��H���LǾ�u����ʚ=
����B�����+��I w��}/и^�2��ڵ�ס�&wB�4=���e��}DD��0K��.;E/(A��2\��Wj��|p� �����tQ�v��N�O�����6�CzjF8B?�|X=�Vh�W�]}�c�u�Q1�=4���12�|F����4��/���3a;����־ڟ�O������Oo�Q���W�d�h?��vܖ��n=(�o�[h��j.���S9�iA�� ����%�du�V3r�)��k'��+ȥ�9�#�t�*�q{�V�M����&��mb8�i V��2��&t����<Ϡ�����Efy�D��YGnJ
 ��{68B�a1�� �$�)Ӄd�*���t���鏓8H� ��Z֍Ex�a.����c����Ŋ*�𾬇<��߰���~� ~��Mw��*�l.���;����mDf��՟cY�d�'�/����?�s�b)}�N.:�g:���	i�G��K��̰X��Ҥ�ؒC(��:�U�Y���M�7�r(-�ߨ�_G]��2��W	gH^��V�sl���(�Q!�v��k�-n���û�1n�V6*�P4?����v�V���١��/���8�GTϑ"b�����Oa�������_*j34D�`�hD�^1"1)�Xm�z��å���T�̧J��G���@�o�X��(#͋�w��������?�\�سcM��ۛaV<�;��ĳ +E��eٹ��zcC@=E��1�t�׻C�[�`������A��� �����S>R��q���ۉ���ׁ�]vM)�ɞ��l�Q�?|n�{�b_���]����S+	�N/��ۑrYZ7�֧>��	^�Es�ҋ�.�)�k�J����9ߒj�՚�΄�!U�7����̞#ݿx4�k��!���u������nH�Q��yF�0=��e�Uq��w��P������r[���~b��fϔ�?@Wξ��p5wj��@�DM-��r5s���\��6���-sa����UT`�:Dҋd\n��u�lW�3/A���z�[]6W��#9�����Q4m�7~���K�gl���*�vu�DzG��/�K+B>0�[5cZ�g��	�9w����r������	���8o.n\��G�%�C�@��YVkOs6�P��_@�������=�c���Y3S��B��4|�j�~�'��ޠO�� ��B�[H�8�D6�U@�=f6x7�*��X������?�r��Aѩ:#nqX�L�l�V]ٟ��O>l��hd"��o���^��7��W*��o3����QC��d���k�'2?:�D`��ל:R�?�K�,q`�V����[���p[����i]7����VV�~O18k�;�����7{�ҝ��n�?��F��E�Ȉ� "re��5�����nN��cby$�#K�0"K�"9��>���W��p9�\��/*�>�M�4�Od�khx�����M�0�#�oi)�N|d�Az��J��ˈ�1��2D'L�Un?<�_�U�^&��n+o�#�Z���O]\p�̕V6�����]i_������(�bi��Я���o�&c�C��tK��.�rq�\�I��$5~�\�C�c�Л�~ϫ�.m��mV_��#��ey�`�|�����v�3%��������?�Ls���|�;�W6J�]j1d�����O�n���҃�['��ͽR�<R{��ѡ=�����+vtJ����o��"X�DF24P>�[��-�_�5��H/��? jIxZm��&�qW�W�o�z �;L����{|9�O��V�nQ���I[ek�Un�k����t[��"��6{����o�P��Ѐ�0�;�30!�J����u��1��7\n%�|��Y9��=R����<�8��5��`$��$A~����%$���鰆FE�(�ߑ]9���\���@�E���nIr�ŞL	�@coYwO�#D<��B�[>s�r=�%�������$m�
��^�?�Y\���˺ٗ\��q+DH�Κs-�V)K�]�1��9����u�o��@���-tWZ7���p� 2��0���E���.[��
SG��T�X����(2��i�qD�4ĢH{6� ��
�ֻG� kЩ��BHS�������^�m�^�x*_��	��ʯG&�ʬ���ܓt%��E�����������؞����@&��&�^������9�;�Xc��i��T�뢀�>���:)�A�I�1QE�J��Z�ٗ�$���)�v��}�C�}J���qS@n2��43��Xi��8+�=]�qEW�VM���YlG>�د�u�7���x]:�D�'JQ��Ak�_cg��75ߛ�/��8�4�3k�p�xz����s��+rFmYk�e�)���?�Bv�D[��q�:Oq>Т��C���'�v������ɗs�`���.O.'L�P�i+�_���	L���/�j��x����5��%�U��$��c�p;��M˧V9h� M�x	�~��>�V���6a�j�>8�d�6�f�m�DH��;�г��+Is���{���F��p�{�+�M��Y*�V�O��l0@��6�~5H��Wʹ��j�~���=W��Z:������BY�t�u.��Bc�7UzTW�}���v|j��/��2��[���e�}#�ל�>���)�1�x #�e�Ab*$���Cw��<[@-��,:+�#����})��:��*A?-���`�Z[d���c�Q�"�T�j��?�O��٠���y�y$�Lu�s �xR��r��ֳj{��R�IGZ������ߛr{�!�D-E��¢������2�	�j�%�9�!b~%���Z�>�r�Dg�Fw%��+�nM��q�'�"�9�����$�����$����'���ǁ�*U����]������z8Ñ^���O��	M2����\;�]�mړJ�'j���%V��	4�*+�"��+�>�n����D8v��*�kp������P���!�t"{=1��$/\�!w�+R��d�<&v~��5�����[5~���
���$jr��O��Z�D,�����Cϒ9�:3d�����Ǽ�K����z�O�����]��z�^�O��%O٥h�0��O:�A�!�K�K+��7��i��Zݑ��z����v`�&؜%OZ���\	�|.rI���ʍ.)���A�<)������H�Î�3<�v?T��>�m�--��?4�\,��6����a�y6��sb%`#�H�r���>��?E,�UVj\b��Ѳ���)�p������S�����ۀwk�9�WI�/��᷻���诮�kJU�:��^#���>?�KJ��|H�p����<�<]���l@UtY-��>�sֽ��+<�=L����L� H���\DȘ1�B�z�!�N�{���ڙbzUvvp<Pc�3��ч1A����}�8鏣���L�͹V���?��!�ȧ<W�й���OO����R��O�VdŔ�0P��ac�SnY�O�ٔg>B��%�����ء�漖%�vbd#;����E�p���)���r��IZ�A��(�A��}ic����@fx�dG�]���y�C��6+�$���������^1/�z�b��u��jh�����~���M�..	�[���=��%s�	F���+�#z9���^��oZ5�qxf�ć� ���϶Ni���S�e�3�f:��'�㬉(�Z�::@ޯǛ<�{�pbL�p{��HZ�E,�EϢ����D�-��QN�"4e,�dN����7&�C"��2#ȚSAc���������4�.�I 5WHy+����� �L�ȟy��r��"���P�������!Ez�P	�H�e7X�)��gM�V+���OV��Z�[D�)�t�E(�}�HX5Q��ޯ��<e��@^�$N\p�twP�"��?GS>sH��7�&0+����oC�{gu�˥�P(��Q`��Cs&BB��{vW�dM�~�O@{E�/��_N���qz	Jwr>n�I�k���f��hi氒�$��cW�"�g�ًY�(32ݯ��_���*^�dv\��֮~���T�a̻⒉������J�Fc��׀�ɽ|go�L�v��r��77�5,�v@��q8 �hV��%����C.�a�n&�FR7#ӟ,�����:�:Y�����Z�#�5�F۔���s�ڌ|D�|r���V�r�V�5_Z=�Gn禦]��X��uj�m�n���v�[IV������s��o����.��k�O�J��գ�5�Rc��̞���Ih��4������i^���Q�vEz�|�p���1R�P�b�t��fn�>��lާ��Ӽ�e+���r)��hʐ�/��0��#�	O��Vl!�D4j�0�� �Sp"�^�Q�3?��� f����. ��B)��	�����y7��1�&~��N*��i�b�b���L��i����U�n�V?�V-�\%?*Emnt8��E6"U9�-a�,�G���{'~�!���/�E{��^	���TO�g3/�D�#������*4��ݐ��c1�;�蹥��&�������\����o����Nn�2��r��8��P�塁����}��e��HA	ͬ��TJ�s�:x�4��X,(�|(�ą4�J�(�ڻT=|�mc�_��e�_vd6?���'>!4	�
Fb�[��`�C��`h�W�ˢ��o��X��+Lvi�G�Z
���C���`<b{.�?���b�Ȃ�:GHTo���� �J��h����@Oߜ֟jYvq�ӪDy����O�K����m@�+�=b.K�����5����WW�G��#{�/"�X��AX/�
��v,O�y7�S&+�[Q.t�i�C��>�ީ驶�X;a�0>����	����r���Z,��/���:��4\�_���G�!������������mnc&I��G]�[�>{�;��3���GH4���͗��#h/O�J���(�7>-U��#�L?g�'T�J_�`���>��i����C{骽�̭}�;�?w;��7�/����_l�o6�R��qx��oGjP��Fw;�9&ǯ�5�&������������f QOf�-�]?�K��s�����ś�?���%�t�O֝|w6�֛�v>8���J�l��ϰ�%���uqܐ�DV���o���ĕ]�ٹ-�ͧ��aC��A�AZ)������W� �L��S����Y�����Rs�~N��A���)wK��MpQhK�;g�������?>f;��Z8�D�,���0��p�.�M���p&	�0�UY�nР���ncqʹ)�@
�v-V\]�][����:�Ż������"B�Ҧ�(���jE�*"E�M/�s��$E���^?�d.�<�\��{���1lw`v���V|�vR|��69������S��3�w)9��h�D	�D�I�N�q�@G�Eb�r����_|�;�t��b�`Eʩ�C�\(_d 6[v�N����AE�.s��@�oh�G�엜LP�Cs��`���X�Em���������P]����F5v��z�A����r W�@{� �����v#[o�"��@�ԭ%[��(d�3�Q�����+]z�G>mb2-h�q��=��i�G��PeX�鬻�h+"��� ��L)~���"�< Q���s�����N��V����g�5<���������ٔ���!� ��i�����k�\�G)�[K��ͺlX6�r����9��q.���aA��^|�0�6�����6Yp���m�iKIV�j�X����K�(��B�6�u��h�ؓ7��e�x�\�=����`+<�t�O�OG���K
K���L��"���@�(��QF��#ٮ����iC���>�-��,�}����l�n�%B*zF��+��.VW�EX�1�B��V>0n��4y 	P�'ZD乪�#$���M�J�,�ߕU���~s�N-^�y��D�S0^�R�j�ͺ�t��0�գ'4Q���=�N�	���4���d�\q9٫���z�C�@+��nK�̨�� �I�>�i��k>t��j�^��(���d�N 1��ʈq�]$ ��ጊ��?�������3�\�+�8:�����-����h� ؔ���<���d')����ߚ���+�5���2G<c0�G?n	3@~e�����xu�h3���spt
�D6����8
�3��l1U��-D4��[�"0c?8z)��cQ ��Աr��[.��F B�t"į:Xw5�j�Ѐ;;,X)��sR�=3��lc���C=���C�	1���Y���w�����~�9<��Ќ�������<;"��%�,j��$��>�`�əa�i?h���t�4e*���v��@Ҋ���DI������e��������7�(��S�.̶d�����*�ˠ(.�d>���,��yv�����\3s;3�{�(�b��c�y��N
'1|�Ҝ>�>Ni=��?-4am��_����+O�)��hd�՚�����l>XҐ�YY�2�|{:��zF�ڀ���;2��B�8�+_�/ �W�\���tpi�7�^$��13�&8�%�S3#Hg���X��s�|L����-��Z����g��h	�7�I��3� �fJ���Ft��n���3��Ơ̈u1Й7�BR
˾c+��z�����Z�i6 �3h�^AY�ό��'���㜭z�Xk������Ջ`p=5e3��� ��z6�i��������,du�d>�M$nG�!��,�6!^Dr����S�xF�&bJR���p�eO;j���"I�0Ђ�܅8��c���qD���wU����:J�Vm�H�m�@�%&���b_2�
>h��Ap��0�����u�se�Htu�P��<|�r��� ��MJk=U�f��߶��9�B��O�2�%�����SstI�W]�!��`�]��t%	���3�rS�ʹ�3''0^��a��Z���������ɂ��
��n�.����P���6H���3����ٰ�j��Ea:�ԛ���u0���~����1����%Dx��3��5zwn�P.��Y��k֞O �|��������6���?���8�F_�E�����D�zQ2��Y��uf�1\�Fi4�
���$�!H�h��N�h�a����ụv�=�"�"�yz8Y�Ƒ{�"}�ԣ�����r�~v�Q`^�T:�p�}.�^���U�?���e͋깿2�,�N�%�w�0 �'Q�#Qh8�˸����،9�v!>匁�A�Xkh!��?�E]$"h-��U�@������bwb���gè<���R��+ER�����>~�.��&"���c��6�0^�}���u�=��yd>��[��E4��Ä��X�X)�F[I�h���� %����ËV�ŤT]��+r�/����p_p�����QV����4��qZ-(��q��@�(�|�Z�E{�k��q�ݚ_76b
��tË�NR�?�$U^��If�[Ш:�'�)��td��S')����;x��	f6]����3��N��\^Hg����|s5yr�A��Ī��qFK&�G�;�Ư)y�^,���FHy������s��Vw$]z�~�-�N1Gu{��T�ڊ�&omF����B��(l�Y��g����OF��K�����U�P����yf�GD��D�SQ�g�?8����⻵\��2"S�]_W}MH�o	��-�A�昕s�N������W|�m6K���'`5(O���T�D�������`���P)3�����V�б1|��0�����p8��`��ґ�n�L�:)�V{��|��7����ײ��%gqL�����'s@��K��`�8ZA̽�9�4J�>��8��tP����$�Q�C��u�<C�R�����\���l孷�z�/����c��*BK��k����r�s�Y�ȅ��/��Sa/>�0ʹ��Nq�����4hc���KRU���NĜn�@$����{c��Y*�۹nX����E���ǖ��+�3l�3c?�Z����Շ� I��XR�9���1���h�����)�dU� ��o&ߋ��wZ*]G����y`;��0؊�	�0y�: ��V�'ϭC_�ݫ�(\
�o��=P�S]�%	��r�A��῰.�s�5̓�߷<���Kp�9X���ܚx-�U��o��ng�Ҕ�������NY8>?�]�;
Cy(�ʗ��xP�����?9'�d�ba�K��ÆD(����?�C��L޽!|��x�������%��|u���O���tZZ*��E4���rb%Di�]GJL�f��˵Lקu���?�@�JŰz�gz�
�J���/�qh=S��M��_���2X��fL|m�J�]>�: Ј�h(p���DO����3X�"���8�UW9A�:;��o�ڞ�Qg9��q��`\S�0��P�}�]�ŕg1�x����ی9�T�s+E�G�ii�e�f�,��a��7��`�~��)�-�X�v.��G^�S7R�-=�(x��t��t��(�<D9��!j�\�H�_-OK�:{��!���Q��(��U��v�u��uȃr�07*���$��+�Na#*���^����r�,�/,�a5�A^|�E��:�p��%��&h��1�LDć�)Q#�KE�
�<s�T�P��I�n�\0�:��$h�'U�=�C٨��|�l�HT���4��Q���K�'�=<�|R�$ݢ�#L��	�9~%����eOv���`�����e�,�q����U�ܲ���`a>�2�aa�V��'�\��?��y�QM;5�
hu�@]'��(��"('�����j����q��wd�_v��nM�ѿ?��Y�}��>Q~��YgB[�C֘`)�b�B�-�g��RDyp�������6j������F��	�Nɟ���_P�<>%�e5��`��&4�G�A�.��	WwE�U���dZ�8�K�ލF�0⪃��%	���|b1����]���q�͟ �E�=-��Q�yg����R�7�rѿ�h���K��a�>�И��V�Gj�;֬�ڝ��d��C����%��4tb���1���6�z��hQ.Nc-�[�-g�[6�QQ*-���nx���=)�!�3L���y�\V���j��8�nC.�Ҫ@h�N6���4v
�	�,���V%l���/�#�6��u�jF<���0�B�:^��w�0�����]���N�yR[�?p	�$cZ��w4�����&��ޮ�tQ�� �6<���Mq��9b��wX�&��v%9�-�H�lU^y9�H`}+�}� �h �����id7C���#Ve��n*�c��:�cXf��	ig��jch.廡}���D4�o�ę5i�ה)�G�R�~� '~m����6#ȴ:g
�9��v_H����GF�m�Fx8�%*�h'�V/EX�V�^�7�$��0��^��缋v
�0�$!�1�@��
'�����vc� ���C��e�B����be��A�b>��>ܞqw����_}pɄ�+G�3�:>P6
�rPu�<�_�bA�?�1���
ہ�f�5���1������Z���h間�����Y���N�9~m���|`�D$�U�&#��ň���=��%���|�3�
t�g5�b���ـH�J﷏�z��|��g�_w����J��|>T���\�!��S9x�1��R,_�R}�菴_��W,���θ��`-�/RŲvF��e���ٝB60�T�P�6x��I�M`%վ���e��`,I�#��Vf{�A�?F�gY5�.F��>㽐<�i�I�oP_ٌH��l|z%w��e�L����@����.����k�7Ⱦn�"K#TэX��#��z3�M�rlC��L��l!���Uݾ�����醻	��)me[V�PAh��t� w^Y�D��a�DP!3Si3K���bN.	v����}���D���>�M�e?���960j�O�=�xMl�|�m�����TP-��U��f`��>P�~q���r~��J:��_=�
�\,E`!�'�;�zl͡_���o
��.�Qb��2�F��	���ʔ]�k(�.j�!"-��BЍ,�w�?T�b��AA�X  Ɂ2�YL�%Ŕ�����O���V09�_�ɯ��.O���\@iN���a�����b:�'"Ȗ���]?�X��G��n�� �C+��Z��?�̂e�Z���=
�vXG��/[t_y`E7s�!�����&���q��&H�1"�+a}�4���>��P��}��|f���5ސ/6X�M����d��6���(uV�7�A�=��j����ޤ��b!����{`��.0�d��`�s's�'�8�kTZZ���$�-�y��i7�mM@@.	Z��1�WA6s��V��6��Z3�(��lǅ�.�_�=��m���h�n�9��b�I�S�����<�p����=-d�b�Ɛu�7��n�\��/�Hٜu����e_��i�b�PW��{ܞ�R�W_3��h�q\q�zu)�5��x�3	͉�������c�ڃ?1_+9n�f�pX�ҽ����{�E<�����}���-�bF���\-��s��k�"4.�>.�>.2�̪D���ˍ�|m�Mz�<��B&o�8��aW1'PG��@��7�1���^���j}3.���2�C���L���%)Շ���4+��	��Əhg�w������o�Ź�#K���7��Q�R���S�l�]Ӕ_>����k0�7Q(M͔tb���a���N�p��]���m��L�Ep�W�3�;Ȣ�j�,j	h�����1��>�H^��	'�YD�lC9/_��b=�Ƹ�,��N�^�/�I_75�is�^O����ѷ�lp���R;w�"�ʛa�p��b��ŋ7�py\�F �O������v{e
��H��n�M�V�^<hD��`*��<���W͂��w�Dv7#���D��2�A>�d(�h���
u��#�n�;PM��6&&��-}��%�Q�"}߮^�@b�]݉(��Z{r�%���Ǻ$	��Ro�j����%<pb:���S�ԇ�h�+��(�zꂍl����8�)��P9vu�?I�^��Xt������?���T�*� �t�.��NV��	���SX�j����B2\�9Aڦ{�����O�]�*����&���O~��9��e�V��D^n!E̓a	���@p��a�O�-(G|;D~K'�Ǒ.���.�,�/���X�i��Ï8ґ���_x2�v���tؙ2~b#��''���~������d���@���wK��M6 ����iK	2P �>ړ��;������G/T�'��eN��bN��h�jT�-��]bB�
�?�XN�<(P	����-8,�-��p��qL�
|�飤�qX| �HqP[Ncܛ�n��\���������ԳѲ|�vlei��T�%����*��o��3�҈��%�rƻ�����N��/HQ�Vڟ��k��k������x\_�is�@Ş����u�o/�U"_+P*��ˍTD�Y0�r�Ư4�z�s������ ?�����K��U�aUi)@�a�b�u���bQW
���Se�bq�U�������(��f	��6��*/��ق?<H,�ǃD��)r1�ER1�2k���D�D���d!M䕪���j�
�űC��B��y�=��ŗ�����,<�x�EZZ��|�ꐏ�IQ�z#U��^V�ƞz��W*�V�Q�n4��y{wg���h���zvSJݙd��*C>���ޮ��EU�E�+�2b�	��Hߥ���_,�W
1e��ױ_7��lo�.{�l���X���:���'c��լ.�e
]��:�(/SݛY>��J3�Yj��H!Üd����W��� ����\��4�����8�7��|n�\�ˢф����ͭ�h;߬�w�����c��n�|��@������U�f�H/����H	��@Э�{��Ռ�Bb�� t�3vV�{� �6��~�>�e^4P�<�n�^�;Ы�p�0t[6�lϛq�(}��UZ��qe�ƸN��,�H
�E�ѳA�()�r�9�<Q�;��ap%�����}zJ�S@�<��$�"gu�� �����r����=D	K��MJ4��h>�~?eI�ۈ?R�t�8�|ZKo�P�ƀ#����a#�2��Z�7�»Ђ��cEV�<z�"_Z]W�BRp�� �x��!}�_p�HV���ѱ\����"������k��v�c)�C�������xQ�z�^���tɖ���+���]+F[����񧊂?f��N�Ɓ�^`��k?r�aeu^���v�q(�n2��R��'�1M��WX�4^�nteB)+i_��^P��$F�����ЕW "�3��!(���ҡ����C&�.�l�bG/� �����@4�����=��| 1�E9-*�P������	KT�M�,C��@�,֭�U/!�Nl0��}���G��G�9b��T��Ղ�L;.1��p��\�F��e%E�ǘ�F�_���b�a�+,���o�� *5h~m_��߿ߙ0u�|C\Tɟ�>�">9m�@�5F~�Tis�p�z��H{�b��,��	R��E�7�70z����Ot��;Q�[�ǚ����L_ōH���:F';����޿'20�w=�x�<���2��N���5�4���胴��Җ0�����K�A��h���1��s��T���}�r�;���!Q-��#�|�.�L�z>�P������A�N14��_YMR�����waS��"����pN9�n\�Z1�3)�=tA�4�t�Yu�s��d_K#�3�.�����7rx�T�c��t$5�I�9;��Ncq�3!H^���n�SQ_x1ڟzv�%9�H\c�m�&o�J��ޏ�L�J�S����A��M��u��]��5�48���Q�����:g"�9���ݖ��Sy�t�FIK�#_��m����w�Ǝ�}W�H��VZ1��5�b<3z`��p�+¤c�X��ˏ$��;���I�63�Ԃ�&�QPT4"d�n�������@I� J(�O�c�p����3D3I6U#�l	��nʐа�G�4"��w��D�	&��׽�ە<,�hv�<2?��I�t��ݔ3�0�:�S�Wr| �<S"�Z�|��p1n�D����r�H�|�8�΂��o>��+}&J�
��G����F3cM&��QB7)?��SQ�/,�A���ʢ�#���a�xo&SH~쓺)�t��6Qy�x%#�%�'$J��󍕆�����RnװN��HiW&��]�y���(�F��|	�N?����V؛r�=a�8\��^z��� �0�0��m	Ҋ*�ٿ�M	3}��e�;q� y*ϖ\ �VW<O����D�˨'���Э��	U�-Q-����#���c���p\�ˎ��M#\,3��b_��}���{>��gϴ �<]��!���?[�Jڙ���e�����}m6�01j��+:(��X.l��<�����z��7	|����^-�F�����O q�8g~��i%�܈`�7L�}f6©!�����(յ�@���z�1+��ys�����N��8.4���sK��g5	,K#�ٻ{5����[i)�j�^�����%��a��I�R��kwx��	2C�a���0�k�;,��Yj�<�6����`#��Ą�u;	�R�J������w� c5i���w�>}X:9jM�L���.B���͡� �[xO���Sac�Pq>�0 Β��|U)?�Kdہe��(�ŗ����_�w9��+�u
d�����=h�]��X$_���52��ձ��n?;���m>xu��B�f�ؙ����A��T�藰�O�$H��yd@MLӜ�^7�2b|d57�\��w�x��8˫s��!�UNЂ�q=��ј���,m��O��s�DV&�e@�\D�%��d�M6q1����E>����]���B���Pmj��$"�ْ����-��,���Kf.�x�ff6ˁ���A6!X�e8i'�X�o�FD������6l/�	��r<����$���bl8�է��B��N%�NZ�&��r�P�Y��K�FɝW?�} �Z���B�>8��zdٲ=&���{�I���g�m�f�؁'�z.=�诟eƮ�0�_y!�L� �Կ���5
��g���p��F��n��e��T�W��nV��ghT_ٞDd- ���1�˓�C�0XQx��|v5�?�'�����lt ⩾�Ѯ��r��d �-_ K��,�����W���m�t1,�{{4)�^��8M�1�|�{�5AL���cps�۟��ʳ�2߁�����a�d�Y+I�)����7���/��M��� �Ǉ�7 ��^h���'����W������H�{A�b�2�}���|!%*>�������F�Ѻyߐ愚�!�]�)5噓�<�-�v�6��~{���s��a��� Z��߳����@xT���5��K���Tm=Z���aG۬�h���M	�l��d�%V�Vi('gH�[xw}
��ߍ]�3��O��kף\N�(�G
c�pj�����{l�zvX�1Ĝ,=�c=!�(��x�DB:�����&[��LZ*&�~���m�o{	�u���W�,	{���`J��717j�Z7T�o�w��1=�ō���O�)��z�v���a�ޭx���G.��9Q4�Z)ǥG����()���5>o�^����0cIp��O�t��"eW>�z��n=�E�I*ms
o�]t� #�I���Eʺg���o�t�o����ݸ?��f��6=� m�G����}(�O�K/ȹ��q���9�+�:���V��/F���I^�`���k?_W���n����8���|�8��4j�D��r�q�I]�YP$f-R=_��L��{q��]�bS^t1��@�7Up��;�
5�M���r�~�ǈ11���?w3�N���sm�zM�+����v*C�[�Qpq2��{�L�ɰH�`ٔy������g����E=�k���4�oӕ�Je�4�R�}�����呋2e�$�|�XĬf�kp��׷!��#2�1;A�.��L^�}�b\�xx|��%���d�G���z��CcSX&��iz��2�m�E�"�%���KP��{��'Lo�"�;�ˀ�~>�YR�)7�ua�d���I��ۺ6'�?/������ʓ�&$/>�.�L^t$/�..�>�n�{FmM�c�{���~Z�5���9y���hg�8r[����E��.y�cQ�b{/�u�5��#L����8;a%E�v#0�|�I�E�گ�s�>��R������^W}ſ��|�Ke�>î<r_\�W4��>y0����^�Ȗ����fb@(�1�m���P
7��"g��B�2��K��T'��U'�WY�v���ґmf��A�s:�u����Mg±R+�i�}����y���{)"3��Nv�d�*(���i/��Hy���"��Hr�S������@�
��*]|\��46=4��i���Q��?�jo)�R�(�e$�2V��ϴ�I�g�����u���>`6!7L�ՁQ 0,|Wr��~,ʳAu��+��E�(C��-A�E�(w�;}�[*ᗍ�q͞,!]+N�_٢�.������:�{�"x6�������[�"�ko�(=��[��D�Npv�w{���+bj��R(����sꋿ���$^�o|����+������72Dכiǩʗ�A<<��;!��Di�:'Jd+z��\LE�b�����&�������>��8�a�O��^����{k�[�R�`�#�W���78C�Owi�g�A��~�
{.�;3�F[�T������6��GQP-�cp�\�{�.HU%䝓f�W����#�������;���p�07i�f���z�y/��":=�f���F�."G3���Oh��;~���� �x�f�^�B�{�p�n�2��Ǝ(�v;�{%��dh(<:M�X���Ѯ��_"x��H����\�����F=�!:]j���~�Q�M'/���ck	��vN�#߷+^�1�*v����À;�ANqQ��fTLCF5x�*���Rʏ�Hx�/�`L�gr~��<Y}竔��dcKw�p���E���t����5��\��r�E��V�p-E�U|#�(To�M��XA��ש_��ap�JA���O��<��_~%�SRkj����!�c��%�����)���pkv/hG_�'6y�ܣ�p��)�ά��V�º_1޼o5��%ht��o��e4���&=NBl����o�?T�H�c���ˇq<�ci�֤�ǋ%�؞()���pS��E�-p�@N�btuǀ��:.��l;�\�+��y��@�%W	������1�������+p����W��.�fp�R���W�Xz�*���^�31T��`D=߇��@�h�y!�XD5�V>���������&�@)_;u:�w�Y	L�Y9a���P@�Nͬl �
]F�1�4��'��y��a���)S��tk��#�u��.	R`l��^{�հ���6��JjQ��`�':`�chU��5t�x�(��%�y�-��e�'������H���}�í,û��ኼg�V3!�3�m��-Ɗ��ՙHy��	�:���W{�9�����~o8 �@��:a�m����P�sp��͇�7�<�$i��$u,aA�0�5�ȡnN�?6<�w�:�9��0�����J� ��r-�X�����tt�����E�~t��Ey�~T�A�-JvuH:�$�6~LG��;>&=c��glDO�̨���a�i�5n���B�ռ4�$����ݚq���
��Yu����7-d��Yz
��W�$�T��e�����'}Ai�wCYb��R�P&�0��\��i�WVF��i\��]У��j6��'�Q�h�
�Z5K�`\A�fZ�`Z���q������Y���L0�S��.���U_wb�GG1=F2�BiO�y�|��T��CD���_�M{�G�
�c^��>�`�F ���nM+�r��^ˌ��?߬��������tӳ�5��.9���b>Phư�#��1��gn0�����^���7�Z�)3
���K1uR����@��7�m-mЭp{5���
3-z��7�kX�-X>���V>p�p�/���!��9���Y�vy���@�g,>��ϒm�H�PwU�ӌ�wi�)K/���ӱ�9��@��Ҩ���]���Su�h���}i(��,;H0@N-:�ٹ� �h�M�+�OÆ��@�q%��F ?,��U�g@z�N�A��-�E\"xC#�s��ªx�c���.Mǀ�9?` c��O�5��u(P4�<�	�S�E#�P4��ۀ���SN׶ۺ�F�VC;»O�@�ҷKwS�b���Z��~`b!���a����m��$ ad�0Yz������^iU�\ܪ����ZU�1%�W��� �l�+ȹW�wF�f~�Xb����}�H�;i�#.�R���ˈ$�ud����t�e�����׾���	u瀢�u�-��ԦWK��5��ӄUd�3b4N1J����r�ȽYZ~��<�6��rYQ܄�Y�F�"t{��{�(b�L��+ �cv�&$�c��w��f?.�!Km���F�Y��#�c$R��@"�c��-��Ei��h`؆U��P�u٩�~>R.q��A��L���0�Ԛ�� ��h/q�Ԭ{D����Ǭ`�@xf7"kV{�4i��RüC�Qo-�X��0�<��*�[[(���֔�^.����L�;S5OL�f�1��[���/
� ;R&�Xp3֖��V'5%ڈ��y5!�>16�� N��K��������ۙ5�Yu�fL�VR���'5C�Q�O2F�lÉ6RN-��{�\;�����h��"��Oe��z��"m/Q��ܔ�D,u���s�S�_�(E�]�Ror3
�YM^���|�(�齱\���p�|
��/o�<��"��rR��jZR�j���F���Ed]��2-��ڟ��6�7)�{t���zx�L�a����B�G\��M�G�7�o@���OV�z"�Q�Y�Rx��+a�"�A=�(�5��OMc<ԺȞ^��Z��z��t��1��!$�rrS<����"m0ei&ʫ��Ŷ�F9[Vl'�9��)o��W��i�������]�����:��^-y��RF2�S�W���r&H��aAo�cF
�Պ�/e/�O�&���|�3�ơ@���~�Ym	�@Σ�5]�����O����0�\�u��R��('W����k�����L��� �ou�������MU�0AԾê���B\���S����tY[)�w�c�჉���С����U7�H1qK"gH�����ŮN�f�-�A;I��b	#;�K���ٖ%��:U�?�'00y`�ʥ�q׫��#�]�G��u�"�3��&�$���'5)�I���N1C��gi2�t��Z|/S��R~�(O]z�O�F�(�.R��f��@�1$!y�mlPj��H!�?�ٗ��s,��%�ƒ���,I@�W�/!+��
 V��ѶQ~S'bQz�g���5QE�~�0��>�fPp�F��ȡ^t�P�����Pv}ʂ�)9,�/o7�ʼP��/����#�4mOB�| ǜ��*������.����X��(~x�E|�7	�6ng«QF�����]Gz5k�?�<�T/E�������Md.Jy?��=/&3v�����ה�S�@���BF�)VX�H�^�'�] �c��[8}o��c<�".��R>)�U�wr�]B��E8��r�%13��H���[<�V���b 6��y��'��ѭ%��Gn� �Ā�)#���mqv:n�gx�_�0��B��X�����)x�Y��{�W��G�M)ك�$�=����JS��U��]}H��g�Q�w���5Lo��Rp Q-\��̔)P>��7qR���c�|w��c�M����V֤�7)�R�jR�<DE�W�h�	VL��Ž�����r�V�����ش����l"���l�o�NR�e�O�T[�L嫝l�G_fl棏�&��/�2�����9%��X�����N�r|���}�;8�s��f��������~��aW
ٻ�RC����<#L�۲C#���6��4�b:�	!�Ш�ÙQ���c���ya��r<�#�L��v�*��Qbj�=��,z�	V�:$�_��Z"NXЊ�Ջ�gnz�	��u�|�$�rB����o�)6l�7V���&��ɮ\�5�����?���J��5���i��,�4�O��*Y���X����'�gHO|/E���	a}�S�3�1�L��H�ف��8������[?!��j���	yA(���Y���� .����*������x1x��DmX.LG(�@m̼��e��F�_�e����i��1�q�ΫLL�^D����[�����:�Ŕ����
�e����@V�[d$�#V���y8�ژ�γ�ȗ�l���y��,�n�	����&�ʏ���	V��G�k��'݆2sa�nG6���������P�X�>0{ jk�Q� ���(������� ��$Q��좲���F1��#�[�-�r7$r�+�d�ݪ_����\1�'�kAu�pӅ��+Zp��dId���p���j���<͆}��&���&�����[:���pʄX>Pq�㶚��*��'��+���6�\i5��l��)�����w�V��5�8];�+�_�B2̨�<�|�pLa)�l�F	�\���s>�c0%g�YL�V?��Z�I��:C�<v���Z��Ijj�D��e��I:yv�'.�9󳎵O�/��ָ�F��N���\�~�OD�;d�Z:�ϋ�ğ'}���.��t��a ��C=R�GY�H\���w�8V~�)?�l�|>X>�x|%l�"z.l�w�������8|�����3�U���A���3�U$���c�Ɉ��SD�г�3�tC	�>>�i9�οb��D��Ҡ<Ba�C o�G�t,�j̪��P�# �,�����.-�w�O��-3F]yBDjrP9q
 ��Z��)3�:�G����!E~�l�����s�#��Q	�O�� �K���;(���01mtj��������QN�}�lpW��������)gb���Ç���I���
���{DbK���P �]�A0���T�_(E��Sm������6>����Pa��I���y�M�7�Z��<�Yihxa�Ŏ�rZ�W%�>�k`�ʺ	q�_�����z)�-���'_ /�ǁp�}��2U�T��a�7濳��I\��8�	�}h3%d�0�F���f��)�eF�n�I;�u1�+ϱ�Y�>U�V����ɛ�>��y�!��>��P��K�;���SӁ��rY����&����<�� �K�B,��j\	B�+1��������|h*
�Se����GtXX�2c#3���H)ʏ2F�Z�n2�P߈��}�%����.m�枩s|~�:������*�TҎ��)h�5,��ܸ�짪M F�}��N��֕��b�+�B�6��	"G-�r:�0Ɣ�˽rZ�x��6W��;��]� �������4�;���"N���\��^Gg��Jo��{<K�#vepbe+����p3�\P��Sj�1߮���Q,�>,rQ�0��Yi1m�ϼ�ѣm]6�3)o_�<��#]�*'o�1��N4R�՛;����>���	V|tɮz�$�)����n�0� ����Iq�m���.�w����4�	��۟ �u���8Ɵ�'���S2�q����׍�afu0!��@�%�d�7�hz���na������҇@��J_����}l�W�&�����y.��Ul������o8�+�WO�4�����k�^|9\2{By��t7�A�N�&��#��7cz����9�k��Cé�1t��&���@�E��Qެp";(����,��{Q��� FYYW��:�!��EW'�sP�=�*�a�����!�����Yf榿�r|P ���и4�^ٙ����7+v奂�t1�)���=���<ߘ��<���O�|_�q�0��m��t���)PƧ�:M0Cs���)�Ϯ��K��NI^/��J�%H|��n�bh�z\H�5�3�r���_�[�ۘ��mp /)&��bA�o&lih���(m�t���;݊�����(��� �����S��=�� �#��:�N}��m;k���"������޳�`ŉ��0��BkQ;4�����S�B�j�0q����(���jYۆ�}�oD�����v��მ�H�%���n��=�ao��%t�7������᳋�S6��"B?b>�}��Q�`�N�>#qL�,��3ɓ�E���r B,�{�5,�;&݂�4A�)�U��Z�,��У�w�At�7�oW��H��L��0������^�uֹ� l&�0?��,v��v�Yyb�C�9b��׎�k�\䰍k�ǝ��ҋ�%��9�4�ҁ�c�4
����Q�H�|�}�h����+V��Nw��[)��
�H���R���e�x�-ui���5�h�Z@M/� bX��K��6�^�ݤ~3�/�1�V[�2}~V�r�F�*�`?�R���;�[����]��ĩ�p��Ȑ���J�͆D'�tۙ.Rb�pQ1=��`]�\ݸjLJe،)�/�W��9]L_[���!x}�z#�ԫ��M3��?��ʀ�,J��{0�q��]X�dy����:�_@�� �׻El��J�VfÒ����;y/�k�2Qi�����Z~O��+�~���f9&9�����	�x
�ۄrG�F&�1���y1����bZc����wr�A�b�к����{�>�Bz�G�����{'� ��N�����<Tq�����0���-�o���6���hYKx�	��|m!�`���t.
��\3-;ƍ3�_�;��n}(��F��r�}T��kXyڞ1��g}>�r�Q8y��%/y�I���;��M��M��?~�ۤ�/|��(��I^��U���(��;xZ������g���-�~��|~��cc1��	JE�����i��s}x+���2�?�>��.�q!�=��QO
Ѧ��?p���y�yF�n�;�ԎW\�C��[y��6��+��+��m���Mnw�p�K�l?�����<�#��={l �� ��c�HH3��fߣ�}Q��H��ߗ�u���������\L2v��>��/���Ҕ��|��b@��B�Nj�K��4ʒz+v8�-?��_����(V�A4�U�@1�03��l*K��S'n�G��u
���RA�����*Jꭄ2����'�A{���� �����R�;(�����p��%��������� q|�f�J>�:��S3�ƭ��|�5dy���M�y�>J�{ǉ���YI|/�c��!� ^r'�c��գZ�J�˘��	��uFڇ��Ú�|�L*�sP�pS�2��i_t�	�/��f%	���~�:F��B��H�`0�F����7��ּ��Z-㝝�3t>/�)R���,:Gx�x��]?��Q⟳�́Q�=~b��i�ϩ8�����rG&���
�|�GRx�r׍qr!��^I��?�2�4s9�u{S8���Sxf��Պ���B�ӮN~��>�[�*h�m�S_Nce8����WƲ]����4��{���������.	J�	L��a������i;��B�"�V1��\UHĜ[P~��֓�9��,��([� �d�ЀL!*�p��)iQQkc�_�w�����O���L����?�a�,o�AI�3|�#���څ���dfxK��E#�Ҋz�Mߙhs-�'�I�B��� c,�ʾ�v�{EK^�?n�I%p��"��f��]S9�]�hd��+K�g�����C��0�}S�:QJ�7U���g�	�1���'�Dy�I���$��w�O�o�N�, ��k;��C��d~kf(��
�m���:~�Ց{�^5��#H
��*o���Z:�.��W�O�3�fbz��>R0�°�=�M��]���>EOA�v��$kMؿ���W�a+��L���X��F �Y�zl�r�ңK}T��ف\<��yDK�d�p��i)�*��5��/wd��82�a���ږ����C��Fw�A�� ��������0��!�u/y�9ηDx�d�~w�v����U�0���{-d��5�d�'!P�
�Xy��W��X�=bi��+Z��;L�G�҉�Вz^����b����r�'䂫�^�.8׀�I�<�@bDw�r�����1���o���&;B�p�O�^��Q珙�	Woa���į�[#���Wؙ�'��ņ)�M���Wr���	㗺∎0{u)ƺ�ߥ��K۩KS2�5�ua��c�D��>�)%0�ḫ��X~'�>�4zP�}^wB��?�l��=�Ē7��RJ�s�Y�#k������,��yW?8�Tq>��{��P^���^�!o0�DCN��?@Z��G����'^�2�EɊ���q?��ʃ��@.��|� ��O7KA�'b$I������O}����$�(����Vo�a�Y��!�u� i~�1/�p�����X�z���r�\T�Z���r�k�)���m�m�C�N(�>����|���svPn����Y����v��h���c\�2��#}d���@��5�b!��Ei�(�6�L�#b��,�v1�*�Ԃ?��&Z*�1 j�!+\�&�d�-0�W_4�jʗ�Y��R,5_�I�e��yV ���j����9x&�&[��x&T�s\�W�
�?n�WFQ��L3h�f�5]��)��Ӊw
| 3���Jq(2u�%B��#��W�Oꄲ���}�`b ��Q�$#Z�Ѕ�o�u��߸�����S��G��A����pb`+
�hݟ�1�:�� �0�/��ש�`C��\�;q��}�V?�>�;~�83[�H�:������Y{���ߕ�s:�C5��A�'R�H��>W��{0Ga�|i?e�z<���vO��˯�}�P����]5�D��A��k�(W�@#���P��$z�͇�@I���
���>�c����K�wn�)]�P�\̯��|��_yy/�	��z'���7��0ō1��%����S3�?
]�08|�| �>�V�V��mů�����=�&#!��.7�\Q�ȷӝX�Z���A�*>��*)����o�ׯ	Y��d	���A��'�*�������WOa+2���Q���Ȃ^�/����)�rH�z{_�������·63EX�J�>���O��'���	����;�>XL$:��������;�<-O�����̖8�4,Y��N�q+-\>x_/��������6\�G�	�:ΨY��E�č!�s(~e���%�}���ӽ��r|��"���a�����?�at�%�Ix��e�
�2�b�\K�Ö`b�+sY�a\ظ��_��p$i3XM�Ʃ�zpU�����$��_fX'�Q�ɫJ���UWb<��?�Ge��҇b��t1�J���7��7#����\����7�f�2�
�ک:nڑ����T��1� Y��a8��f�#��T�zR|�|���z������o�e���-�L�^`AWIw��{Qt�R��'����(�-:_p��C�Y8�_.G�J���IQ�,a���Oa�t&R~�����yě��5^��k,.w�K���U�9�Ԑ�6[�'�ۜ�%F�@��m�#8�j�����5�#)_T~P���#Oqb{���� $[��u��E�z���>���6�GpL�M�L^�����ŕ�&/�V�b�{�|����󁿓|�	����X�+�5?���ܕ9��M�){*1���������0+��4�S����1�+}F�h��{|R��rK�<��1��46�4j� ��bh�c�,&t��.���Y�듾���WA��l�z)�_���O�"�i�*gü�̳��z�����vL�
@#>�[}��~�r�;��'z4�u�]������z��M��?'��>��D7�ʋ	[[���1�X� ]��zN��\�p*uE�6��� �^E�>�=�C�G�f�3�.*,�*?�b6%/�2T�C�L�"�-��� ƴ
�X�j�H�'�� 	6oh*�^��kHw�^y��t8~-��B%-�'�j�c�]@���`��dP�;3T�1h@��$�K�ѣf���'�~�F�Ԋ���!Z�Zro]�%I�+}J�������Wn��5uR������,X�(�TrP�ΰ�~���g��3vN-1֋a��]Y�����dM	�A�5=Si)�����;��d;���*���p��3��.A)3E�#*���(�W��)6�������ca���v� e�؏�"Oy���ũ���8(�:��7G)���siƑ���Bo�K� /b���N�4/R^<���צ%(X���2.	�D�%��P�C�<�\Y!������g#�^P��H������!�HڀF�)d$��@��OAo�R(wp��"���X�OP?����?�s�%j�G�ϗv�I���y6/��(pџ��ǈ��Zc�=�{,���))�kAy�q⎩8�`�I#
�����<�d���*V�m���Oo$�U����s
l��x�1'��<z�����z������r�H���?i�z�k�\,�>� ��m����	�%���q`��q�.�/5�W@������?�%���c��%Z"�m�YC4ioM�%�e�͸֯3�
F3`Ƥ37��EyF��kۜٳg�B��|��"D:/�������.���3\b<�m����N^z��T��u)⧌�~O��jR��%s��j�wߑ[C�<���P3���U��)���g��⠶֧��=yN�d�O�?�Gퟡ�#���j���k8�^�<����dkav𴣅��hcX&�u�f�R�p �!J���*�X���ŠX8!�UvS�h���~Ƈ��e���Ĝ�d�=�R�p�o�>����B���\����(��f�"3s�S�%Md�"���:�3��_%s)�1WN%� �x
Z�[u�n�Y�M���r\�r\b�׃lR�Zr���A�K���������*t9!�.�r��s4Nr�������q}��Sbh�r14���l~�;���.�I,Y]��)�kQ�8�N# G��k�c�G����&���٤��9��J^򠛂�F�=��i�0�f-D��	���1�|I��X�[�(k5N��W���=-Z������Rx�}�1�8t8V���̗Bى"[&�HnlT���f=8��R���ү�Z��|,b�s,��:�Q�������L�0�g���kR� }�"0���3��W_���x��&OMG���JF�Y��_ʹ^R�ܴ�u{,w4y!r�(��0������	�����L����%y�ة�4�ͮ�.�WK�p�hH����P�g��X�*F3y����]_�{Qc��	#�d\0�x.��K?0f7���������*� �
��2-�x~VS�8c��J05�F���A������� �n2�'㒉���Ņ�����ύzBn[�wu��^4v��#|�p�9W�C��g*߁�'��B�Q�?�z4��u�fB|(d*��YǄw��(Bz\�����91�>��Y}&ۭ��S�/.����U��p�X���ͧ[=\��C>ԅ����F
%C�aC~R�M9B��g{sF;*^����"�o��DM��%v�&��8��u��kk�lWMjBZ�mw��i�v�A۝mw2�..ۅ�������8�kC�1J:�M���7�:�S�ۭ;�W�d�MIG��4��.�I��5$�8Mִ�J�7��;�٠�� ���z�@Tάۆjjd��4c�ۘ���N�!���kA�����@�LL�J'w�$Sr^b;"b;ϩ/T�f��83�&�S����Գ�E��~m(��������L���1�������bi>9g!ǕZ.������-!.�ꁂ�^$|��3yV�>�X�_-���z+�ŷ�q��W����Ls@@{�[1_i^�1�S�A�|�i����
������s|�o(���/+��`H{�ziƀ���(y�`	詰�F���m��""+L������&S�yL��p��;�,-�5�׆�Z����e�4����Ya��0#QU�÷�#I_��w;2|�qe�H�wM'D*t��w�kf��K��&�ރ�A,X���%�Q���Un"�n�|�|W����RD��!���h�NHn�"��I �ł������� ������?-��"�{�G#�aay���b�����Dd;Jam4/�H�Xa�t�ŋC��Nv��Ǭ��IY�8V�(�-�e�{�[gY�Y��\��.ٺ�K����z6�	�"{�#[�A8�w\�X�~!�-G� |��+V��R�zXhu jbj�5�������%��(u0��B�hE=�"'Ƀ�t�A��Q)�k����Cr6B׋��W�?���Wp$}�a���~�ɘ�R�?l�G�W#�+e�|���&�K�&����1_Sc�k2�(���J:�?�A���o`��Y��Z�q�I���0�'�ρ�@�EafCFE�����7�o{�gƧ�4�݃g�������Δl�]��|A#t_��𸚁ow=4/�$�F��"����?ԓ��5l��W�����~]����(zݒK(�N��Pҩ|�#�%��Gǀ�N�B�Aax�f��m
':/u}�6��f?��s�ek*���
�w���}	xT���,	��h܃F4QԌD̄�0���� F�JeF�@�Ό��2�,m�����Vm0�$Apa�" .�"w�$$���˹wn���>O%s�s�y�{�}qIY�?qC��7�@p�O�2b�ݟ�un��]�c�1���]u���<b���h��ฎF���'��!��Kϋ[��}���ch�K�W7�-�}�@�����E���N��������������?3�i:!�}�с�&g	���l�4���[Z� �����|� ���ӛn9�"���ˢ����*KDX6����$�;�^eIPN+�q�RM##`����&�5��M�l���Mcc�Vů����9�s�����a=��~V�9 g.MZ�Ō�ё��ڃI>ks���C?䈯"9V�5�Z�w��qH��K�K�?�Ӣ����Ȯ�eo� �Ej���o��N7�M�[�Ǚ�f�%�0L�Lv��Aw����q��"��Aa`��ѣt�U��okC���*�2)��L,�_�G��O�K�~�u���0�u�<�^}
ET�h�Q�2g��ԇ�r��60��d��@d�D
O$�r�r4n���o��G�q���Qz{W�.�[�	�s+OtP'��6�P�Y@��~gH�(���.ɍ��"�O�ϣ$�{�]�^�z�I ,ט���v��� *E�N�D��;Y8e��OR�yt�t��| ��i�ˌ-8�%�r�t�#���\:\��˰V��]��H\O�'�Xk�r�b�j	@�a�/6f�n����a�4}g�NW7#
�Y�N|�؉A�{�D��$�)1�?��	Iz��+)����FN4T��:vOg��<C��8GÐ�V�_��{��'��?�z;�B�����p�mM8�n����V�܉�?b,��������ً���R#z�^�˫�!BK$+ϦHsE]��2(�c�[[`�Ȏ?�I�����en�p�D�!ݼ�p&����/�X�ѻ��@6��]O���6�<~?r;)�50T����'��_pq�W�s�Xg���al� ��u��X.5��C��"G�Z�������3��e�U]��!���(���m<�'	�lL��R�$��S8�M�o����cj��(��&�[p�0��a3�#�I뛐��}���d&-�l��L3�e&^;	���f�W��z�O=���b-?vQz�(��t�f=���,]Y� �|R#c��b���.�?����ƚ�C�-�>o�Y��v�EoE������.��1�ʷ���"�3#	[Z��Q�l^8ي�@���������ۿ�ݒӌ��Q�k�
���;�(F{t����i ����Y
�KʀN��kqV4���ܰ���^5��1��%�m��p�m��i(7a ���Rs2N����k꒳U�h�X#��)�咦n�=�	.���#�8@z-��C-���t���� EU4�0��t(g�P�ҡ�%���Ǹ;=C��@+�`�4���� ��v� �Q-�j� 󎙛��&�M�νբ�.$�`��E��B��']�rz,[ɜ��g&�4������E�Eɖd)<��V����Ƴ�� Z0s!w���9A���zeR9�6f���V�n�*x�ʱU���0E��7��Ja:ց�f�0���S�WV�ْA���㑍�}"Nޥ����ã:�l�tjON3L���?.��֩�2	Jw`��f��N�����ջ3��}���Ij6��ZU�6>כ@��*��z�J�ӑɨ��]O�k�ϩ,�[r���߃S�s�P!D&Q��#E�[�5qA}�C����ki-<d�l��6�Ɗ���~��	��g|_�V�%,����_���~���L�|��y���-*���J`f1֔lU/�ƵJL�?d㜈�j�*l5���(�ʋ5����
�8In1]-���gVNs4�"���*���-ݨ�u檳�5,���?R!�:�feog�C}p�X&��33�(-}fx�ےl� ��{��^�0����@Jդ�����b�!�p@~f<��������si;�f�5��R� T�I��p��A���f�|��@���ش�j+e�5�����ҸṘ�iB{X����&��C�١M�������v6=q� �S7����Za$pi_"E�<%E�w��4=�\7�/�i2s�֣�����iVf�K>-̢i ǿ 8��W����������C���C���hta���{���N�|Mh�1��C3z�q��Ŭ�ZU>ܡE�Y��mx����Vy�1~����a�i�:�8�~Hn}�f��c_�O��Zԣ':5yc�Q}��6��$�Ih�@a�zO\���tܜ��a�[
?�!������ �^�(�$���Z{(�37ݫ<����4����k'���M��<�iY~%)P����d�����'�����j`����iQ~N���;���(a����&�QȆ�Aw��
�����o���RCA��D�D~e�֏�l5��/�b�"��z����v���W0C;^�rB��S *up��j�ޱɋ2RWJ�*������wکx�<��������,q4^�J��H�բ���&���o�Œ/-���I�k����Ib-O~�zo�+� ��Y�}�?%t&)I�����I��B+>2)
ԗ����hyg�85txr�����蜚h1�(W
"����T�\�\�g�Zz�i��_�iT����~@''ٸ��õ����w�M�D�߉l�S7��y���I�ֹ���Ѱ��NC�5�崩ݷĹ3|�+��@�͘��\�>;4�$|���w<zq ��Z����*K4x���{MK.�3�r��t��D�w��
���5����t[��%I��c�ۂ}Cv�ٻ�s��_N��[1����jo����ȑ���
t4T����y�H�.�L�q�jY�PZUΎ������$�KL=�jGn��ɖ��ԥ�	O-�m��� y�b����tuʃp��@�H7(o����KO��b�����Kk�L��<��<�~o��ߣ�{@t�(ٶq���h�s��S�r����v�lB����?!kn�]ro��cA;6�����#�'@>X)�O�Z���?�	I��>,�S�\�^⸸���Qu��J���.��;N�y2_��~N�gG�Y���F怎���ɿZ�����]�4�m\��/ ~WU8I޽X�*�$��{Q+��m��x,t�V��_I눼��=�+Q�@�7Q��>��nk:�|�'��zo')T飓2��B��[��w�A��Ƹ��{i'{NѨ�_��O�◛jsj�>>=)ǐ�}.%A�����P�b� ��v��-��D�P@+�h,���`�j#,y�~Na/��n=ex/N�θnF�G��g���WG��܏�j��O��}�"́�(x����* �@[��^��B�7�R!�>h��S<a,{a�� J'/��wMP(<e~�S���|�&��Q�G�Ep�X
�N��tt�� a"ry��hf�Eh٣~��|�M"�n�<Х���}DO9,�+m��vo4�hsdK�C2�3�[��	�VN/R��-Y���M�'����n��x�5d;;�n�ǋ�n5����r�KރB�0�ݍA4 ���1�])�*R��u���Dt4�4��@�i�,�B��iE]h�ӌp�.XH�۹Y
�i����ͅ5�L&��'G�i���U�l!򐮽 �XO{���t�j4m�d�"��S���DG\m��R�.6
��H���¸��ϲ�p�i�7��R~����;�&�g�w���S��8@<F �
�LO�5()$�.DL��(k5�,.�ԀX1R��y�l�:V}+?���L>θk#����P�c������t�{�����a�m�#��6d<^�B�W�<��Z�:�\WHd�E/�1�1�b��!�m��r(��"Dw8�7�����D6(**=�U<�ڃɕ�W!ݜ�������d-�|�p�����E$�P�,Á�hO��.h���t�꒰sx��z��1�mp*~^���e��%-��M��c�#��2������[��OӻB^a�4��n�L��.�I���y�RX&@L�Oe�n��䍫���|��[�/.�\x)�ʀ��ü�[�n�|���N�=���*�^���&�{�w �J���	�G=�݅�Rd"�-,�{\r�eT��ч���c�P��%w�K���"������[>�l��_���^=J��5��a��	oV��W1b>�JK%��V�5��>;f$�}'���'q�A��{O'��=�Lè_�����d~G�|	�R��U�9\κ����Sd�'���N���e{��Њ�Îi)��&�U�Qka�X�N�UOw�@�p:�K�J�΅�\�A:�}�yK��/��U��nwT�*�}��Uw���n�7%�m9M���IΗK��g�\��CR�E�x�����K3|I1u��,�/6����@a�%b��8�Ն<V�lm���R�X*֡fxL>ݥ�,]�H��%�}�!�0�)�	�H�
q�c7�j����|�p/m��n�5m
<���X�Έ��i�D&�����,���U�S/�������>����d��d���f�'��%w��࣫.Guj?��?{!���.��F0�����ي�O7m�o\��b-�i^��V�gy"{+~�U�e�F��LKG�-�m���ۍ��d�����B�V�sO�pQ�_���	ы�a�J~�]��Z�?)^�������o�K<2�� ?��L釞^.�᱈2��m{hs�l���G=�*L���`5���H�/�+B�Ё��do4b4y�:@�	��"w�����R�.��K`�=ʀLh��Q]Fx�EZ�E�tcN*��1�<�����Wv:V�ڭ��[O��R3R��5���C�@��Hd������|)|ʪ�����M�d�C�xg�^�^�|�/������}�}�ӱ��<�z���6�q��9:SZz�U�[��7�0HnA2G��PXZǫ,�����+E�L�)E.�DBX�K�4K�aD�����	+�(�-9�E�Q�,K�I�m
��p;��0]�b|X��GI�ڇ����tXcQ40*�IǬ�_�S�C]^թ�n��Vk֧�	S7ʟ�y4���V�����?�#ͤ��T���{��7ܥ �Y��]�d��q�������y`q�<L�� �S��ׄ;h\�O��|��^_��O��ڍ9r��'5/�ݠ_m�S�����pq�WY������Ȃ�r�{���z������v��gu~95M�4����d���|���z�bV�xҼ(X�-��]�������Y��X����ӊv�bi����y�ѩ����/��A"��'Eɯ\�>	���p�sϱ��A�2��^:Uz�C9 nx�m���EZ]��z�����$��<)�j ���vO�����F蜽�C��Z����8�����Gk*m��E���vn�����ǁ!��?��+��<b����z�9P���a��ID.�*f�a�r˳��k�y5=J�#gKH��g�^�E�)�<��K�q�8\ P��oQ���G��gM�2����s�1I���Sk�vo�$P�S�#�����@i��N����g��j�|:�5���
����!O�u���Y2����%��҄Z,�A�N0�ۤg�W��o=v����� �+L��DE�SI>eJ���X�ƫ�-��^x�)i�g9mp�T;��zւ(�V���RD�"��ívj��!�~\�j+�֧n��?�y��ub�j	L��PHU{�2�^��b�}�������`[�T|T��Tiq�����xLH����M>���	�ͼw���I�� �s�����Nž���y.��gd���P�âJ���#�|�|?�:�\?�Nj
�O%ŧ8�Ճ+��M��	��릋�^9h�h��)~K�v�ܠ�������PyK �90���a�mg~f�J<O2�V�G"����of�=CZ^��J���b���{<�> �3S�X�spС�%�F�p �����/N�r'E�=��rД\܋Wѧ-h>&ē'0��/8�IK��I��W��@�8=/ E|"�|�>-؆�t�=QL��������<���"evF�R�E�8�M
?*���15�׎�U��j�?	S�V����rZ>�GK�B����<�A��'�@t�CH�6�X�sc�(/��������@�3�����4��(�S�.�&���vn��d�\������v���J�V ��uH+���W/�s�3�E �Q�����_c>�����+�"�6��¼��u�`v�S�5a!���|҃/��`�����Vy�2�����{ohS�s������)�}Q��sf��uR�^�#�B��1���;���R�V��w�V�//̩�"�O�>h�m TB�20�
gʵJK����F��2~kg�h��;�{��b��N��Z�(�%rq��=�x��1�0��5!+��EV�aD���ɝ���Ty��*��l��Ĺ�Oa �h�"b'�9/�Ʉ5���Ȋ$HrR ���R�7t�J^3�G�:B8�5�"�M"�K �Y��u��ؼ�?B��H�k���]�-��؀Q(��C�q�J��'����������k�	v�W�G��?6�nQS���N�[16�&F�,�J�]m�^�w�A{]X�=x���BS��-@��'�N�.4YY*�OM��)��_��4�\��W(ZG�^�ɱt�$��K_�0緶�������A�R�Q����Mwa�r���}�f��C���b�J���m��p��ߢ,�x�b��(!�I��"�kj�: ����*��H�RX�2d"6"�ѽ	�x_`� �xI��8�%����]�L��X�����.��qs���Ǚ_Ͼ����E�������V<�I�za��.�h M�>\�P��bٔ(�D�x��Vn%ֶN����?Ԫ���K��Mk�U�����廹�ܻ}d����k��|��_;�;EA�u�AT8<?��֚$��	�A���<hR�X��+���tdi_�����s��ca�Բ�A�P��!|n�v�/��b�W��~��b�}���,$!���적��#o ��O���p�Q���)܊=����ϳSu�5��7�������X�@�U�v�M�������wP5�Y�d�])�{�:7�:0�J�-�۽�L��G6ÑS\~�=��+o��_�X�,��UV�LR7Z�+���B��G�3[b��C�N�l�z�=e��_��� ��Ǜ{'٩}4M}ʥpyA��׬o���0���U��s�#[*.�j������R@�v~���DN)�UE�~����Yoe�%�`�X8��#���l|E�O��긫�M��I��q��*+�G��W~*%���ܽi���]���d���2���蒧�I�:�<��p�?���~�*�}�r��rR���E��w��A��년��I���;��í{�B/���
���3��/հ�,ѯ�x���a�X�'k��І-S��F�������l&�<iC�Xn�uG,����U(��P�g#ք?
�ݹV����x��HcŅ҆Ɯ��j�!(�js=q,���wE�ar6u����{���Q�2�L��z�iZ�9ej�@N*P�m�뙌�$_�߻�w=�{��/�D?��g0��2
Ū��d��ɰt5�q6DM����ߝ选�x�M��{I���LT���);�r�W�Y�M���N����T���ЪΜE\�[iÝy.�(��O�����<,��q�&p1J��DW��+������)z�	熀�%�����䵖�A�?JR*'���-�_I!����G;5�R�@�M
'�̣��k�r&eJϢ����}Se�-�L����E��eh�(PWgǗUϙ�QZ][����$7�zR̊k�wzB��Rt�jx���Z-ʺLnt��\Ҋ��K��WZQ����=a���#$ư.��_�hl�����i���_�9|҆��dF��j�]�)�66��K�6@p��V`K-�������)V�O���
�g|h)Ů`���3Jh�R�vx���RK0��
�H$�@
�}���Ƙ�p�-�R�Z5a���wt�����!��+J�"�7³7�D��Я�u�U�@�!�����\�[��p�F
�(mp����^׃��C�PM'�:Q`yo ���
�Ȓ�Hb�قӬ�j���T0�\X(�բ�%���Φ�����B�/�=��¶�2��B���w'�8������:I�S���M�| R�z�����J�\݉}GO[X2�AEĭ;3��-��U�4%�9�I�Ptp���3Ѯ.��r0�]}�o�up���k	���8Ax��I�Ą�:)���M��@,԰�B��u�m���A���>�L��v(���l���$n�E���|�{�.�!�kuMk���I�B��3��� �P�@r\�Ϳ�Y�E���;�}�iׄEr/?�]Y�dE�|�����}�ݦC��o�E�r�ڛ��	^�۬WG���£�q�-9c2�yV�D|���E��j���;�+�ݠ�G[a 60,�J�Xĭ��c	���{�3)���D�Sd���7)D���ҩ{�u���{�u��W?�,}U!
�K�C�h�(M�i/�#��ً|�,�q�G��u�'��i��߹�/|��M��'����|����iM�$6Yu�*-���?�>u]����˱/�ExZ�nsg_c��EU���7�Sk��W��5���Rd�I�T_�%���h5����P�����`�Go|���N�>K�-�~4���y�!7�H?���{��LY]�����vt��;H�wӱ�^�S��_N�g<a����z� Ōk:}L�1��ɶs�J,�f�Hޱtj���Nr=���@� �R�~,d1�G��Q�	,^�/�S���N�~���_��.��:K�R�'I�k�LZ=��~{e����da��&�����R�.&3�Jv�!,Ѵw��[��.������/���z�Q�]f����+: EfĐ'��.p��T�M�]��N�M��;�JE��@�t7F����1E��0�����w�ǂތ垄FMN�鳡�쫫B��F}k,����\��ϒ@m��pg���W���/R�d��۱h��3�p��J�1<���f�>��lۑ7��MS�~	+�M�d��݆�y]��5���0��$�ԭ�BI�7�6�l��_��Dj�η���a�N�ᯭ8tӫ>PBEGt�܌{��`�E�К4�e�����q(���T-�Q�r.�	C8\�W��OR��� �.z� |��ty�N����ukp�ðk��"(=Wa.A��C�%u[��R��D��Sfh�Rx���
���~y�g\GA֨HF��ذ�K�Ao�+_ީ%СB߁-Tg��o1vx���:Y�Qk;������Ӯ6,��P��\t�? �,(�%y�"������F����,V"��
�����+8B����;�gH��ޞ�Ŭ�9[ҫ��� �Q�E��As��3�$O�s���7]թ���yN��O��1_m?�s�e�`|&;�Za���r��Y��]ɔs��ܩ�W�9�.�6���{ǐ�w�Gm�o*�7wӭ	f���W(��:<r{�e�狯$���'�S����0��(LA\��י��ȆWU���;i�9�Og��Óƪ��I��]�d�����H~`�UU
�mO=		\hR�`�SO3�E�OI��N�b"�v
�j`�ba�/ޕT�,��gG�K^q����#h\֘��L���/���W��9��F3פd�\M�Ӿ��MJ���C�0�͹n&^��!�s(!��JH!�OR��Q��h��y���7�L��]間��?p�(#Tɭ�Ze�,Ć�� M�}��Z��^��J}�h��Fl�%�㹖�R������a�H>,� <hQ%+�4F��#C�Q oT.c�Qjrr�\���<�v���;��4m��X@�`���i�b+� A\h����u1 U���S
�E��h���wR�}�	�Nq6��t(�Vxcp�?��Uǲ��^`bW��/�Iқ�G�u}LZ�	��ͮ
	ĭS�f<Ih�Т�[��u[lz�}�ƙ	�j��y *9 �:F�6ـ��S� �y�^n�p;���Z	oG[(y�5!��Fx!ꎬN-��8ff��e���ǦR#�>9�m��:��['t�H����zl��<aHBf�%���ѳM�.N��>B����w��n��
ި.��g��zf6�|8����	�PBe�Y��Y<qlǨz/��x�}W�Ĵu�n��ٰ�[��1Z������W	��wy'6��iK��U�'��8��r��'ED��`��V̈́�j�@�&|a&8T���-�K������3�V���y�edЕ��t������c�x�8<6l�ug�o�^�r,������R���0�N��$�-B�x�)r<����N��zRm�4i��m&�Yn�YUY��a! �<X����Ӵq�y���{����}�����i�'̨��o!�����ϗtj�k��9_�ܙ��p��OV�sj��+��١�V�xVb����P`�>��3�]! -dX���:D?�j��n@����D��I0��?Z�k�!��k� �[�߸��¹�ܠ�6��n��z�*K�g�z�ץ��Oi��v:5(�a�����o��l ��M�H����c��+�ne�'Ҹ�Gݳ��<�%F2�"H5�f��'8���X@-�F� �l�}�=!zM��g1��~:����!�$��O�}�by"t��XX	�)r�]|�G�����3�R[����YԮ
#���!�@�Tf���q>[{�Po���{�?��%w�e����6���G�`ɒ?�Ǉ����o�����B�����N���J��cE:;�� q��)���:��>��_|���=�H�nI��=�34YI��4HD,����ω$`@������z�ol8s���I�%�w�����}zgO�w�0|�߼��Ir���A�R�fOw�����n0��>D����T�6)Nu;gb�r�Ӓqo��@_�l����5n͖^��ݚSD=;�gZxD���F�Lq���}��2������Yɹʁcb�K�1�a&[|Q��gr|}��߶�bYg��>x�W��u~��bE\��t��!�:�nr1���3����bXh*�T
�Ş��Tp�iŁ��D����\�t	G�1����#X�����c�&���9  �5%e�PhU��i*��U���� ᐁ�P�C5��.f��9k�ؒ��-<��k]n8�}ӏ�j�e	�",��_��a^�a�Gr��C)�/\>ב���ȏ0�!)����6Oa��>�\��E��దK�x�"��,L���V��gϳ�\Қ�iʤb�"ry6���-��\B -��m�4L�L�MHЖg�IG����:9.�U�*ԋ��#�\���� �Iw�U�_�[c�k���̹���	7��L·��!d��&atP�~:�v�Ѽ��.Cϓ�b4��a9�C�#����HHR���b`��X�S4p�H��0po�d��'�ՁI7�E�PH�Ŧ(�������w
�㵄�=���UD��a�<,E�c���q�/֗Q�L`'XPә���ꏻ;4cs����Un�]QJ�OX�:dP?��=f��
�\��曲M��Q�ׅ����H�*��I�,���6&�$d�5׸IZ����I�=y9�1^��u)��E����4a�/R���8�dߘ˂ǙȨ�=xZӣӦ#hp�T�Y�h]���#�
�l�)�l.��
�	�]_�?�jZ��pV�j��
��/�*�*�PR�ŷţ��@��=�I���� P!�1x���t�J��QXc�ІpBFA�Z��-H�ԑ@T�a�AspooۿK�'�p~\���	��'"Yq�p���49�⡼�әM~K����?I��xE�k��"̻��ElGU�+\""w�?�����[9��|b��B;����<�xUk�q,w������r2�g��l��R�����)����G�I�
��@������2��]�mNç����#�{LðH��l�`V,����8��0l�YlC*��E�ÕM&��L4�d�cWg�A���o0h�\��2��'@��\�;mT��Q���È8�v��x�p���jؑ�ˆ8�����n�~xR�7���θ�G�J���</���� A&�,��Br��m�՟�	\�%a.?\�~�*S�� �˹k~7��n��p���0��*�l8Y��N������#����c	u������k�����kK!�@�(����y jv���-Ų����i �[��+�ꅰ�Xn'+������s��Y�P����ф���f�7?�M��Ďy�^J>Vߐ�
��E�2r�2��2�����UF�����Eq�Q�+�s���N!#8Z������������ud��{���S�6]���)�F���T�K�Oda�����)��bȷ����O���ƒ����f�o�|�8�����0O�����\Ď��|OW}h�|Q�L=��N�J�F��SCp������� �`���aE������^��J����Q����7a<d;{p�Z-W6I�3M����g�['R�l�H��������J�����-N�p����t+$gP0���}�n���,r�hf�{p��������\�l�n�)ns"~+5O����Y��I��t�E���b_r����Q��[q�o�[�V��CWv��X�Y�[�I�_�P9��cT����qN�!�s~�N}����A=T}��~�z4���V�+�#Y%�d��m>ǂ��\7˵&�L8"�d��,��������P��ߏu3�=�ҩo��aۻ�i�Z��o[������H3hU}�Ԗ���N��ܿe@M]�ԗ�uhʴ-@��7�����@K�ǺE]���� ��*O*�V����8Tg~	 �m�/(t�~�8�Mj�b��bL��ϼ���o�U��������V�["���@ ��4����unC�<Ϋ��֠ �B���0)������]�h�7�X�Z�{�/�5f/�hШ�]?��{ԑ���z��i��9q;;?J͕:Ծc(�� �,q}�o�q��o���ہK�U-�vK��]��E��Q:,(t��T烎�2�qαE#��D%/?y��}��~d��a"1�E���BejzY��0�;��ĳ��'�DQD��D��[F��A`��9�i/�ě��x���(:�V��n�Q���y�ڊnD��N-�&O��qH�)uݙV�[�D��,&vp�^�,2�D ���s�Nv!�/#���'��)���x�~�Ɏ�-1���ϡX�9�~u:�D
������<X�}��䎸�jt���Ko��ي2�Ę���>ܠnKa��,k�v�0�-7�t/��F6ߋ�@��څ�N-q�<�X�B�������u�oAv��wty�hw��d  ���r��R�I���z�g�AFi9�Q"Zŕ�S;p�N���!,$�+�[9[0B/p�W�C�5;RS1b�_��uA��S:�u����؀pɶ��;k���gM�Hdo�*���K��y�����@X��s�a;�u�1K�C�����Ek=0�2.�����J��ż"�boC6�Wh��#�0��O+�q�V��03�����>�ΨA�� A	@}~N��, �bX�b��h�4��'ݷ����D�W�(¤���Z�����ژ	"��̅��щ����ȝ� hC/�y�Q�R��Dq��h�U��%ӽ"ULw��8n;�C��LV-Mb�ֿ,E��w͏U�k���L�0[%�5u<fD�ڻ㽏��~�<4xbz��m��z�=H��R���ϡZ3�{��Ě�d{�hl��2U����J��Z�Wn!J��sY۝�R�O)��WR�i�#��"ӫq>��5]h��ե��@
���`�\W{��0�|��7���)��ͧl�>:��~f7�����Q-�z�r�� ()�:���֨:�K�O-k�����z�D�>L�Pʧ�63�)�cVm�^�?�Ż�w�6^�ˈ��uF�ƹb����vcG <�0�?��9�i��hQ��Toi~�|JU�X�gZ�(N%a��4	��`��c�����W`��Ⱥ[O`���c����uz$�\r��Ycc˥�(�!~1=�Ja7{J��U
0E�|�5K�ēi�w��P�^�K}�ҩ�C�E�	u$��K�u��a2´�� �����ge1�����0�^<�@1�!���ZB�(OED%�ya3ŧu��z��z[�~�O����n�{�٢���m�e�ɨ�P�'D�,X���|8��^×�.�z�gȇѴI\�V���HV`o�}�ᄋ�ec�VM3��WNj�!�����0��8.�$e����Ȑ�4�^7��Ef���"�쫻���$͞G���G-�O3l*��D�үŘ-��q����9����������x��y�8Y�H��鹯�i/8����?���Y�_�?�b�l����΄?��OT_=�g���5���d�ȵ�s�-��)r)}�Ɓq٭���5�	j>��5��V\l~���3��um�B�:����
��ۊپXfI�llM�q�H�r�?V��ي5�ܞ7������olM�e���=��B2��_��k+���[�c؅!E�k֝O��v`.�}�CZ}�WnI�)�A\;6�R�+}��q� ��R�G'���Q0ӻ1%�BƤ�5��Ԏ�]�@N-�~�� ��̥������p$]�~ay�+6�9��%0��I#m1<}J�Ī*���迎����Gߣ������S"�J���H�+C"�2��������e��Ifx�:�j��W�crS_o�!��<��)�X�[��ֻД��[��GM:>;:����L�H?b�����m�~ ��H�+��f-vW;դ�V�"oi����,�ܪŮ����r�}�vaR��
�v5cv�@��g#Qw�aʍ?'V��?У��WO������S��㞋'�Z��c-��"Cq����~�%�ߧgc������w�C3{#��,��5�ʴZBϋ�m�l&�����#�S��o�y i�6/��ŉXMq�~.�(2�"�%FDP!��Sx�Nm�U/��e�~H8-��͒��u#X��Ԛ��@��ES\�n,��քܫ�O-��1+3�m��8��g�Z�c��~}��FBxB�>ZlU+���2>��K6	~a{2~�i�t��U�����v��;N%.�a�0�[P��i���1��u�_9�-l����+z��w)��d⓿��[�ՠ �mx]��L,��٠��W�9��7�Xq�O�8��MC��]��EC�˹#x^�X4�c5K�C�u��c3d�ZI��~.�^y<n�!9ゲu�A*3��.���9M��g��F��.a�킷r�b/I�ԃ�M�%��Q�kX��d�8��i��=����B�H��-��5!o$��\����Ыi��/��|�ʅ�RT�u-,�?�O��|")ȇN���]�1�sZ���ߋ�,�WnP�=�,�Z��N��o���\5�&�oZ�di�v͖w�������b��؋-�f��^t�Ҙ���B�!�@Kb9ޕh@0JD��0�ؑ�l�>�,��'5�H�Z��F��y�ZRU�Bb�E���fݶ�j���/����j@*�M^�D��E]F�L���&_�{�)iIl!�1 �̀m��LԿ�_�2m��4��=�!'�e�غ��v[$ăm2�V�j�1�`i?�n�vV����{[���ㆶ+�����O�����0����ƛ���iԿoU���}p�L�s��ޅ��Ξ�'�Ņ'H�Zwb�N�����Fa/���yX����jp��S\�)=�J�=n\L7�TtG4��-lK�ni5��^��_��8�*�W�S����H��3H-)R�O�a݂�����Y��%�+� �ԟ9m�s�@n�̥I��g�u�����%���T���E1?����Ϝ�e���
+4ё����L�����wcAX$u���c/�d���QsM�)�g#h��i�u]���R0���a	5��B��^	<�z����~���D5��A��/t��W��Y'|/�/��x��^a�dW�w�7=�7��渎�H��ղ׺@+��k�%[�4�/��f}6\���4�Έ��(�wf�'VY8��t�A�wAz�K��N&�S[�u)�GKB/�����HM^(� ���ڭ��t	}�H��~�����>p��%�'X�]��yDi�+�{�8є�]���.,®]m�1cir�*,���!a������ɷmL&�����3���h0�� ��/�m=F���%�RX�$2������q��m�$^��O^m�P\5�Թ}�C_%,P/�@��&L��V�M���y��c�y����^f�.?����d�Ǡ�a˔�LJ��+ug��z���_�5�	���H�����_���x��*�G��U����,3�zK�T�T�Q=N
wR��_���W
�"\R��L�3a��*we5�eg�;�t��{�UZ�Au��#OM��w�֦[�����n�\��W��>�ȹ;�KO��ݖd	���:�}�^���)���w���8<c�͕��D�1���G�1�)����&eF77��u�_���U]U�H��&Z��7T�
 x�v��L��A ��q3rfH�����p*��j�6������o'�X����m��-R���;�a����~��e�S�|�C�[���:5���0�U	��a+B�ޝj���d�9��i)|,q���GX�E��j�Gb���^�I�>�/����S<1��=fTuw��\��»��	)�'O�N���%����l�}�7e����K��~ M��tE�/K���lXP{:��?Q$�{�[=���c�ʸ|ot`��e�2�u�ryw�����N�}Q�簾�W�S�X�����ᑿ�"��rW�|L ��b=R�� $�LO����^8�v��ʲ���}%?��,�$��`��\����k����?PMD]������`�';4�t�7�JFu�$B��D��39� �ԏ���߈�S. ݖXYp(,3I:����<����`\��	�E�����:�PKet(���6Qo�W<S�7'�)��[ՎE��R�Or0J*�3�&��pCa	�Wl�PG\��(y�T��H@���R��¤���P�k6����}��'( �C�����/=���bC�"�)��-��h����O�����jі�.�6��b����u�&.8�6q,QY�X"��5G�>ӂ��}q'�"���,�sE_`��u4"��g֊�m�Z��cN��8=�Q� �
_�_����,3�`a9�����[�S�oK�0���^Ŋȿ-q�1�1(�0���M�G�
����x47��*�Vx��ѓ|�� �	J�����ݿ��5�O+�> p�_L��2^Xg��t��՝���1v3T�ʅ���K��>� �J��:Q��5���92eɟ�䟛D�X�8��؊� z�� Cw̷YvtzKOxkJ�Z�b��r����-�n	�]��;�P[�T��.l�xH�_�	�1���U�=�Y���ҳ۰�p۸�V)��(4 /t\�h��'<����@����#� ���8�d��#@��\b�Ğ���.i�PnK�N�e^�vm�/��iq}�!�n�s2�Y�~1��y�f�ߪ��<�W<f4��j��n���������{S�>�g��,g��h�?YM�5��z��Y��scj�A�4K�z���n�ݙ�p�u8R��N�UbuX�~��}�P"�hF@�w>�N������f��ҋv��,��E��7���p$%���l,��l���#wH���gH�*}F�[���G��-�2���`���y�� �¯�'����SpF����,��Ѡg��FC�뒘N�b���b4i�-Z��<��zX�G5��۽ʵ�jO�s�~H��g�h����Uql�i0_''LϣF_��Z�K�QTbwf*��4�O�/���ܙ")'�u�h_����5��"V�^����>|6r�w-a�A��7J����"��z���[ܷ������Q�O�}�.�����������̳��ة�v�*�R���4-�LS�in���EF��c)ݓ�E5[o+��< �N�F�<�z���@\3���K�Q�""���9�&K��	%6u�����'���0�'_|-�7~�#x��"�J�'��	J�k�m�il����m�D�$�r��wt�`���h��;��H�´��Ɗ+H�68��ࠦ4i��J:ch3�����+���ѧ��ߏG�ϙG�Z�{�;��S��'������R���|E��'�,k���g+S+���$t��I�vT���y�Λ.�teZ	����r��[@@����@X>U=��|�����9�|'����9��}��S��E�d�c�S� 7���iAy���@��Ѥ'?��KBo�b���Į��ѿ����▫Q[�T�s#��'C���a��G|K�T�;���	� �+�7�o2��g<҆u"\���,$�؋S_�(��G��{1�X���b�j�� ��H��vp?ɫɮSL����W�a�B"U���H��{���_����Z������{�A�W/"g����Xʁ�����6��*���D��~~?<� �;�x��l8��HԘ��C
׌KS�|�%u4���sO��QI�"!x�~�dk��	�|g1��x�.'w��%xT=�b<���0�9y|�[y,�:j�����_��_nGѶ��d��R$��]^�;�|ħex��s@������)�p)�;"[�����?ӽ���E�uu�����{�B]|���������$U��q*���W�[F��1��@��(�h��SK�c�������x��
� )���ǹ���l��㍎����	�i|� I<x#j�'��:^�︖�ؔ$��(�����s�%	�����j�>�ǥ'�s�Y�ZC�}��?`��?!�ٻ+�	.V*�zMP �)uӎ/%:��g�C�K+{�sС"���th���spہ�ƍ�z�F���(�T g@�^O:��;�%�~��פ���y�t�2�\c��T�]��ڋ��z�n�:�_�	��_���A]a��wn��.�d��{�U|������N��sMjO
[�K�9�|��#��fTj5�+z���$�D��.\��ixt����Ѵ�`�� ��AB��C����V�Pc��+��A����tG�O�q&�Y��-\�/��$H�ա'�,���6�N�!ƞ9�ۍ���whn��YO��+�	����dg�����E/�#��.%�AJ׏4f���\uҍH�6d�۫��\���a]nGc+Ӷ>��2ï���S��X���`*�&�%A��#����5�_q}Gn��崩��`#�z�@�,YM>�U�����"�ܢ~ڗ:1�RpOw�`�+�M0���q��O�y�Y:�>��n��A΋��rs����:iAwm?^����ٖ���{V��;6�f�� ��Jv��xX0�V���L�Z��V��l��g�o��j`�;�$�'����Z�o��\��U��<���_:���Ba��.�S�AYG�p�G�zY���{$�T�ݵ��p�5�D_"
?��3��teIKW''�.B���POQuE�G��L� �|�N�m��/�@�(���	�lTk��u].��JM�)s1Ь9�B��V���]�� �E����m:�@gQ��iЛ����7�3���p�.26)�g�TTW�7dW� ��勷�(�����-�#��t+�?��ÐS!��K6��������
ki�U|<y\_�wG��u��M�/]� �4�]�&R��I<�/����mT<�����96�c���{�:r*��
#��~�I᷻�roj�u��G��ݙ�����R�{!˿���ʹ,�^�������(6��Q��Q&�J�=��J��\$�p������ ,ʤ������I�DQ�=0�����}��)��%�
HR/գݍPD}䋄�C��E�_�ѪJOE\Z3srښ�D�e$���i�߆Q��)Z�Iۨ\��e	��'�B"~@�'������hi�[�t�%�*��#]� q��@/oR�m��"lPMӾ�Yt��+r�U}��Q��m	`�����s�? tַ�������4��7�Ȣoxԫ�f��̧�R�#��B������R��.&��|s(�\WBe�i�*��0�_ck���0�Ԣ����(^V&At�A�����������N�=���/ۓD{����ٓD{�����	�O�����H|{Y�*(�m���zxv6H�$W�F�������Z.��������o7�q�=G�r�{$8��U.���o��gK��4��z�]4Z�i4�5P�>��x�g�Wz���<2V/��UB�dKn�.�m�(Y�H3���҄y�էPO�]�)K�[P�s˳KH.�̳͓�G/�uԔ2R���ˠ\?ԡ_��`�?�b�>�l3y��ŵ"�U�H�{�5H^�)���.6��4�N`��v�8w���bC���A�ET{l���S>����o	\�,O��/R�pC�"[)����I��b���3>kQm՝S����%�SK�" ��` Mz��cSQ�6�qɗ�]����I����	e�y6q�WM�%2� {����= �صm	��2�JY����Hh_2�D
O=���\p!�M�]��C�E��F亏�ey���I�#y{����]��:���]W5~R��w�� {珚��ڢi�b��oR;�؁����K;�	^��9�߇��?^0��nד�Y�Z��v����ĩ�VviԨ}�ITS?\��0���L�@C�t��-p�3j߃Z���Yu�}����p{�ؐ+^�gF}yM��������%֭? ��W�<ϱig����>3�����3�!=:)�'9�l3��ޝ-�67���6K��C-����vB���Wc����p�,��C&���Yҳ�a���HXr���.� ��ᆤyNT�k��\��A������&72]2��%Ӱ��ɩF^�a$�0�z���3�K��]�����4���B�bb[�ƶF��]7��m��77��m5�L��k<����Oh<��'�՘�V������}z�����O�}��e�0��%sp���8�-�I-�~��mj���y}��[�m6K E�T�Zot��3/%�.=�T=6�V<FPR����4|�MI�ڃI��-hxm1Y��;�l1c��Ԟ���qS��	�Iל�B�Ѥ|�8�wϷ��۾P���$<}Z ��B>�#��	�݋��7	�U���i�� ��M9룋L���GA6)�nc�ݡ�q����R�>�S개���t�eU�ˣ�e�V���`C�$���7*/E
��[z�b�o���|[���yk3���E�?���&n�#��E���+�M��ыmȭ��$��]e�p[T��Su=m��g2g�z6���YR\~B�8����xߏo=�I�uϪ]DK' -M��=��R��*����Z�2+s�a8?_���0��uq�(���&�N�!�� ��@A�&�r�+�J"C�.�\,I��+B���@�o�:��<����P�V�Hu2��V|)=C��o�j���"k}�����*U��x&��H���O�gM_�i�4��tP3i�y�r�1�j .~p�F�ɧ��
�X��W�q��[��o1���`�\s"�����0�;�r�~�((w�Q}~Ց)������ՙ���� :��l���^�2�7������i|
�LɜX�ԇ�5�Q4��{x	��{Ln��P�W� 	��Wn�R�Ni��t� (Ճw������}l����qU=�;=~j/�r�;��XpoO�_��!�_������T]]�s;-�6@����#�h��cA��Q���/�+��Ę<>�n1���z:������b���~I�;굎��+3]sG�mnx>�M�?�hNMz�췡���G%|4t�*��PM2<+���ڒXvl
��6y���R[��Z}�.��I��л��~kL �= �M������?�Y�f����P�|6�|ze������Q�\4�Ol4R�@���ͣ����\��S���ĀT9��k猥�:p/���X;�P�=e�E�.�Yt�~���'�������2H��!�:��= �����}�c��B<yc�Hظ�6)|�@�	��D���O�g�)ԅM��;�a)�^����	�z����B����z�j�9x�=X�Xy{��]�����m����P�P��=�͞�L��J��O؆{����%8�E��ͭ���vq)=,Zς"��C��UC���jŶ��a��Mæ���7٘*��� zm��� Gi����02��M�s4���xAeN^OÔ;ZdS_���"��8x�UW+���[.k�:�F���wTߞ ���V��a�[v6��z�{p6%ƴ5&���e2���n����Rߤ��q��2�I�C�s�/h�^!�H��� }rH3A�zC܀��i���u����\�Mt"��u?d)��u�ڻ�\B>)�fa���S��Y��C�"+��l��O�5����:��YL��ᨇ�qt��$��S�K�׭y���U��`��q�5�Ӎ�;�P�k���a8mP����ѷI�v��B��jfJ��"DI[K2�
}HC�?sP��{ԍ���OC֭9�<Þ�K�s'
���]sCo�3��?4z7���$�d�����Ś<yVe��� *������P�4L�+�s�s��!�e��M	��l����^���6$e%����gY0��~a4�6�3�&Դ^�y�����W~�*��F��K?<ǌ������$��W=�"j�p�\sv\R���=�?M�d6Xt�ah�lM�h-"|lT��G�0�s�C�ԇȨ��ߍk(݂哕;�������bO��Ǉ�� _�Wf'������Dڪ\��DEYF�A��I"Ɍ�X襯�_c$W���e5�O�+x��V���W��)���;b�'����i 7
�KH���ۦ���	:���L_z	�A�gr�ƾP�)��J,���L�3�0�[}��6r���ԭ)�g����JXG�)9�-�P�N�*����0�4F�h�y��ODз�jV�۹_ 궣�m@���c�ێ�?#%�36��џ(�X�hV����H:��sF
s{;S�����)��j<�p_�֢F��A �s����?	z�����4�@qE���@1��Cb?�k��?��7K�?�}	xSU�pn�� �[�"��AmՑ�Vlڄ�@�G�b���$��R&	��%���訣����2���@[@�ԅͅUϥ�hi
m��}ϹIZ�����g���ܳ�������J��>�h���R�8C��;|q�D��b3T�Ʊ�{��l���X9	�V�߲�]Z�rz���p�z�$��@!mT:{�}�՝�=4GZF8c_�b�]��p�3)�0��`i6�Rcv>,�	��t�-��c����x�^z��X��H)ڤ�*H�x(ބUXa�נ�is�e�폹�8��cqaE�֛� tK�z?���
�m��v�,�;�~��|4�H=��Ct�F�D��u�m��c#ʩ�+��/J�����Is$�.ȗX�o�(k0���-���*�x/��ӿ�Kt�p�󒌼E�fs��E�'�c�Ҕ��b�����d����ӌ���,��?3�}A3�:��rK�O�>��)l�K8=>�+����T`�6y�=uB��p��Ite~��,�ì>�ۘ���W ��rM�X�v���T�U�.�>a�T+m���$�P]�DE��_�m�8�U���PZD��8X��Y�j�	��)����=�-��{�\���,� ͸��S�1�6�g�su�Y�j�����fq���)��Ǯ�J� ~9/�V�2���Ba[Е��8�H�|$}�|�A"/�˾�@�7>Ƈ\������<M�Q{��s����|��B���En���x�T�7NF���;3��w��.7��}12���|Mfy�}6�
�z���mOJ\;ٜK��Q��Kb��BB����mدK	��./T��.����&���GMۚW�K�����s{~}����/��!�I���T]��5�3�q��
�090�J����9��d�ęح����E�k�h�`�?�U��Q�Y*���� �ط?N�W�q�,/�k�2�����p4�p�\wPO�'l�/��+�����5�œ���&�'�V��;6^�����}G�t-�m.�~ͳ��vȎ���qo���}�Cf���"�3A���Qu9]^
-k������g���n.cx��5>����3��܋qٲ�����8I����K��KQf��kSz�P�؛j�U��#f=���:���D���߮ᖬE�I'�B��#�	���e��I���I�/>Xp~����hR3=�8 O!|RW�o�r�B�A���ŵ�Q����.Y{�8��}����ќ��� ��s{1@�ˎ*���"=���k)�$!����z՜~�f���cHSh��Ǘ:�'`\��qf���� gv}���Im��@*�k``ď5v��DS=�����i�hL�[�1�(���$�����Dߑ�F�u��90� .�D.��M4�o[�����#�"�\�%fOz�o��<�u㛚�bL):�S
`�WG��Ŗ$$,�1 TﷅnWgܮG��v}���mʢ��x���X:��nW�a�}<��֓&���Im޸R��4�"�#H(���"ٝg�)�w�=��kY��D��v�h���S2�����V��މ�F�/�&���%(�fle{;���G�'ct}��y��&���3���x���$�O�u�u~�� �.���?7������e�;����e̌sRϠQ~M�vS7P�8�a�5}EÔ���TJ��p 4������G�����&��0����з�!��n��O�e�M�=v�� +fr�#��7�\ި�TNN�Py�t�],]
߹��Z_��k.R{�O�GUUQ�Ry0^	��d/{�\��#��*�s�E:��$�H���%�fX$e�f�T��;k��\ci���u� Vo�D&.�Ȋ�Gz�$��wDB)ک~�3��F���I��9������U����gj)@����_s�9��TU�k�v��[���C��\��LR��Z�%���_��I�
>���/�O��Xqm���S)R���2��y�G�1
�Mo��1&�Ey��$�.`��K7��-�7�6������D���L%K)!�I�KM���������| 
g�hiȠ@!6�Zn[#X���P4��~�:4��+���s`��� �F�6�{�e#�Q��H'���3&�s0�c�8`��yr��y�7q�Z7h׹�j���{���ذ�K�)O�h�Vi�0�x+1�y�Z|��¶�	!X~-� ���l9����p���M8���R��rv�q�e�U��2�)ࠜ+@Y�D�G"`�=a�"I�>�ğ~FnC�p&�^
?y/�k�ҨU�o�V�J�l����a%�X_s��{ �X�zG��σ�X��q�x�ն�����X��������s{�e7cz8�U56"��[��Tm����a�hs�a���č�I��7~�ߎ��	��@�b�;�j6���A��D+q'���IJ��pn�~�%����/B��O���R�+Yw��|wO������^��[h��H3�CT��*�$誓ѱ��O!��x+~�
:jE���-o�����΀b�g^���/����Yѥ�S��������L��:d��H�s�z�3�I�9����Z�筙����y[�U��f�^�����ja.�m4�\�˄��s����i��&�)#=/`��X����)���	�D�E�NJh�iBH��_(R/)e�%����6�9Ҟ)�l��}�k2�
v�Z6'����wf��ـ�le����p81�����q�X =1]̑���5m��w^����|F��>���XER�Auq�$�E�36mu¼z��7��������z�"�w�	t��Zc���M>�t/t]&�&+/�5��7�ś`V��%�[�l�����#۹�z^^�jg�I�l�k�Y��zv�l~ף�G��v����JCU�J��J
��?v�)����o]E^��T��U!����-į�aF)��8�gE[������F�i}rI��qq�j	ެk��EG�#FcBN=7�����7�ǾQ4�6�-v����^;��!q��)��Xb*l��H�VVq"�곿�q��Nz���ůC���GSz볘F��L	�D
G���d{E�=��]/��_�㳝�3����C��/]�n�wn���I�
��`��8]8�{�;��9�A�O����.C��cJ51��zB ������Ȍ��˷2J�Wr�(,�#���g{"3F絺�e��㎘>^j�G��]�����~�t�������Q �Fw��X d�&��5J |������ ~��?J3�����R�C!ᥰ#C]q�Pu��P����C���C��1���u����~i�7u�'��~�6CW��������{�[h}�C��>�a[�]�!ݨ��7��+?G��Ư���Fp%��HH��Oƿs	����(Ć��_�� �_�ǫ5Ɠ�x�nIK��݄�fa��u�/��x��ږ�!�!�0)��~�v��}5��m�\��b"{���N�t{�X+��#m|R�w֘鷺�g�䟭查Č�Ĥ A�O�����%jΔ��R4��tj ^��3�,�����Y}�OVh�p�Hی�cc��}k%ٟr=��δ����s��,L�"�<-SYJ�=�C(���w��|�]{���Sیz�3+���܏Ú���2�; ĩ�J0������+P��=��Kx�Ĉn{�Ğ�8���Q��!g�@��5mfޕL��k��mߟ8ͧ-8=Ly��d5�����?�/��!����8,��v�O��֭��g�A�i��/"������V�n��ɚbb�����Z�6�
�_+��go�۞��M�T�ӵ��b��!j���ӭt1q``�S�o9 ��pu ,F_۞Ե�^+OE$���ǜ~�1�n�Ԙ*er�^~��O	�����G�u��������!�8	�t�3�%Dv�G���;���Ύ,:� W�E��@{���㮥50J8��Z�"H~�݋��M�O;Uv�	���I������-y:�RG���;��*����6�)\���67��|�P�'�6�N��߼�5(��K�T����$��\�&V�xߥ[���5v���}��Ǻ�*�(������#i[���w�=w��&ŧ��݁�.��ɞ:�s�Sc-�/���D8�Bwm�a��l*��ئ��1o��to*�"���+mY˩�"�ҡ�rFx�A.G�z`� 	vtͥ4*M�eNEqs�"L�sAn"��lR��<!h��ߏ�&���pDk�8��:F{��Nz ��H�^���B83$(4��f+z��)����jd�����~�A�L`x�g��$��=F�{����y�.¾�<M�x��|+�(��C���"\Ƈ\.=��	K�d���Z��o�cym���ଢָ��$�t2��*ԯ@lG��.��$���Q����~����4�ŔgV���6D�=���h��CG#��7Jף��WR�s���n�N�&S���>m�Io�u��1���NJl�	d�+���׶Ζ�ЦS����:X��~���Sz�E�B���R�'e1�A�Hx�(���9l�=�"#`�N�q%����7�C����Ń�8ƞ��P�,�sS�:�B���e�6n �Nc���sLM�<S�z��`@
��G��?O� e����z�VycǬZ/sc!<mD�h�u`Վߵ��C/ �?8�ch=�� ³�)����t�G"l�g5=����!���� `��j�U���=a��q�e���n��k�©�b�P��qО�b��+S���"FX��+���/�k��a#��jk�Vu�98~/��B���O�����0/���_�:
�y�?���=�?Z�J�+g��$��K���G�p� 6��; �g�vq�#�Ѡ:��X���՗i�NN�j8������^^����z~/�����{���dv۬Pظ1,afR�x�ɨL{hP(\V0���������wq9�/���y���6,��m�#�z�G|3]pV��&ëi���T��6��]ؓ��v�#W0~p������c��R\�|f�(�VRD�;�\�������9�o�BC�J�
�d/@�4�;-�.�<ɑ���=��J�)���nl
lA��n�d�<G/Y��y�O5�w����و��E�u3Ba�3��؍���My�8<h�L�o��6s/�R���-	_��9^<؍�E�S�i�j[�cQaΘ}{R����U��^��u��.#me��'7Н�@>˸�v�C
�.c��{,�\��щn�c�ɋo��ZC�����6s������!0��ф�Ǻ����xA,�եcI}a�.�#���! ��\�&�����������1�얝����x~�;�Q��g����ϚI�����T��W����7W/�<�o�k25OB����W��$����å�Ƙ�]0W����E�Ԟ���>,� =�����r⥷�{���w��=���MɊ1C��ў4��j�g�p q'���"�Sa�;S�w�ż3�{�|�Ӑp0b�`����CP1Z9@-���=ڦ�f�@X���6�_?�XW�H� ��F�y�@��,�A�z ���j.��4�/��ۧK���;5�S�IugpLX)�B�J��g��kP- >�ɮU*����A��zG<�n�U���8B�/��������+����9i�\��
Z]��&�+5=rGGX�����a��!gr�L�b��~�m�ض��2�!�tY�?��R����-"�
q��^Ӛ�������UbMJ �'��&��)����"*��t�'x�%!�~��gE���S�<(Nlln�+�����7�
�8&:4d�����~�P�8��Q����Q�V3��u͏d�(��c���q�|�4���_���Pr����bN�7~5N��^lso�s4�d����2�?޶}�#:@j��y��hu.�Ӯ�N<ue��]�����{��MI�Bv
zk��Щ�1�b$!��!z�_�׺쇶r�>���r�����)�H�C���G��9���.%. �d���5`�㈂�w.�{~�����\{0p�\�oGDK�R[���QD�꾧K��#����s(�v���A��~/bU�ƞżL�yI�y���0���ڍq�ow�W}�w�>�xz*�F�>�HLh�G���E�YJ&�˅��^E�'V�w������l3EI��]^�
���ï)�>v��vc��&�k-�}��LcQY�4�woM���<��ƶ�k�&�F����\�}{~��`�h�~�ވZ'^o/Q����1W����Z
.��'�t��{���(C��ò�@}��P_��m����Wv�.��=��.����n�7�^/ݎ���m��#��헲
�^Z������ұ���~Ite����V�>��O�#�	���]{��~�Mk.�Ԣ���L晒�m��m��)�F��q1����T)%�ܲ��.�ee�޲+vs�;�I\���~�����7�}D٪�@L�F+�Ф��k	I��_j�d,�o3@Ѯ�B��߽��g�*�G��Wh�_10kO�V�}|h��RE`xhx�rx������E�|�J���@B/�i��ߴ������E���?������P��N��%�࿾����`����"��w�P�(z�pqX�N���{y�a�ϵq���;��yb3���O܍9t�~*_J�ֈJW�7��?K�+���_�h	Gd�n-��V(�	�F���$S;I�0E�UBW	�|�>�<�-��6�Z���@z9�Z͙�l��ȹ)Jva�7���⫠�=	�)�+�I[��I�Z"�a��s�CEy�.{�V��8�#
���.���O�=�=�,�l\A�}�S]B��k��Ժ���B1�JR�IϢ],����:��b����+$(�܊?z�*EĄ5?E��P�K���o��G3sT���t5L���o�������AtطĴ�������7W?���8yBq� YZ�d���s��btja�����/��r�g�v#�f��DzT��_�F�F�F�\7���Z*��d;���UX��\AK��r��I�f��&M��/��ڬNԖ���Z�`�\`;,θ1��*�X��@oh��Xc�s��_90��WfTT�q��
�Y�mO���_��=���4�|�%O\u����d�λ:�Tl�نIZg����W�#Ŀ�#va�#�����zE�������<.А��8��d������k�����E���ɁY��������7{	��]�KC+ߊ�z�S76*-+���"�i���4tR|U�vD2�>�Ȫ�w�>����'kS������M��.�'�>��h3�g�dG�@:r�tL�=t��ã�7�r���xP�oAj�$�pk�]ZB�z��V_U"���WS���oN�c�޻+L���,	�=����Ed����(�(v�Ԕ�Q��#�c�.{GQzΊQ���d�6L�0�XZ45��M���lpõp����' �'c�^[� �@ȣ��:IT�L��.-�~���x�p�%������S迳~�(_�O�94�p�O#���M�li���)@�66�P��+B��<�IF�.�:����F�)��49�Y"")RŖ�|�$_X�ˣ��"xtO��O��}���͕��ޢd�kGh���H�N_e&[�� ��aK:k�v�O����e�qJ��+\i6)=�{��'�a��-*����2�d~eW��-�u��ʗO����W<ʪ��,<�UTRz�]���Y�A �v���	�ޟj�ڨ�Bc���K�}���r��(X*+,�XF�7�|��N�F{�b�ޔL�%��k��n,jȗ�R,����m��b��+�9���Ư�|Z��1L%9�'W'��[Bs����, Q�g����B�y޸P��)_L��5yb��O�Aa<A��~U���"�J�O���[��!����xZ �h$����tR�ͥ~��|�UG��"ǦM^UIi$�D���4���-����5*��5&u'���������Qq��w�fq����T��o���w�A�軋��p ����"Pk`�s�u�5"�æ����N�38�t�&+���G7@χ�&�e.rsy��(���u��e�[wu|�5�{�u��a��{8ֿ�gͰ؞����˽�L������l�(v�V`)=�Z��Y-�����[�uE;�[��W5��,�o��a~,�`|�59;��	l����n����Ba#�G�|��\Dl��6�-f������|�_P:3
��e1�̫�6�c#������������-������0:;
�_c���^s�_�snإ�mSlF�	/>l]��B-�tŃ��c�x�֨2�O탩�����}�z'E��R��j�6)]���S{�?�l�`�,r��f���nVhkT�����*�]����뭑8=jq�ɥ'���o���<�2����,
/i� ��%_�+,�=��I=?��f���l��h\�K�0�;i�!vP�:<'EF��f�����c ��Y0�ͧ�3q�^�	;���� G�&Za#�(�L�2h�}���0sҊ���;���!�gW�kH1�H(��	�$Ŗ=��;�vV=��~[�OS�|K�d��I��UM\���	���f/�cn
&镟��L�V˵��\TΏrק����-��K`*���_Ml[A[�AIq�C�	w�mъ���3�!柃��9ԓ���7`�K%�rӱ���;	�*��ĕm�vkH���t';��ڤa��� <Ï٥��i�(�L��͆uٲ_�Y-XaWO(j�CmQ���J	&���S���&�K�4������: <��O��.����69���k$�X�J�vM�D2^��
�lry��F�f"~�%����c�z��S	�qP�EH �;�s����d?r+��æ����#�U�0N���d�
��e�ks{���#:�q��k��.M!�r��<�|��@
��Fb	;͝����>#'��*x���ρ�v�(����m���3��AG�hV�=6�w����U�����TBl��hO�~�Aw��Q�7u7{�a������%Lr�;��o����昺o��=�3�͉ɘ��M������8Bt�b�}
�^���ӌ�B�J`zb�v����]mU���5xZ�(��k�57M�LӢ�iC����Pw���zU��5��q QyW*Zw�[�;x��-\Qŷ.;s�V�9xO#�	DIj��,^Z�����A�G��������v]��4����5h�~�}�������?&�?��d�{���vզ�x��m�(���?������_�~E5j�N)q�O�4O�g9>����6�?�lBy�{:�+�����)�	���2�]ԇ&+V��%�}�q�@�q�`�`��%����)�U�	3�x�2S­
���0qOK'�>45R�!���=T��!���$�B��yP7��Q�/_�� &�c���b�J!���6L)+���O�}���#m���rnd�{ �SI[v]�����~U�SG�f�(�[ȀV|����7oqSqY�?��2F>��<|9���o�Oy�,���6z�W����G�x�����΢U$�P�-<HloT��2��E��q,��'2t�\ �Cgb=h~�j-L�a�6,y�a{jcCd�d��j
H�#��$`��y�#��H��N����/"��~�4��0�O���_s3�tX�N�\�ȵ�on�'ݙ'$ZX�<Rxj�%�r�K��R�MS�[]�,j�Qߙl�⾵�N�
�{ܮڅN����]���hsp�Q�J��krs%y���0�_Ue���B�Kв��fQ0�,�f��Z�ƕ:�̍�.���^B�9ĀR:=/�������)��gT�3�s��طx0KF��C�t�_���
MD��ZR{�Ō+���b�jIžI��4��l�a5���C����U�۲jH�`�C�q��+E�ޡ7<Δ�%m������ }�JlZ�B��(�կ���׋�_�>�ҎR�w�)6�1l�S^~A��7�=I�����	n��0�oMA�@�����#��cu�S>�d�W�	�
>���R+���B��+�%�:+^����0����$����O�[��(��Ol؆ ��s�1�U��t�����Z�h���)�����ك'c)t�	QPyli
���h�C@��P(�Q���9G�5�x����?�����P{�P�M��ĵ1�ω�	즷�f�#��穃0�}��_`	˩�^%������S�ѭ�x}��n�\@��w����*���wʥ"D�`��s"�����l?�9.mR2f���O+�@���/\�P�W��"z�P�/����Ba^<�<;w�cҽ��Y4��kK0��ʬ�E}a��"8����͑�E�P���`�/�v�|��g�J�@���;nxv���a�H��YP��?��L�@ǪO����JP�SoŨ����@���愲f=��g�����d�6 ���׸����޻\Q�ʙ�o��7���G���k�%�����ehU����E)�kv�7��p��p���m�z������i�Me���T0�4�8u�R�K���6	��2�h2P	ƿ:�L*�y /�"�u-?��w�l�`��7�Ap�|��p��Ҿ ��^�L�m��?���[,��v2,�X0�1_���Y��s8�?79�s�)�P.7Z������G�(_�2��A���i�cݳ��j���.�҉e�*Ļ�]���?+E���}������Rwz,�6"kj����F*���zmc� 7n��'���%�=�������E*a,p;��⿼S�Q��ҵ�ZȎ
V���{��IkR��.�ZffI� m��v�@1|�$J����[K\�l��������ȩbi)��bM���y%F [0,�-���e�/(��&�h��O��@&�eCP�ݰ��-�4B��k	�����Âu��g�8����r�`�Kk8lp��Ί����ł‵�����hn���T��kK_'={&V��T���z[�O8ܥ������D�o{U��y��*E��>�C*���XfO�ٓPMK��y���E�:��Z��%(��=F�`\�KQ5�#g�/���Շ�䶬���%qd�q-i~� �u�bI����x��͒��R��%�WT_21�>��D��}�pv�q�t`_���b�L�k��ઠΦ�k$�5�� _c>!��͘�k(�e�J262�zPt��9V�1�'�1]ǑIē���ѧy�7�g�W��契j��a����'��L�'��ӏ�.���4��i�ʪ��-��̻8D�B	�|K�iP��mS��i>+�F�zf*��V���Y'1~�i|��I�̰c�$��'�^{�~���9�Q�I����`g���wwQ[��{ ���6Oj����S�Ġ�Y݆��9i�Qz`���߱���Urg����F_¹�yָ������~��R�r;l/�,����'���Js��"̆�F�)x��N-��5�(��[�&��`����0k��Cn��/�LC�~��kĎ>�����6��1��q�a�8֮�����o]{:E��}/�2#�>%o��Ж�a��|��}�f�a'�"W#n^�q�G�t��]ܲnA~������`0)���V._�~!f�ux�N�F�gD
�/\�>T�g�U]��o����+��ܣ`�D�	x��h�֔���X}mC�`��Ѯ�Nv��[1�d/<�_�xpF�7|�	��Ll:�6+nZ_F���������m�%�-���Dfu)�;�M�kJ����GQ1_ӌv_�PE[*b�<�K�c�^K�P�U� �&;y�Z?ꟁ��J���#��"�iz�2-6�.���Hޞ~�k�3Xo��ՍJ�^J� ��lm���rp��n�&D�9G�	���{Xx(��Ǯe=�����ӆ{]�[2i����!�	�@g���5�v���t��Ma�~����`�8G����Iz,C5]0��l��s�6���a���/PN�q��T�@�o��Db�M�l�5����Z�NƲV��F�c�EکV3,5�t��Ղ৷ �q�u<~������]T����͡���AG��h�����Yh��#yD�.�s�¦������] ����~��D<�+�u�����d��)\��K�Ƃ2T��x�]t��}�S`�z��s��_�^n���.؃�g�a��P�i�^ؿ.�f�x�T�.��>��Zl�X�ֻ�oF#�D�%+X�oM������i��L��Y�+��p���e�a���ayE��8���=�_�[�j<�[�#��@�n@:E�g
��7K�'hq�SF��=�+�j2��~.5�ܕ��`��
����۝�	V��i�B+��;�\>�ɧ��Kܸa~���s�1[�"��+��7��z@�a�7�!�ڠ-��'$5�@���:�wN�a6�yaѲ��d#�v#A���·��䋍�&e�Q�/��vm�-��9��r ��,ٌ_Dn-�t�^��P`����P�ن4 �4�*I	~�R�'�Va��4�ɳ����^�6VK*�9��">YwK�O�t4u�$���*�ȒG���*hEuJr`��Oh�I����:�RO���q	��p�'��Y_u6��!�u��3$26�<��R+3�a��0�ޜ�f�u�%o��WI��E.��.���W�V�k{��}_�y����a��{�Y�C	�=~�N0�J8�D��pA~����C�����w�����$7W���>$>cg�����^	n8�~��Z���}G���b����;ʅ�ai��$�W[��~�M{dFSD�x��h�u�!�9*s*�D�)��K�������E���M%fb��m�O��g7%`:�������!���Ř���%�����X�0S-o�|��o&*�d���K�]�֮�0}4�5����Ba��>�6�r�cx��X5��c�WA&�.��H��-!J��B�o�%�(\�{�z| Z Y�U�8��zRӱ�)�3ť%�G_ل)��)�]a�v����_��2���֡n��ۑC��#6�4�S�tu�W�0{;�x����10��Yةb";�	)�݀Q����K-� �n=�i��2���������&)k����ў��Y?U�_~=	ҏ�?���HB&;rV��(-'�E[�ȳ\���m��+���v+t ?S�]��n
��,�Ar�/GCl�,iE��T8��ET2�?�G>k����_t/����S�˳��[��fk�x�����7���6�[��㡯F��V݋�_@��.[c�MVOO�[�D�����)�A�)��=���nyR�Ö����h����~�$��o���\�����7
;e�&D���RV9�(�t��}��I�^��l�7:�?�"�k��B��W��P�s�b=]����	z��h��v�Owlb���^�z���a,&<A�Ǹ��ƼGZ)��$���ѯkS���&�UJ�n ����`�Ԓ��9˚�a�M�ޯ�F��bߴG[���J���b���x4{�WE��62�ȥ¤���>��ۍ}�Ak?ڳ���
�O����=�.Z�"�R��Z0hP �*��zז��˫��`Q����Dx`@�#\�̙��"��翚ú~>l����>��'��tSb�^�����l���&G[��o�f��G@?�x��E�o~
����3[f[m�,Wj�+�?,֮�L-$�\�@A���¬���E�-�[��:j8��W@em�Y1���@F������5���ߵ�W��>�(�a���es�uo�b+�>�gt?�@d���Z̬
?�Z���3���*�� Q��ZCE�o ���z�A.�u���b���bx�X���0�F 7K��7ߡ��qq�T��|�f��MN����q�SL�E��@a�G�������`°�y�VshyFi5�66��&��?{���|)��󆘼�in^YD�yv�S�i�6"�/��1*PC�+Fe!�;��-^�����1�/r���Z�|&�w�`�f��R�bl��	UP�p}T�̚�D%ٓ�I��)'�mmmE/L$W\ >�S^/K�?i�E�p,*q���O�ߝ=u�\�%j�6'�����@T���<]���UU k�?��}q�N��Y�H:/J��i�3���ߍ��WkF�������'X�L���
�:9B��G<s��P83��7#��'��K@1��y�g�Q�۳����1�\���r��)��q9f�1'���5I�����e)B�"�>0��WY�!M��rK<4�_�"��B�B�:����7[쯷/�P!/������u�Ч�ArQ!��o����ĝk0ZɁ�8}��K��97W��	6��Wa�܁n[Y�����)���"~��i���Q$8Վ�'�Հ��a�G'������{�	�s����ҩ�%��}��+�	����K{�<�uU��hGwt������Iq�mL2��+hK���z�g�#�ʩnQ��)�A� 6��axA?��؏.���E[3����x	�I;���D�]D 2�ks��cD�ga5���a�,l��2O<y�O���B*П����XP�.@���c�rΚ�oE�'n���%U�dPbcD�A��Q�M,Kf�jFX��G3Ϣi�3$��of�1�7�
�ͷ�s'���g�S��h�f���Ej�Z�6�Q���U���Z����� �+��������6���UY��f1 �IÃ���.d�7ֱ����`��Ϙ-B����ȼ���Y�E�
��pT��+�&O����h��%;������<W6zrǺ��)�?�Oa�|�/�gZ~
7�w ��0�IQ�5�&x2��TB���K��VVp�/�W��N�������s,������wk��vn'^Xѿ#�9���CQ�-�^�5��!o\�:s��k�ێ?y�	6߭~�������@ʄ�I�g������F|3v.1�lY���ܧ��Z�����ͪ4�yV�
�=Ma{p�d��Kmv5��S��b��S��*0�f����[�u�R��Rs�M.w$$���e���屶�_-�M9glS�+ؒ���Hٝ��M��#<G�q��.�`�ud���V�6�:\^;�P^[06o�;h�w����0�
��0۲vz�}�$!�ڂca�*)�jA9"��C�<Dd=(֙����(a<�������; B\m�3 ���	�bW��?���M	d�D��G��I1@O�SmuOB�_b�!͂6֏�;	�ϯ�1��w�x��5����؏)��B�\3�PU(����~���RQ�׭-�P�����L�7E�9XT�.��L��s"ս�9cmP��Dg�y~gm�19*���q��)�������9���7���,J�_X�����&$�n8=)��cm>����h�xyO�X?�voԏ5ag P+�;�!��4K=�i�K� k3!s�\n鎀k/���o[�w4�E�nԿ��jw�%m ��
A��z$*�0"+������d���-����f4"�B�޹�Ia��9���H�?�c/�7�D;4/��@ v�}hQ����&_e
�n�C����b�a�G��a=��P.��q�ZD�44͟��N�����y��=���hy$���� ��:?���5�p�)�eG]�I�F��1eܑ�i#ݼ^;;!��(A����y�jO�#Y 	�(Z��C,G��xyX�-�e����&��_�$���� �Zz��X�[���q��6@>vu�8v4�9�����)����ÿ^�Z{^�ᕌ��V:T}��������,�g��o0�.-�m�]O0�/.Q�`��2����*�qA�:�v�.H
g�� 	�u��]��MU�vbl�D����A_u������Mȶ����'�"]�^<KXv��n��L�h���봳��'�ۯ��B�?���z����<�b�-VjC&���Q�+L�
��W6^:�i�)S��Pm8��ͪº��)�X݌ʪ" 謴��-��`��S�{�qd�����w*y�VJ�i��JWT��w��wk�Ө�������'Ŏ���?c��x�ĭ@{���Q�M^۵ؖ�6y���C 8��g
)o�*�Gr�ꉌƌ
�pm���x0�ĩ�V�w��J��{���Vԯ�Z�fg�	������^��W�	�'ou��|�c�;��a�@Z'Nv����Ѹ��;����*��`���N�A9�d?�n�����Y��氭t��Nr`;U#)�l++��c/�B�h˄��s�Ϡ�tǥ^�Ei��Q��Q�����Ŭ�#�#"�F�ت�M���j�ԗ��I-ԯ;˕�����&��h'o�iD
�}�hOqk�h�CQ�����*P���������"ܒ���j-J`_�m��B�/�d��
�2�'!t"�� �7��2:�����ew/* ة=f�@7K�(mf�ػ-%�$���k�7Z_�2��w����1��3�)���Iqf��}��L@8"y٭�@u�4X�0
¦�5�#��G��l�����Bh��#c*��,��Y����w����^�m3�NAC��H<�6��7?AW+3 �c��[�n@�vn,/�&>�@�ib�����7��v�L��Sx��j�`�6���P2�X}8��V�J*��YmñĴ&��o��s�˖��~~���a���r<��1���a�0��8s���:.u��6��}}C+��U���7-&!�)����|���?9�	��ox$������t~f#�S9Џ�]�	�Y��q<�u�u�ꉊ�^WD�Q��)k��$�@:�U_R��{�^�ɳ + V����|,��Axm��<;Zd�pJ	�?�U�����m�i+j��D�'rL����ʃfu'�2������|;��N��7r��
������X8�� ��p~�UZ�+٢��Tq��H8ޒ��ځ�&r�Z��p@.�ط��V90Xn��-�k �6���� x*<E�q���q�5�U<쩒}����d��_*$Y~e!���_u����s�o?<Vd;��'�}s���7Nі�v����
4�j�N��
G��.���j���8���U��|k3�$H);���F�Yj�#�`r����U�ڴ���̓(���t�\ZM��1�S�����.s��{��)<��#�|Q��~Mm	���=�WE��@�w�4V���D �۬vm��"Uwꑰr[Ñ��֧\��	���<1�t�����>0��EQ��Xj�q�m[�"�8i�(���,���K\���hD�Z�-� �^����K=-������OC��8��Nu���d�@���u(�336`�_:��f�p��G��t�I��%ۘ?́�,�J�� aڂ�aWPI����c���,ni;0��'����+ӷ� T^%��A�$���L�I��Y{\j��/�ʪ���
߶iewGl�MH�*fڊ:��/d�� /_KjD3���řl��5	8f�k�=�8���b�6=^�{-�u&�Ȯ�i6�9��S|I�4�+�!#���q�ī��� �\�,"_
�Ÿd�[7�MF��{�b�#����#��a�0���Y3��O~��	��|�f[�cJqM~N8��)��|B�����A����=5Gt��NL'%o�$��B�%dm��M��?�ά��IZ~�8nS���6����EΘ�([��@�����Gͳ�?(	��87�p������ �yt��<*�s���đ.�.o��U��7�vz�9I���⯑�����:&9��a6h�d?2$���|�/�͉s�>&R� vvI1����N�Í/�G	�����z'4 �;8��ޤ�+��j ��D[d���S6�]��,'ހ���o2Jh�d�7gв���Ձ�s?O��CW�E��ڃV���~�v��� mܴ�R	M��8��hӋm�Y�$T�:�#����#�6u��}kȕ�������_��JTwE&���p����A�j��@S�W�E�W�����F�緒��p%�흕�E��V��?&�Ch�����W8���+�����'ٲ��'OƁhC�W�C�]��R��~�����ڳ*�:bn �X�C�~.�O����:��m ���s�Fh�U���&V�=[E����#���Z��G�D���qߊ� cQ�P��Ӊ��q����i�� �M�Z�A�]�@�um�,6�o�D�B�A��kH���
��'��=�ӷ�6@�,$ࠫ�Do��Wi�����'�&��k΀a>�m6��GU��w�8���~P�=o ��tա(0]�)�ߢ �ݔ��u?��.��u@��8ZX{�����ۄ�M��Cx^>�bKf���[)��è��2�fm\�_��
�xQ��V���Wn���x��j$�ttP%ti��ԁ�����	����`L�.폙GhF0�����|
��>fS�S����Ia!=��h9�.%�*�����w6U��{�X���Kt./���jc�h�(��`���I���	�/��.�����u����>��-;j]��j+(�����јI�\�y&Dੰ��9P�p �� �3����(Carb�қÍ�í����) )%+�y% U2|�����¢�0V~�����|�/����7�����dmmS�KI��=K�a�wXm�V۠��Y��=N�R�-�j8��P��E�c\AX{r+����B��,�XmD�O��O�#k�X��d��V�.�7:�E�-��u��!�~{�Bm	E���r�y��~�V��A���<D���n��7AϬqN3�6�f��ƚ�K6�låo2����Wk"�9�͛�h��!��o�����z(P�#�a>�w(��\�J40��Ч6�o�6â��`��JԴ�|�ˎ�[[AZ\t�K�����K���~J�)c���{��;\��v G���&�D>��s��)��m~to(p)�B�Z�^�ٹ���oܴ3��>�n����&�IZKٵ�&ތ�Q2���VH����`��ߧ}���F���-��9ۃ3��1�)��o2�3��������������V�o�H�g�38�{k��G_t��՝�a�����9��v;7��)ğ= v�E�/��)���|X�Q�s0�9��G��g��V�l�����5�C�,I�	�53�w<ם�Q�^�F���\:��q84GZF8��L��)�lg��ܵ)��V���%��� U�gU�鷢�bF=0Hz��-]���Cۭ�%��IFa�z�!h+%�䳦�jĿ59�)��#|$:��P0��9��v��J%(bb9�" �����< �c��ɟ ���'��'W+ڔL�$����_w{_{>��G�::�x�n/��x����L�d���;���eu	���Q�O�a�>v�s��L�;R���S��D���L�(V�`��'۪c��ؒ�OO%Z�NS���'
��q�a*�Z�x���6�=��˞��Bء�����MȰ��5T�9�es�d�`(L�k�C����B ~��6}-�m�����l��B�@��P��X��W�����~������6;�74GV.�Ǣ�ZKk_S.c_��*������Ⱦ�L�8�D����/{�Æ����ƍ޳rtf`4��wᩳ����[��va͓��v�߻��n��9B�-EQϰ��	_�=�n�i��K'�A��~e!������s���)��QHi0E}�p#�D�u6zZ�&�	;w����|����C?��C�?���VM�g�\/�ڃ��1��PNU��h�S�1P�T�rו��a'�X)s��)@0y�%t��i�F�	��>l�fᵶٚR�-dh�1o�2� �P\�E���K	��!�\�f�����񠱱<�@j�Kg����z�)�4�����"�swg�lj�:����|U<B�6�����>�@�	��'ߡ������FMQ?h���n�PG�V��p}VFf���5ɩ~�hc��R���w��pG�Ԉkb�~E��"i�����u�����{��F�� ��P�4��]�҆m9m�@R�R>�7Ϸ~����
҅3yΟ�z��yG�~����Ǭ�<ˁ���b�]�S�-&��H}V�}����G�����Z�u�g|�,��(㗑ҝ��ޤ|�����s]���������7�c�S����wF�8o2�8s�C�p 
i�OG�ܷ�W�*�@GS$k�K$&c_�a�i� s�g�����=͢{7�Y��m��y�E�o���JKy�h����15��OC!��o_X�t�k��B�r֢�ź~B�#:U�����/nρ�ɀ�� �s���(ٵ�C<����x9d,k�)����\��I��+��E~���WU�Y�hJ�RS�|z:n0x	�]�6#c��D*���ე�>��D7`�R����gmB~�k�|�����$-5�dJ1��xU��n���Q�[^��Gy�A��lÛ�-y�FB�--�ʿR[�7nm(▜�y�L`�$$E��O���ђ���ݳq�[��@}��M��܄�>���q8!�_�n����O��KZ�m���ˏ9�ܚ�M�{�w=����h�u#g��=Il�Ó<7����܁F��ٷ{:�������m�� �XG�i�4 D����q#�C�=�F���3�v���	t�s R�F��6~�b�F���W%�����NԛO�f�_���N��*�i�ۭ�_�ԅ��!鏴u�u�
g�x�,F�lA��SK�mS�cL�RaS�q�MV��@0q�;��@v�p���f�y0��In��l�J���� qT�x	�$F��V@���1�K�ss��fc��@�2�-;T9��S�o�\��Z8@P9�&޸�Y2e�[�����x�Z@�l�pr:�k�K�d$�l�T�
WgT4�F�5��$��}(�=��p����V#/M��~�(��C��L���giPE�3�T��gd�F���M��ֵV>'`�hF{�C콩��|��fOg������<�$#y<����v�H%���T�#^�a�;CW�U^��pq��kZwqK�
F�d�sf�Iv�[�A[�Wn����MSNiP��S��"F\8hZ%���(����3�q��73���fY�gaS썵�W"-�i������P���V����q�X�c�$��P�$�g0lp��`�V����(��*�/~�b�t�����߅���Q�M��q�%�I�Ol&Â�u<�����`��Q,"��$��F��e&ֆ[�12�B�"F��6xe��A��Ĕ�-��WpLC�V�]*�6���FK7ɓX�K����{�`HD�$� p>wZ2�C�0��D2������BI�݋�Q���,]�fl��DJ��P���C��)SO�=���F&G�~���I��6`T���U� �[�m�<g�٨>Fѯ3�0��<2��b�+y�J�L��8��?�"�b>ʉQ+����������g%��n���hS�%�e�5o:F��$��5#y��\��i�d]��IK���S8E^���\��=��L@��� [D<x��]ȴ0d�7y�Q����x��k&v>����)=���?/�}B&{m��&��m	�A܆nN.�f�Q�K�aqC�<DTa��D^��¸|��4�'���ZRz��g�(D=K@6#�1Pw��bL֎&���3*�}�G��q����� �\êh}֥���	vƿ���S�5�����CI�I:��鬲*l�>G�/{��3���k���#������h(�*�w�/H��2|��g�_���o�����H6UWg��AqSzct ��&nQ�Ə��KI�J"��V6��d�� ���#{��T �{L�[Sq\2��55|�"�"c�����Ոk�߇�	8�]"�v;�EP�a�d�~�2��)i��4�Q�u`��eI�t�h-C7���Q��4+�Io���7���1RU���M�Q��|xh�����|Ƿ�س���x-2�. ߾���5˾1<ʖ_g�SJ�[還0ܡ^� {�L��;1@��8�= s�~�&h�~rE��9��k��_q>MʠS��s�`X �<�P
������ī@�`�&G<���֖�B"
G5`3���}�Hσr�2���Wx&��u4IouV��d ��5!8�k�xU��x�Jt�F'�GAP�lt`�"L���`k�N,ޅ�<cD��!�|<c����������7���U����~���@�DA����������9���׍P�T5�+��D�(�ml "B{�OY��?|g��=1?������CR8�,��>���������*>
^�[B�2Q�d~
�t��:JKLc����vT6c�)��|�2Ńr�:�h�Ɋ,���j������T#�	uB�qL���F�o[R�@B��#lO�Y1����EI�r��p��o���S"�B�5%x�t�	��Q���b�d]µ�4{*=ĻƤV@�Ғ��<��+=���i�;��@��a�A�֫��� �(����7�8��%��y�� n�V$������(����~�Ñ?�Ca�Z��*B�Y���s�ŀ�D�gޅ�}�@MC_V���Ɋ Q{Gd?C�C�v�;�a��Q��9T_��')~$&�ϴ�$/vC���Nq�!����4��`��z���jۧn�#h�Sx�bS��}��k���S}��f�ە�����q˚1��AC}Z��EV���	)�]�qp7V�'�5�T���x)b
`B}�Wxg���.���<�Ks�L�Υ�$��Ѳ�c&G��Ňm���!@�i�$$��L\Ws3q�ȵ���m$��Ҹ\A>7S�}5��q������'����3�e*�a���U�$�R`K��X�8�ɀ�%�~��4Mkc�#z�
��At�Oٚ@�T,� ��\�d#�Rԩ��\�є�=�[��LX�K��)<��ʠ���B�Mo҇��~T2-i���ݻH�#?�����I�(��� ��m���F�ݶ=Yձ�o-���o������ɋ�4Z�h�B5�լ��M��	D@�56�Ҋ��+QC���tX���Z�Z�Z�UT��$�b���P�,+�q����|Ͻ����>����s�>�=��s��YX���p_�����[[�pY�����٨�f�+�zK��&�X7_k�jW�t�g�ߒf���+��Hy0�)m��.p~8�p^Iwl�����������	���&\��������B�*���-�{��h�w��6ͼB߸IR)�*�qJEZ�����(�ڔ�$��l��a������I��IU�vAԓH$��(z��a��t���>�/�
���B�����7D�诤�l�!��{�yU�X�f�l��6�ԑ�AD���K�{Gtn*��+���ةi�|����C�b��j���>O�����g�O�^�yoD7�|��I���2o) ���ġ�����7��u@ ����jH�}˥)�=��n6�݅�e�(�{��ib!�u�O�OT�u�-�p3ιZ���Z�l����݃p��|�	K��˻u~_��B��<�q�����x�}�c<4h�=���Si�O���'�p*����:ѱ������8�r�ɣ��ji|����9�����?�5#9<�����>�u(E�>��Lۘߏ��%�K�z#::����������v�������o�w��c>�IS<(`��EE�}�Z4�0:�yt�5��hu�R@�^��HS�q!�ޝ��[���J�D55Lw=Dx���U�=�ɉJ�sV�"����P�蕮o���e|h�q9;�A��v��L ���[�\��g��s1w�aKDwW�|��ğ+������C�1�^dys��, 
Ld�"��>�zh�P�Z����aU�lj Z-�SC�g�>e���@��&7+����p����"\i��s�����o�H������vU�"��OD���S/�p���J9<L���Y��Ӓ�7��&7iV�VI�b���q�^Mo����۟9��`�M�V)�`�H5tK���AԘgY?S�����Q�6{��C>�˔����qr��4�fE�'����Hk�4�>���nr�������y}A�R�¢���"p��k�/R���0���-a��B(ʺ�
���kĉۏ�dO4?jh�n��_���=���6>�87����b��kx��z���>f�=�5Lz?� ֵ"��$5�ye�?sE��\�,a�s��a��jM��J�_�4g��4���ct�P��L��Y��g ��3U��P)Y�/�o[��j�Ȟ��ɞQ��#�e���8d� >S���/�6����Ĵ�$��N_�*[�__#+۱U�����jf�.1L3��Sht5���K��dJ>���3�ET)-"��}
��Z�fΠݸ�4��#����[�}�D�>W�{�M�gQ��K��������I�0��܌ޏ��͘��Cл�R��F��[�yq��m�Ni;iÈ��"�c�u�z	���؎%j��Z�oLy��ȴ�g�����������͟�I�N�C�@�ƅl��H-|a�Q����"N����k�;�h�Ic���+j�mD��૲"�>#F�|"��u��?/8��]��E�{�j�y����(���FX�4Л���'��mzPU�ǩ
 �Q�B��öׇ�X7=���Ȉ����kl~�W�Q�����\��]J]��q���Y=���%�S
`��O0�a�[�Xz7`��sFF������,����uI*I�\k�sN���wiL`�ΦQbmR�Q��<
�[�|��?���xW76��6���D_�/H��0d�!Z�H�<�H�L��^�W�uE�u�Yp�6���s�b5��?@��T�[��^���4���O������%OS�f䩡�B�.��{'. Ⱦp$n.�U�^R�!0�i�;�9������/�F�װ�f���b $ز7Ӛ����Eq��>�KN��F�!,s�)U8ヸ�����a����Vߎ��Ս����]+�@�X�������8�XX�T9˃v���-���pxJ�?	�x�#HR����uᵃ��rP&A���Ã>Ako\�?_�w�5q�w��Ql�u�j��O4y�?�!�m&�k��Z��_������3K��$�ez��߶1���l�ɏ�u�&����mW�����J=�!E��d.��Zy������8�`1�o��[@#�ǕY���0�������;��3������G6 ���.y�Q�ii�)/H���e���C�3�э���!�����f��>U�E��|^�W��,Z��}�'ӳZ˟�Rk���4�V����'�'e���7�} �f�fפI�qoӚx�9���Gc VS@`�ϱ?���?>gύ�F{n�z'97�Α�ɵ[o���o�����s�1ۭ	_1�f�h^�)�O;�N�DѦR�HSh���RSڬм��l�o�i���4k����.� #M(c]���eSL���$��y�)���hR�4�=�{?��?D�6dk������7� ��yP�ŃY��<��p�9'Z��ˋX�Qi8k��ǜ���cⱆ�?���'�)]�0��R�.��Y���n=k�O��Ƨ�)V�]����r�PI�z���k��
r}#� g�Q�m�pÀ��yW���_��_M����Z�>E���F[��4+OV�Y'waX�p���AH;D:�$���_
�o����ȴ���$^�U��u�3�p�����_(~��67��e`��ރ��S5ك�X�������$0layzc�m�s5�� :��%ɣmֶ;�r���#��һN���:���7���i�S�L����͏����=8h�dkH*~�k����/'���1�:�Ȕ��E��ٜ���f&3�s�|�	�u<�A��8#j�����P�L&�-vGMޕ��,���*���qM�r�a�\�,��&v�-?�Jd�XT�����<C>�)��	�����7��=���_��zH��[I��Fz ���H�;S]7*��7�jS��2r�R��$�k�3�p�=���8}wIs��CD�<r>C�.�Ǜ�z-xw���V[�϶X~z˜Y,�Rms�5ú���
�ы/�p�3�u3�ݣ��vw��41#���̜�߁ӀA���9��5����V�e�@��O	'���mkٵ��߳��3I	�A�tJԙ¿N�wsR1����)���uX�F��g����i�P��]e4%��jw��Y+}�a��e�эVZ-�=2I	nm��WD+�v"j4��ѫ����X1�qs�5����Ńy�n�sPZ�5ѹK��<�����Y��OFrC|��62j3�{�"R/w��v)d��UY��v�;XvK�Ď������x�k0	�m3�T�z��M����ˈ�6z<�[��+吶��?)b�bk�Y�Y�/0��"9UZm�����>�Ь�e����aާ�nQ�w�ơ3֢��x�Z�f?L5�4�XI����t#S���fEq������'W�S�
;2g�<fn�ctz�nq��5^��e�ݎT1̟kv��wus}y�O�(�h��u��>ޝdf�����5}l�����Q�',"s���_����V%w��'�Hx�(Ĵ���C��iQ������'�-wX�w��?q y����2�)7�(�=�,��J��:@��)��*��>�/y}��D��!nuU�p@-/�x����Z&¹`�V-�����M2���� ��?��\9S�}��T�8�bt�h	�rn� et%zǱ���%����`$��Áa�?��܁׋Qn#��A�p�:筞D�-�*щZ���)А��b��ʝ#��q�:�uކ�/p�C]�#l���u�{��F�]�LZ3r��P��А#ϯ��~�cpj���= �h�t[<�Y��(��V׶C%<J���f8#J�ym\,��N,�r���;���ܸ���"h�Y��b� "��'Q��c�n[���O����s��H������PRbx����zһcE��p�fum�/�I�/N�]ӊE�y�K�0�p{�/�/7qR��G�-���y}�Ws8Q�P�|��"�$�U�0�8Ӹ�٩��_��s-��/$j������ϋH�jObv��'¨�G��������i_�G������9�9a6텙��ͪ�p��,�Þ��k�������?�kV����o���e���p>�Bg����}��' ������&��p_"�k�9���$�7���9eO����AvY�8��@�J��{��g#�_ŷhy��/a��wY$xa-.��C�`zv��N.kUҐ�߲>��g�����D'W>"�&p���N��W~����y��L����w�gNx���7��6S��|�^w�X�"���C���si�/�kk��8��8{�M)�V��U��Uڲ�~X�nf7����"��UC%�� Wr3Z�dY�m���������=^x�!0@�L ]!	��E��b5�2�����=�D=��_r����e<uyD^��	q�)���'���P�y�ay�Z�#HA��Գ��kǠ�<F��*�Fy��P�MM�d^A��b��p��?�-A<�n��<(�+���
�F�6���Ĝ"��ӮQ �q"?��F���U�F�.���jV9�U�>\�Mқ����<`7|��|��Ĝ�Y_87�7�>G}��Ā��#�3�a���5��}�����M��&%�9x���,
*�f�d� ������M1kz$���2�8�_Tn��⦿c;� �$6��d�ؿ��z�SE��3�\E˷5���擨8q�h>�8�R[�ZD?��{ʭ���@%j)Z��0�ߊ�+H���Q�VmGO"z��͉Rۏ�ދ������G���[��H�3_���##
6� *�9f�P}s�1��Q�g'U�n%;h�F[p G]�ssp%SޖNԇ���Y�4��@5���n���<5B�*6���H8�E���D "��3��5��+�<�3֢�XK-%����}(?Þ���ޓ���F���Q�iJgb�.}E|�;��'2�1X�"%���R���R7D��9��O� �Vc�~�	Yd#j��\!da��R��>$Q;�u�hJPN��/����$:a:-��X��\.SsԲ;ӧ��1MK����c�<��ħպ�/'m�=�gr_@{���c�6��E��A�̋T���\�1 8_C�6�AR��L���w˱µ�v]�v]�v]#��7���v���cI�'m�O�So�>m;�ʚ��V|��Ю�fD.���Y�'kL������i��vXJ�8F	e���Vd�~6��
M�PQ8*�S�i��q�ƞ_�I$�����'��
�� ����Y��N�\���Pi��۱W*��
�Z�ܕ���������t�)u���b`�F$e\���|�����/wf	�"��`}5c��g�y\oy��Q4@w5>�,�Gi5[r��w��<.K��$��5�VƜv?����V�ΰž��<_dZ�u]э�rc�UI����k�����ֆ�TaMڈ�����YIKH���d�m=ŉ�7Z���Ҝ\��7'���F�s
 dw4�bф��O����Q�:6�v�v�7��n�>�q(R�o/�l!�ώ=8���n������R9��Ǒ%[���};�4a���4]=b������Wr�OH=�3�#j)c��;����wJ76t��m�t����-�.���}��	��B]�@���Ӆ�7åUp(�Y������N���)�j0�5����z�VP�Vll���VWFX�����VC]�S�0c�!��k<�4)�o���r1m�7�AD)��"��y� I��"W�i��|�L�`jy#�(i��/�"
�LZ����J���]q�������W�� .0$� '��f� ���]�Gm{��L�Ц���!�b�:K3�_O��ϙ2��&�dVCs�K���DN)��.�ܟT����?�d�s�r�jxh�{��̔��g��0ߦUooG�T�ޝ%b�
�Ȟ�7${���A�wr�3��7b��hk��:B%
�M�ʇ�ֆ_�4�;�mǾ�^��F��b]g�9�'|�W��V�+{�����>ѧ���.���_X��� �,�p�n�G��,YEV�]1յ���Q���T�hUN U?���P�.��S�>���~�6wJ,�Ei"	=�֑(.���א���j�.q��Of h�ǚ0��I;�rK���2*NB
��b��yN��[-S�"7a`�qXz�;Gu����P��<<c��ꟷ/�r����i��L���y;��X�Rd�"�4cM�b5˩����Ld����-���,��_
E�����s2��=\��"��*�c^���06p�X>����C����\P���R�c���M)�hK��mh�I��!2hs�s�^$fꤷ����ڷ��P� Q�9G�Y��H��T:Y�dk�Jn�8Z����ڎ�»�� V	�WWou���e�N�t��d�����0Rg�Ǚ$gc��*����w�EgA�U��ry2��vz�6YC�%̈́GS���|n��Fd��?��!hb�Y�#���}F}鈝�~���^�E�Jp�,�%^é޶J�_����+-rr7zb�R�R����&f�N�Q��K�B�i�uCs�FU�L]+�Y��&�R�$<o�0�c�i�]�O-�Wz�"ͩ��ď*6��n�"����$̶^�z���0�0���@Oܡn[gP��y+8��/��w9�ݗ�Լ]�q���9��g�f�����CZê��;���D�c0�i��&�4�����n��i;�ܔz���N�g��m���Nk��n����N{��:i�c(2ˋ#U����<�$!�{�9�����|�%feqē�:Hc����H�o�籩Ԉ���/-���F�q��m�'��Z�U�r/IXwn�'Ҟ[cqVi���ٓ�H=ɲ�K��Q��\d�<k>^����8�-�&-���b��A��D���%�YD�}@���s�p�9�x~�N��o��,�:��ƌ)QZ�<t��t��?���(n/�t�����l�f�.
U�,����G�@�U������$<�_���s8�$֓�t��_���kfq���l������$�__�5ĝ<�����V���*TG�X�	Ob���S܂Q/+.i����3L���/�:p�'�=����-����-n~�u���W�F䉟�F�ۇxL_|��hd�v����J��=4���#�������4QD��*ToO�EҊ];T��NQ�:�����*���	Dj��K9`ugp7���M�<���̰��Y��aֻA�uZ_����<چ��#���n�e���?�2��"�L�Z}��vkem��kz$ĥH�d[�u�	��Z�\&7��� ��`�T3r�D�."C�+J#eG�֖}g*�o�+ß��(�dm5��W����\Ħ[#F(2��9�����Jc��E���y' rO�����$8�xə���K9��G�b�:��2�ʤo�����j�����>��*�0h�=�;���`k���!Ә]���w���i2`r
���o�"@��
N�Q# Ԁb��G߂�|� ^+N�c�~���i��U�Ñ氛�����Fۺ�)�q�yܓ�՟Ô7�����z\�r`�[����hzv=�Ӂ��x��e�@�G��g�f�o���RM\�z0 txl�I������?�3^Z��&�I�����b(��BE�f��E��-�hY�B���5������z��1�]�z��TgzBՀ�`; �������`|��v�uT�枇#���'����"��ܫ�45S���֥��;��L�3�i��Ѵ/~/=��YO���-T0�8�q�l�X�5���$?���T���r�K�к���:�j�~���@�d��m/��k�b�� ��f�r�<)#[<�����r�_��t}������_�!z�KRC��}Y��	�qDt��{	���� ��;����$o"��������k|��T�v.�kE�Q���s��]��41�L����O�k�xl
�\3����K��GµO�� y,�?X�+{/�iψ!����L�J���Dj�h���z��ݛ��>����R_01ϧVv7Ԣ�������Ka�غ��G���M/���M���?�°��B�`�E�Ő�uҲif NB]W����6f>2Da��H�)����!JrIJm"2f�AX?��_%]���P�(h_���g�b�*������9
��Q[�7蹻)q16�O]*4����Dd?~K���*{��5�Gr���֖t�[�e��LSgK	5��"�b�}���i��c0�Bo&f�|m㥙K���͙lC�^x�r&^��f��$���(,���IWn��rz�����{�w<c�!j\���[_�X.�v�c��L��d;��h���p�-���]��niQ��	A͂[��ɹ� ��r�ld
9d�(�vv�}p�#_�ì��V��)F�J�9����AbAb8�"[�'n!i���@�*���00��oK����t
�~���8n|�T���u�8�kf^9�Y��p��f��u(����=�6�I>8A��,�S�h|G�ס0�Sm�f;��V�A\k[]O1������6X,8[��8�Y~LIҝZ�5����ϒ��j�2K$���N�5t?h���vp��p� �
PS�l�hu��1q|*��Yd��E��-{2-�ɕ�VC[��x�ЍYM��ݙ֯��)��`?����|3�����HUgS�P�'���Z�nt���)��P-�k[#^O��M<�PW�r��;��tz��C��Pw!	�S8{����+H�� zd��qE��yɕ=/�^Odf���e��������Yq+��g��W�����v�����c�'gB�:d���q�<�H_W�%��Z@�d�_����26F��Û��1{(H�d=2�/�16�1�O��J�٨��ΆY�L�*J�s�����O��=���α�:c��@�2�2����!H-BR��V�E�fZ�7&��k�'5V����1R���m��AgY��*"��ð���z�~����G4n/Fw�9�8���c!���J�;a������E�r�u��N���~�nN��$��$0�da�����4����B#��g?�0���=�H�8�����q�#��څ^�p`gw3������	�n�u�2�ۛi{����K�	��{tf�~ztR�LT<��X*�>|J�D=�v ����,�X�>*�nű��q�s�-���Ud��-Å�l�;<�C����a1����yϦ�~$h�и��������ɏƥ�z��Z`eȫEV�qUc�Wu�g����?��	Zo�-�ï�K`��F��#|�#��/�\)<�f6���I���q\O![x�.����B�e�u�Tl~C�W5��3q�4����b�E��:�dC�ȁK��^�_
?AH*v^"�z���گ��A�jzd�%n�|���UZ�R��*���
��H�^/��ؗ���λ*k7a��p0-�J��k�o&�u��h,��K۬|��Wyԏɚ����;; L��\C�3xP����)��}T�T���M����5�&�8���f�=�'��Fn�+cr��h?��Ƴp.PW!��aλ�t�F��k�N-��B)�;N��=T�:�|�����`�� �o�o%��ڧxu����)��nݸ��gV���-]�o��c�W���y
O��d��4v���в>;"�N�J����3�^�K�.�U?�O��W�j�������%�l�Oa��t�1��~Hj�����Y����5�q����t�����i����#�탖y\��#�e,W0pu�A��X�D��tµ9��R�Is��R��� �t���{&�g+֌�ᔙhnG�)�J�x8�@�u�ߚ�#s�Y?��k��`R��0��L�*q �����fɍ�r���촭����5釃v%�r�K�'z=�M�'|B=C��R׎��2s���Ds�9����e��ܮ����_��H�� �kCRr������$���p���d��Vn�ӻ5��w�T�KHT�~'�6���㢗s��˴W��7��j�j�\�cd��F7J�!˄/����Ӫ��;h�-�o%���34��-э�u}	���]�p�l`m��o	x����=d��y��!(�	�-���D���(i�D�}��5�tכ�c7�	U'-�������>�H��Ȉ�H3����w2��.?+�4ـI���",/n%��4�|����7���@���L����q��B]��9�^aW >��I���PM��5���x��ӱ��X�űX��O�����j�Gצ+��l�#�A"����?)Y�>K�	��_S��:��(%�Ւ������� O�)��W��A|�s���;캬�/�O�C	��r�PM)�g>%�[�M�� ��D脺j,<�Qp��3S��4��i��־?6�$�f�����ndep̲kK��'��r����Xyؖ����K���~Ṡ��dG�����h�D��f9����L�Z_斪�%�2�k/��8zM�ƙIX��.>h����Z�=,4�E���[�WR.7@.Ě�[鰃�E�#��&)��?Ӗ/K�����H�(��YE�
)�ZK2�L)�!D�S�Ȉ j�dR�>�OF�\� �2��X��)�Q���67�/�����ƞ㬟��%͖�3`�<E�I��O�K�pdA?I~$S���'yI5j'��쯕Ag�}Q���u�M��sRk���gMO5p*q�`c��0ɳd�yQ���Q���P#xy�A?�
��Ygc�&*	tQ5⋺9�X����b�!7���ٹ�·��l��5�~,ɨ5���T2��E��F�E3��c^)�z�w�Bލf�<��Y5��V�g�P���ݼ5_]�<i%`F�����ߺ"!�a��k*Y�㕉��H4mdW9aZ�'�W�.,y�S�?�pK��I�.��k��z"c�G���-��0Rd|�'ļ`��C���0:^=����r�V!J�Y�������,���,H�(�jf�$L��ͷ��k��7 �o9`)��d���CP���O���^sIqy��a�����ڝDRK��� kư����m/�W���m�9�c�zS]��e�-�Ȉ���ޭ�����.�䘚s0	#)q��^$��(��iV����w��x���W�;oS>�<�v��É�0�����cHڏl��|Z�<�Z$�T[Զ#�o�O� �Wє�����ݼ1_�3Ӎ�8#5ݗo���S���@�
�V�"��
M�Z�?�����;L�k��oa�߄�>?����|�,�:�:��qˡ55��\$9�}ۜ�fQ�w��k�]4��i������Z6�|F��C8�hď�~^���o�&}º����q�n���yՍ��ܒ��Qo�J�V���W,�3�4�,Ϙ�l������'�TW��$�(|��ડ��P]S��y�專5�;^���?Yb[0��Od��ň�;l�{:�D	�eQbtb"#X%S��%����<ifǂ��V�թ�J��k1�(��Y��-�(�k{�珃�_��l��6����̑�k����yV.�b�~�Ȝ��o�v#c��j��"�3d�e�E�I�ch<�{c��J�P#̺����~��Py�#4l�0��R�en�L���厓y��!�`G����5������P���,5�����hfwk���?��$�M�#��5�?t>~ӯ��^ş�>�a���q.Xg��M����N�%�-��w�	���;��%�:w�yjx��O���2E.�|��z�=	�1��4a�;���t ��,yG����d t,����O_��`�X�z��b�Gݸ���������h��%ݱጾ�Q�:�T�LU'"}���������"��f�����~7��`3ܵ_a��֘S��[�F��f~�-{�\�����<ȷ_i�'���*��y0Q^��W�K��t�J��,iF{G�]�5��ǁ�-��+M_�x���2�PYJ��k�3&���"3Ml�s��ȃDy	j��H�Ʃ�rc'�a�w(�큯�IY��p{8��V�`l
��Ǿ.Sng�:�@���pA�c�8N���ړ�?B��Dp�D/�q�Q7?<b���(�� �x�mh��fV!B�Y[�s�7c[��Vcu���	��U->��zc�a��j�f���rN���J���0�!~�g�}94���5��1T��e����Ӵ���3İ,ɭ4n-�*�욮x�K���4��m��֘�D�u��HX�m�4����������*�����e��tf�����v*�g~���s�����*�x&��}tD�<2�7�NB0Y/���X����7q]�2�U&�mqb��?an[|��+3?F+��>��O*?ݵ��~��eҽ��p��ן٦�I���a��~��?��O�1�fsd��Fi4�8Q�V�}Y`X�x��Vp_xV�d$A"��?�"�]�F6��dZ��To�>���7a�8��tKg?�i��� fc�ޝA��6�:s�4X�g8�J�M�*����x��Q��އRP�h��@�/����~Z��ʢ�_n�/�/�D*GY�O�n�Sϲ~�vC9�4R# ��4E�[�O�6K�[k�/�>�\lh��B;��ڊ�n`2h%ݖg��k��tdx"� ,�8U�J����;�d-v�mQ�Ċ_���u3:
���0G���������gB�:�j������=�)`FoN��8j?�����5;�/��#���̈́���`��"� �=�#�Zyă|ӧє�,Kp�����\�,#0Ў�N�W�_�)NV
��[8]��z�|O'����18���+�n�����r��g2�F/Yd�v�De�{��6D�hĹ�x � R�K>�;��uj$k�]��n)�O�U�5�P��G��U��	�����:丫�
�%jm�&m?=�Ǔ}����ze�vW�W������͇,�e�����@��oM���2ت�XrJ]u��8�O7�FIs�[���y,f¸���f�IM�����>�d�#�"�<��p��CV�B���(����=��ן�p�xE]u>�o�9IxR^sj2��:�ǄH� �E-������vl��l���>�Q��y"2W�.x��:��k%F��̀-*���;���vc���>FK*z�	5Ʀ7B�J����?K�xb�j�V.9���s�8U�\AvD�3�����I�_e���xܢ7H�⅘��b��蔔>*�6�$�D�?"J�Ӎ�V'�����襒�_d���>���&4v@�t'':�����dgrd�z��J���}	�d����Y�_�����e+M�э>�������>6�C���U����W�Ee�Bރ���tp�
�j�3ߘ����2�@�8���B�
�{1��*���2�$��B8�<�WO��_�5�i5]�If&}ǯ�7��⤣E3��T�A�x�3����O7�-q�^��~�vL�Tc�L@qm�׼���j��];3) �r{��5��C�.�E&S�3��e&F��&#����SJ�1�I:��I>-�m�6g�"�8O7kHx�S��c����1���'�3�{\;��
5s⇤���hSc�#�f.qj�%yK�b������s��g�67a���]�B1aI^�m��+�R�tO��E�u���)7��m�z%(�z���	!��J#��6>פ*u�' ����@��&l~���1��]�w0K��Ho_@{��5�fJ�ce�i�v5�>�O��b6�t���ex�iU쭨���hS��D~b.,,݈�N�Ȋ3�QM�jN[O���j;��a�ժ�Ӎ�Z�<��sI��R���8����İ��I3ʪ���I�&��v��Ϣe���%k�S���>�]����Ү�35����ֳo��(���	{|"�'k����L��\-�r�z�_An�k���H�|B0tӝO���t��<I�-�L�j� %�85��3�h�ʊRiQ��3,<�$bQ���^�$����Y� b����[چ�T�L-�# H���wӷ2H�a�\\�i���1{�4=�t���Y�xv1�n�2e5 ��ON8�_y<Z��~&�#Q���,[�wZ}G��
N0)�g��ŠҼ��mӝg��fHt \+$�Ȣ���pJ�	�ލԗ�<�dgpo^�+B�f���	�[�Ŀ�O�_�Z�jG��lR�ɏ@�fc��j(���[z�V�F��fG�]Y@@��m������c���u�ȫ��*���K�^�;<��mA�!��9 [�g.�Ź��=��q����3n%n�p��.�����g�-b��o8�{����p�fl��~$��V�w*C�̲蒤��/�N?',���/s��ĀyT��v�p������O�)^�Wj�+���<��?�J���Hͬ���`O������`q0��k[���.!�K]��Z�-�V�s���%[ġd�:đ����rG�zn����f��\���4>Ujh&��LXB�Fu��za�З��C�t�T�s�!�4�Ҟ���C��mՖm�s (���˺W�b�we۹;h?��dW8���N�oVmv����[��O���F\(��X��"���f�MҞ�f���?��M�O9�9'��{���9xV3mq��{k�ƾa���ߵ���i�\`u$0A7��J����'��M��S��E����Ч�Ч>`Aa7C��В�}�#p�W�1/����,EH�����LJ"��f�,�]
�R8c��x�5���K��i'��?L~�����U{&�)PW�`�f�Ϝ���s`!��jtslxʟ~���C���_o��nE^ �ۨ�mY��0�G�ƀU0�Q�hid�dE1}��0}��s �^���&��6]E���n� ���~�_�-)�lpu�WF��&֜�[�e�~-��N� k��~N��2Tnz�3d��z(;�!� L�N�הV8����;�k��X�#Y9pW�c��y>`� �Y�7�$����sT�c�n�BQã���y�u�F��8b|��skbcSuYO�U�su���r�617$9)"�l8�(h�R�J7��N�����@dq�^�ۻ}
0$b��Y��X9v��[1�	�v3<Ek�j��T4i+�*���p��>\1LTB5dDG"���K$��_ _�N4үr�]4RO���B/)�(�%:�;8��n��\�2���1����Y��x@��Wێl���O+yb��t��j�_��w���jp���ۓ�e-��X�G��U�ƀWV����E�^6��v�	��U⑑Q��.�*���E��������ж9��Â3�h�gP~�c��!�Լ�A��"�T#�)�Q�����j��n�41�zmWIs�����i����S�W�h��;���p���:=���~Q�*N�W�%8� �=sԣSҥ�+^,i���S�̛�u����|�wk濘ے�īNk���;P��JD~F����W��NtT��*���
�i������&������.}��Uͼ}4��;v	�g�>�����6nIoG
��Ep}K���nc�ϋe�+{�ڗuo����A�*��š2]6ܨ���N�SpG8������վ�yI�h�f���bn�[�e���`�>(w3��k���Bg�C�q����<R���#�x��v�� w2��E%z�'�q�XcNf�NA�?��ί����Jk���������kޅ�P^sR'|��x���É�섬C��S��E$������0���T�����{�:Ζ�溷P��������	2A+�K����TdD��q��kMO��I�'ɵii���oT��ߟ�����9>˜T�E�b{�Y��;ɨ-�ӊ<%]981�'%�_k��S�x����]��W�q)N�
�[���S���$A}h'�VbqM*Vi-ٯ��jٛ!�m��������f��s�#�E�q�&�Y�����1���[���׷�'?���R�G�%�i�e��M9��m�<��ʔ��գ��-d!ه�Oa�����a&���A����N��^���\T�#�k!nm��X��A�B�m��55!��V�Q���F6��_ N=/���|� F^I����sj��)�4�7�����#�I*�5�NH�'��r�i�u(���>c��^>�_z^N���q��
�����{"�p/��sQ_B7��$G�zex�$qG��b5l�Ex����L��d�
�B]�/�t#��M�Y��[ցٌ�O͟*�����F���̺غ�#��m�:����o��V�5�Tə�\�21���G4e���w�F���<T��e4��vأf\�+w�Fч��#e{�+�U	�ӿ���VU�v�*-�,:��@]%������TM�{�ÿ�sg����O,|.�#��6>L��x� G��v�-����L�W3�6{�2��uup��cϩ��ѿԣ��jx
l�=Y�j��K[����FF5Q�ߩ��3�X����#i�C��0��"�����O߿��5aNql�m�DKU�u�^XLM��U���k$m�oe�o+q��"��iv#�%��fL��j�S�d{9�j�׼��1�i���W��f��'�\�)$ .b��|F7�|Ί�;�[��_=Ǣ�4'��d��a'|����n91!�\u��y�����gq�M����V��S�Q�Z�������g)�*�X�09_�Q�&����2��!��uڹ�c��9��(+�u�X�ȩ��`�]��f���kМ��8��k�=G��(��.M"�w�!E����!�C<<��<�X�fYiX���;p�T��~5�M�޶:HՕ0�$@�!�4\��N�-)��j!�$s��g;&IG5V���]Oģ ��UV�����	-4j�D���u����WG�[TI�rG�|F�����^Q���Oռ#��p6l*�J߿���7���5s(X"�s�Ά�U���R�9�}�w��xiAI�w�(��Ĩ�cz{ܤ"}��b��F�ɇ�ϋ��)4liQ�`�����.l��SH��U;����T�?D��M�{��b����Oi�cRklPY�JY}����.5�)��Wp~��WKF.����Q��5�!~J��
E7�!����4�L�ͻY�^���������P��:���%]���'LPh]���]*��Y����"k�8YXX ���H��4�~�t.�F�������E7�XZ�O}���U�u���he8��OV�w��*\ l�Y���<����$����(��z�T���x{o��[��}Itk�#��l����p�M��Yz��V~ʄ8K�5M�5�b�j����J����P˛�B�FS��K��%]�m��Mz�t�&���iT/>��3N���h����w@��e�5삖��@O���VD����x�4e���؞;j8�ň+|�Ʃ��1��!$�:�%}�����{��Ō�zi�=D�@�ˊ�(�rAb���L��C���Â$����;��O$RP9�bpI����Yᬄ����"DjH����E4�?��"�Hl����\��>*v�9_�C�������J��K�q����$�Il�)�I\�څi��S�����arQ�|O�/XG� ���z�$>&O�)>k��ejNr�������fMLP��n>	\����Dj��09����Oh���p��`�J״���^��~y֍I��4�!����H7rR:��޷�`t�a�;����Vi:h'< O����)
�����,6�~�c�FS�ּ?����/0��n�H��9_��$xS�K괴E��i׶��cʼ�b�
wk�r���yl���9��}���ff#�0���7��� k��"�z�9�h��PD�ǈw���1'��T�U7�4<z��A��0KQY]�	g�*��K2�g���ͱ�I��
�A/�䉸���.w�R3��ͼ5�*:3."v������v��i#�,~?D�V�T���H����Իj��!�[�-�ۆ�u,����.W_k��_����)8�\��3���â���P�$��K����:�(��y�ho���ΰ'ወhk���k �}�޼Ʀ�-r�O7)��G��8$z��&L��pwv��8�,��ѕ�ѿV��kMiM����}z�8��opT7�P�'��ɶ�αa;���Йj'
�q�ۊ�!�f�=g�N��t���'��x	@�
#g��ӹ9$���4�Y9N��������ގ���� �����3L�t�dhU/�E}�V��C�q1e�t3/��,_$�O�,����=���h�25�V������d4����V�zO�t堋#�7�-/=��ݬ��������Io2=�b�S�(�o��)	0�=C�����eȜ�o1�1�}���#o8�Y	nJS�U$B��H��	��x�|¡�_d�5'��[��V'W��bE��m��xPn�K�O�ш,Wg0�|�!"�r��'��k$���?�q�&܈2C������^��?�RN���P�:�v8Dp{�5��&I�(-eo���\�~^M�yp�&މc���)Q��?�'�؜u�i�&����Bp7i�Љ9��y�#L�F���t���sL��R���'.�M�E��1�x���隸�~�o�>%�$� 쎛�/�I?*hjH8�F&�/t�mk�k8Fj/��W(�V;�����8�J�4�֏7:�reJ$���H��Q�?]�%K� �b�õNˣ!5���t4}�=�v�%u�y1��y���F���-�O�/Bq�~��O��\)}r,� ��+zS�V��^gg��Z+n�OpƉps:ђ΍p�����F�17=��~ٓ��ۛ��� �U%6��aX��N�-�]=�=��0���jl�p�����RRh�x�~� V��A����l�	��F���JM٢�הN�H��^�}�3��^Bb]{�w���?FOʲ=~r9��I��0��V%�+AvVW<?zn�A�� ���0rzO��
�_Jl^�V7z�Kl�T��?�݉J0�-�s<��΍'�'�譑�FB*���=%���葭�^�?�X�o2� �xN\��Ļ����Γ�g���7�/��|�W��9�N����1	�N����K6�!z^�<o�Xg��3����D7���4�aN�jٓa]}F*]���5�p��k�B�?�~C-�u�,\�#�����'� ,ُ\\���Х7�
@7�(7�x�oV�r������y�`��y�;��]���
��#��~�?�9�Ns�`�z`D,,7��G��R�dW���:ҜK��Z;�kjq�K��_�At�C��C���΍$O����9���b�ל����$վ-آ��Bi���Nͼ)�^&�F�]�YQ�`�rǸ�ef>Nt-ĖA�;2��o}�Z��h��I�_ix	~�|Ν�e}�ϩ@�p{����x9�˰���7$ߥ������U����3��9���t6���u�ٞ�Iƨ_pS��ף�l6�=����ȑ8fj������+�6�h�ED��6� r�'�Cg۷��!>����Ƞ�Q��	.�oyL`D��Ͼ�5��.�����3���X2�H��;��~{�w�g��^dv͜]P�5v2��-8��ij�Q<����2�C[���*�Y�/7�1�YG��zgj=��+6gtd]��>��F��
ŧc���n�f�Ŀ$	Nd��RD��v4������p3��m��s�E�^sf.D���4>C����S�̙X׹Զ��S����Ѝ�`O"�ϫ�g,��m��Ӹ�F3ZU�E��@�p���,_fu>ZlΨ2HD{]3��Tj,��@̤�_( ��M�̙��:�DaR��|x��q�ei	r��7�|f>�$���*���i���2�
������R��9���9��a�9�Z䯝�e�q���ȝPQ\��_��KK����^��6�Dû>���C��h��,���!Y������	���wyT3ˊ+�/�[:�vFp�o!b�Ġ>�$�VT�<ű���k�P7��֒.f��u���C��g��<���ٺ�ן�x�|��7�� ��/ޚ��4\�yRi�Yq:4Zfw�(��mQ੕5���lM�ݚ^b�4 N�8}�8}Ip�C	\ �?�V�zp�N�Ȱӻ���'��R�&�����G�-u��s .��wE�X4G��K�}ZZN��tT����^ٟ�',-�?+��7�70ؿ\;�9~;������M��,xY6�Qg���5t��9;���Xm�g^Is�]Dr�5�"���B<���P������I8�	�8��XRk8��(�h���ĨM�O6�6[\[Ե� �k�紞2���T7ς��-��L��6�����=b�_D*�aG Gf5e#!����P"�"���|�57;?p0S�.�=��h���܀cJ�1�����V�c����YjhbSID�@ͽ`[7�l.^ĉ�h����x�>r� � �&z� -^�vb�c'Iy.��a�%b�=����b;C�@ �^��
h��'��M�G��k��b�`��*�m�Ɉx�%�;z��\������LWWM`}rH��JQW!)�ka�54��2��9'�kN.���Ҝ����5�c���Z��8��;y�<��=-�g�J����>~�I�n' ��ǵ�)�;�����Q�K����0���e���x��:_��[��B��Z	�࿴�����iD�����]�Z�YS�MB��%یL�C7�f�'Rt5�L�f�k^��>�J�>��a��0�B�u�C���8��-%���n;����2��R�]�5�sؼ;�JGi�v��Z�[7K 4͆@��f��v4���ڠ�2<E�!�(�������"�2����w.7௫��\^ X������?�=5!̬�#a;񤧭��Y&�I'�tz<�]���ӛ��H�z��^�ڞ�>e 6B�3I���q�;v����W�pz��������bWm]0�?���і>F��ծ�\*�Fy5�1�wqhhI��~�c�ϲ�I��P�̫g��̊����6 /?.����1| C$5�hbkoՕ!�jC�8��&��H�m �j��v����8�Y}AI�4s�n��v�i�*��~���Ե�Zd�o��[�u[��[����-t�O^����)��]z�|��8��x�i1c����#����1�C`Λ�2�t��i����?ҵ�����>�);��O���<��I�Q�3���O�pt��a�:��E��x�~���UW-)��I��F
?�%[��FZ�Nym����^ֲ<i�l�+k7��M�����gO�_M�%ѵȴ�����t(���3|n�?O�Rp[�fEV�`���)�4���������|@˴��
��.������np��^�{�k?��$���Z*k�k�߽;��h곭��P��F�n����"�f�f�M,��O	20 SUŮB��`6]dNs�t	|w��R��ࠡ�[�z֪1�A&GqHHy��3�|�6�;D�^�Hv�9�.��$.ĺ�=	���ݷǝ�ԝ:뷸�%� �䱿�&��?����D�v�|����u���+�ڣGT�s\,>���d۽"-�ċ�l�Խ�H�s�{ V
6^Gs�9F��hE���4���!�4���aÀu�T��E-0z�M�'��G<m������0��f��CD��d��c����Ȗ���ň��E�/���;�$� ���6)	��]�$&]}��R���Y��כ|G�WZA���>�c_���*#��w\A���G�7�x�I�H�X�I�<�Vsc_���D�0IQ����$p��(a;��c�x�ێ)�[�(%���D7��!C�3�=zmQ-��H�#w+�Ͽ�����i��2��;������P�\�8
��X.���U8���)��P\�:9ydB �wg�0Z~j��tuj3b��Xp�^d������U�b���}�a��Zc�I�����t��nW�?���:��iVl �.�� �<�&�>lYJe���<�	�"����4S�f7p��k+E����#�SY�� ]�s�&��3;�t��������đ �Y��k�!cL��܇a��2�V#��[j��� ��D��]�K��r#ќ�5�4ַ�<�zb��o.f�f��h�C4�e�D�k���'��b�1ahg�@�$0�f���#e5^s���D38�.˷��C�F�F<�FF?��ّ����9�|��/��8</�$�^���`T�1�/��\1�w��7Y��Ѝm����`<K3g��x�_b�� �=�}e����xm>L�C�r�Qt�[(�SefU�rJ�1|�O��u���F�{��١��J�ԑ��vz�9����^P, ��L"���b9�ۼ��Wn���%��bC���G�U"�v�'3W(V�{d��Y�6��Cm�c2IiH��T�����}�0�:�}.z��.���{"'�\(��>$�4�3��7����,( �T�i��W�V�_��\�7��rG44�<�J�C��f.G�� ��l�-�:��b��K+
���t[��B*���o�n�?ƭ��7�����K�6��~�qND-�,�{<G�%��0�U��sH|׊8�0�\t�9���d?nf���R��^���s`�+�:�u���XݖVƈdu֕��&��{N�(��1{�,�f���6{������c�C�k��O $�9��w�h�_��D��^���T�������t�W][��o���Nu�[���?�d^@ZA�3d7���1�8���|�(+��o��i�z��U7g����MM�ˌW���W�>�'RZ��e���U^������\��k���P��Uǟ���� �e�����u.d��d�{�^��M-Ʉ�(���~>׾)?�Cy3Zi|i���!]C��cC�ņ
���\������F�x�'��H��	�˔��6=q����]8�����%�QY�ӓ��A	�4Q�eM4C&�rt� ⱊ2(��H�v0�x��~^�*�\*�$���b���5�%9�����z�'����?���U�u�zW���ۭ }�07��Sɻo�8}�o��������D�64"V���N���:�/����ϳ�66�����۶�O���|<W�v<��4N>����8݈�H��c�"�*�SӾ}�K����~<��g����S���ۧ�]݅'aLBV;���N�4��� 	H�����w0?8���0��<��m'��y� �R������;�m�I�Z����$�K3����t��V-k��Bd�d�:�Ɓ�XV Ǩ��U\c@v�M�vum)%�`��W�O�u���ZNޛ,��խ�+�ۼ��LH�/0���W���V�G{d��!��\�<BP^6��2X5�(��u��K�����	���;(?�r�l ��r_| ���UB�F��K�^`L��(�V�KP���r�o.�fl ��b�oq-�j�<�2�]�u�ϕtU�ŁQ�
���G�l�C�����22{�A�^-�[��&Þ������d�7�i���<]�N꿂�����x���Ec�����F$��TⱧQD$���;M4��ܘgKp�N1��N���l\u� O�Oe$ZoY����{ri��,U�@Sz��@����c�u�Q����K\��c�h׌�ޘ����V�b=&8�e��|�+�~x$2eø�v�-F/�n����>;�HEn
�̊.�R!>g����9!��nn���iT��&c���?�AtyN7*7p��/I�fډѸ�(&����rI���9:ҝ�}�<�ptt��+sw1�;��eZ�X�Bc���ȃ�(]h��E7��gw]ć�oY�f1�gDyz�pS;�o�}F�Y�7�/�|�� ��iz�Y��QZ�"��~��`�Y��b��6�P�D��{VҌ�G��	��gB�d
x���5y�����Sx��-�mɼ-�c��K�����]�B�a»��?Z���O�<�SIQ��daw����/(�zsy�)��H��V:|�I�CPR�����alة~N��~8Т;�Sy��!]��< �:�פLn����ĥ�ƀN�P[�ÄLV���(���1���A�ŽX����hM�n���Z�[$�t�����>��|�x2�o�!�"b!�ol\+��9
B-[pڶH#Ɠ���)��$��]���1���Rԙk|!qO�8O���M���b�{�Iz��i�K<>,��3��Q��w�	�L�k��Lڮ��2�+�����W)�P�*��Q�esC���`�ƶ�FnI	�~c�N�N|�q���Re����' �}���*�b�OkQ|��wڌ�}���݋l���C����6���ɥ��wq-ڤ��;�8wR$A�M(pg��)����>H�>'���S���5B�{������&��e׷S��c'ˣ�L/��gG|����ż��9��K�aϙJ�p+9�J�< �m�у6椠�@���� K��vJ���%�F�z������^jP؏���n��7dbf�Es=�6�y�� T��G#�U��-�Xީ-��x�{���I�����d�+usWc5u'��o+�79�*�"���ҷИ]�l;k�y2�_f��]�T����8N�pȝ�+�L��\�Fę�3캐���	��,T�sa�P�_���qE�L���*F~_�S�S](>��F����*F�\�V*��dqd'y[�)�j��,��ӒuG��Й���V�ϩTk�w���a�gd5d��ʦ�0Jq%��	i5��	�TYP���ݭ��j x6�����#�1"�۾(�1�9�<����H#���gG�.Fn���&n�F�����,�I��b1x_���b�b���()B�Q^��0�y�#P��?�u� B�h�rr�ӌu8$��/M��'^i�=],��2m`��v� ��d�k��" =�2ŀ*HQ|G$�(Ų)����o��{7#��\��s�5�A��������x�D܁\+r^�N�͘�#v�.���]�� trJ0�k�e���T	v+hF��Cڍ�	�D�A��~ŭ�~>>�T�砟���g���c���n&�,�v�*x��)�)�e��$}pvC�b��S���V���C0��0���r�)a��|�~�D�j�=�cH'[d�>�ѣ�!�g΅�C�9��Fa0����?����!밴\l� %�H@��Rw������.
�x�3�:���:H@�5vr��>y����Xʆ��+��ӟ�+j�)~�.20�`2�<`v��0g�R8��)#�)�����a>Ə%4W%�bܬ]�?"�B�؁��f	�y)ї��O����������Km\!�I2_�l��d��Y1�˦�a=Bjg���/��"R�1�Iv�'0|���=z��` �*�ŏ����A�<Tl���������8�pw��Xw�"[����C�c�?��g����4���!۷NlþfAv�l �V�g�&��W8o,f�|�$��@	�wv�u�4��ڷ�ٝ1�LT]CQˋ��5�q!s"�Q���2 �n-�&2X�h׻�O���v~�n�P!�r��
���5��wR���qA�^I*�����8
0`�_�gE�e��p�qA��	J��uL@@��yG��=�*ί���u��c7e�c�~���zw�������k�R4%%��ĵ��*:95�M�B�u�-��
&�8�A�:ٮ�M�jX�6J�j�]\�?�4._d��xc��Ļ���&��S��B*�R¯@�0����;��&;ԟ�cR\h�]}5���l-����m��1�GxLT����Nm�/چ19���D�&r�~�OQX|z�) GQOa��	YH�ڸ���o�Bp�ݭ�Mqj#� �05��b�񣙑�\<�CǑٜ�����b	W#�ggqW��Ť	�ɨ5�#���"w�O��c�?:2[B�`��jG����!�=�^�§����Hǥz�*x)�U`�|�Z��a�+%v×��>���C��Gί�H0�qx)�߅[s�����IwF]YwyX`��'��Ja��-����C�vQ�Ny\1��])~�7����A8��fPm�KO7���.���D�}U�ٴ/�a�R�j\yF����B��(ڇ��8�M����|u0�������� ���۷X)ޚ/�9����T�5QS�}0T7Qy<xes��b�Qm��ܸ���	W�(�pmk�y�L�	���(�p�)[bz�~_m"=-W#�	V|��F{F.b��"��������z���U2ܝ�-�
�nF�+�: 4�A˖J���m���h��#S^�oɶz�FC)"�Q`$�n�>";a��'Ȏ�9G�Ֆſ7cn��-��vc~�i�q�T�-�*^O�:UJ���z��=�/텏�zwC����="��Y8�2S�R$�6��q��Bֲ:��d�J`��x�~�ϩ,Q ��B!mB�S���o@��*w\^JA1P�*��	�n呮��
��C�X�]P�pgT:`�9�Mβ�NuBjA�Nw�T�~�FQ V�mT�qp_�C�(���Y<:0q��Y&����VuL*zHōIa�O`���TD�x'�y�C~"�84��䇦NH*���sٓ"Y�:�dO� V�3Xm�o	"4 ;��t��=�Zla��:��ya��S�y$�;��<C��I�E,��[�J�yK����[����λ�!�DS�;V�ѱ�#�jNgwg�a��LR�R�f"=�<�F����C4�	���n4�����܍WKb�*��rDV�W�Aq+��:˺��	K,i'ہ�n!h�=ќE�b`�Q��^��<����śؼS����D�O^ٮ�?B����z/�3��3�1��|�f��x��HQkX�"�C�Z�����	�5����4q�����i��Nv��h�N����:�'@V^�k�`�$��[�ӇruM�N�����U�F�H�r�y]P
���`O��ĳ��SZ�A��QZ��,~*����c�����3�}�(P[�2T2=d��L�yW����+�[%g�A�2+/��>k|��?��U������}����g���i-(bq5�oz�B+L�m �WO�+��=C���՛�c�q��Hy���?�׀�z\f%��
�y���ȗ�Z�	�@re�=&�+Hb�%��b������Ռ��rI��.�ćz�g�,��Ct~A�Z}��Cѹu+7J2Qε�F)'H�_��G�m�}�ﳸ
�#.��� �;S2�hA(w�ľx!Vyg�ǩ ~�I�����k��
�'�=W#ΒWv�׵��p&�í>��GQǦ"���`�؍M��w��_��<��/,�]_��ś������WH޺U��E?wA��5���*��}2��J90:�xH��&��#��!Ԡ}���8�)��J�Q��k�=�y~[���p�h���}NC��P��^�K
.8��%�i5و���He)��)S�B�b�RC����ml��g�����>�<�ȇ?A�9"s�������2��BC��$�@P� ww� 
��#��FE�<�*�b4�1|����EP[�ռ$o2�6PC�K �A(Zy
��8LH-���P��Xt��ڣx�sH�y��N�]�q�r�m^Lk�8�Zŗ�21�̎����f�p���񽌓��4l:��(�fĻlc�c�+o���x�����0�M嫭�?����M��ZG��%x����+��6m�ԍ��k��dfn`R�;�D�����B���C�L��.���������S؋�/��W��:��+�۶�����7k�&�����Qx~d
��vv�GD�=E�0��	o�Y����1T�/���N�@����0���ZE��6��O��CZ~��4S��S�I:ܦ�;E�_�wEu�v���֨}73��Z$�RP>�|�����vD�8r��m��gp�?}�Îf3[�i>ԛ)3F.�
�hb��k'�c�V����d���F�ό�7��&(-%�K�#��*�ks�����zo*��[����A�0u���O�O4���ֳ���G�<�s��٬O+�g7Vo�`��1��d�B�� O3�R���:A@R�F��M&�a#Y�"�WO���Mt��:����ӧu�)K��b��}:�u��C�R�� ��s���l����ق���[?�r�Ed�p�-.�N���P�֦����W��6 N8�SL	�(���W�y@���Pf�5�tu\�=v�b�TxG\��Z)�N���ϻ�҃"��_ʍQk���#SL�M�@шZ�cMd�/%��P���Q�٣o�C�j�.tΙ��5�K��Ƭ�o�,�o�q�J�'�]N��ec�+�~!�$�^�Gz�YY��\�R���}��y]q^�7k��:�z �!�=R>�nC��:�T_P�#��!1�Zo��<�̗���z23/�u�.�c<"T�Hy�Ρy����1��v��qC
��J���ikJg�x3����)����\ �q����)��nC�
���u{Y/�/
W��]R�+�{%���|�'W�7 Rg;�#�-��ޛ�|L-���n��E��.��Y���36���;�v��R��uJ'٭Тshq�z����Wqf!��x=`6ߩũAt/B����[��)���?�mh���"ɐ4#�U��m�L�M�Z�f��s�5�K*E�'Xh��d�	,sx��*d�F&��|aIek�ЧjO|��'����7f�Pc���"~�lp���:�{b��I�KS��w�=E�\��,�i��3���,���T��<�0.獼��B{�zʥ����A������xEڄ$�T��Ȅ��0�	o�|�.=����{1L��lWo�s���у]Տӳ�ޘ�/�s��v�I�@��!�!�N�4���Hq���1dE�$�50���qG���
H!:�[�6��E&�'K����綛�pj�ٰ�ŤU˥�`E߅!ծ�W��&b��A������⅟)<���m�!>��-������4�64B
0��`0?�xG$R#���Pq\g3!��.����e�5���"����we�O���'o��|lj���� (��DFpK��0� �(?��JF�Ɔ~�i����=6����]��Ԍ|z�sU��4Q��,=t����
�K<�8r�E��S��U|��-����x�m��9r3���PN��vRC#M4V@.��M���m���%%6�3I�iD��s�c��3Mf��ћ���0
�>m�{�<�7�R.����_�S��+��s� �t|{qӱ7o�8ɓ�SӠ���}qKX ��l�Ta��
ͭ]D�����|%mn��v
��n(Pti�'Q?� ���v�G�4��h���;@��(��uӆ8�v�j��M�U#ʮ����U��f��[[Y�f E���Q
�����u$_E�jǍ\��=��n�?��u�`M�������|7��(��
$��B @�C?jy���c� �&��.�{gN�N�P���_�?F I�	a�o	�)˞>F)%�T����I��S v�F�)s�x6e�
L�|���6��-����Ǐ�_�I7�
�ڎ�'P�]b�zmLQ�0�V��vu��Ka�\�mL�3��]\�n�+�-��pq��h0�������:a���,��А�c�8��P@K-��m8W���|:��Ck�FO����2,f''<@���|iŨ��p��8��l5��݌�� ����7�)�rDg� B���3.0Rw��p�]�=ۊ2�]���lwy D=ߢ�7:j/M��D8'�wI��'%_|�-{~Y�`�?�����������6��3:�k�1�d�$j�l0��>�&��_��e�~��?ۗԮ�H�ӱ�3�=;L
�D�9�_�N���I�-Y��*�C)(I��˥hOi�d���9��T|
a��_d�"L�R��c��:@ ���xm�<�eԷn���^B��5݅EcJ]j*����S�ѡ�0C�4�H={��P�Rw ����aa��~�L��X�(��K���G���<��F�%G	Am����s�A8�\�3YF��^YQ��B�g���bQ�!m	C�֒C��B[��l���@��IA�@�����)PX?胑o�m������|i쥿r�y.g/���F�y��)E�oA�E�	����������ge@ݝ��f��1����G����D�яG�Y�d�N�j�s�˔�z�/@�z�����`-�i��@_q�L)O���P�5�9������tA ~�C� :� n�l�Ę���2[Z<%T�=�{	�j�3��{�����|0<����v��LqV��x���i�1�b�x.2�",Ms�>���d�Cձ'mZL�X\T��ЈZ���Gf���:��5��q���ۄ�.RL�f�Hh�#��a��F���ef5��٫Aѷ�c(Ǳ��n7������Q�,J!����tnD9��d%Cag���x�l3(ْ��R�-�?w��7��#��\�cNG��ŏD�Y�+���r�'�(�����\�I�Af}U:[�"����vU(\��;֯�t���Wx'<g�Z��<�_:�=,��s=�$��&��&k����:��tͪ��y��b�k��Eړ�40���ڋh`ۢ˼B��#�_�	�B��r��?�����)�V5=8����]�޸��h��Т;�C��_��|+�t���4������ac�6�``�~Ҩ��b�wM#�]_�FL�Co}�����5�X[�H�w��ȣH�:������_�,�H�����d�cg�������$�Єnfϡ�8V���M��=FP^E˦����]$ �x&*��i�_���f���q�\�.8<c��6�<��%�M��Mz�&�n������w�K'����'��l�����m��ۉ�E:ύv;����up��_P�b��|'I �G�7�ү@�U��g7����IF\�;�c�ֳ��.��K#w^%`k�#q��$�6>S.M�6����k���K0�\���2	[�7a�׆#a�G�#R*ΤH��a"(�PIC҈�TYclu}�Ң�?y6�ND�I��@�GE� ���98��j�ݷ���d����*�����$���4�zA�~����w�Q�Y(��Ô'_�(������C���n�B�?����)ś
�uIy�;{���KQ�S����>�	�$ְ�[pb��Ne�].]�?�ʥSPfo�e����wݍθ��wj��f~gWzYD/���w���0��]^�CO*�C���R�ӱ?���3L�5��rr����a��e=��wϪė�����#��}��Kں���ך��M_lü�]�a�GH�Eh�S��d�\Ebx�o..T�u�BpnK�hS��Gy �y���!�.�q�w�>.����_ڣ7�m@"�&�i-���5�`}H}�rGCԬ�	��N~�Wn�����d;�w�6kp�ȕ��K�^2}V���Mb�b"_�/�u��un����'��-�����Cf�s��#�9'Ź<U��'�l��gY
%X�:\�����8'��6`Ӝ*��cg�J�����9��.�٪ �[�+���>ĳ�T��8�#I��~�C�J�03��U�P���R�bh���z��G:��>��C�j�|4�T1��3�'�!��l)���Q
^��(�N�<���t�r扸Cg[~j�<a��ۣ7�ǵ�'Ԏ��5����N�]�nw�͢�8����V����ơ�����+?���d�@�r�tN ˫��<}�̱����M������?�0�!�x�̸�;	�"^,f��X�щ�2
7x5�3Ʃ�B;N^v�,����1
<A���qň����·��)ch��"�/�楞��Y�"H�r�DX�"�s?�����-�_9���Һ�S��:���E���vv�:26���F�' k�������e�cpkH�b�����|cv}�Ys���^�
����ҋ�#�����0� �M�k���ۡw��q���!�,Z�R��ӳ\�����sd.��W`�DR�/�G�0�����X�m6>���p��ʊ��V+d=�h��VӖ�j������=��F`�ur�d ��0��S�0!>�L	�%�V��^��D��P��:!sQH,IP%m�<{,D�R���u�"�E��+�E�m�<�_9���%��Ӌy}ׯ$BR!<!I2IIx�\:���%}�;0��Z}Ma⒭R����\��Ϩ�U֭��������	v�E��a�i�����b�E��b����������*E�S��}H�#裂�=�ɖ��\�(�x����6M�x�	���|���Z#�itC؂� �eZڟP>p���(\9#H<�QP�|u�Z�A��@�fWP���<��1�R:�<��Ӻ�:%ka�,�׷�Oc��	���&�+�Fp^+��U�OҪ���3V@�X��!���H[�E̮��6����8,��sNoG�j��;�q�e<L�[av"��l7���B	 �W L"�\�K'bJQ=0�kl>j[�.ɯV�SƧ���,h�Ŗ�/z� �j���4L�G���l��/�|��:�_�F���|�o>~��r��cֆi��������"F;1�r��X���X����'й����������E��+���A��܆�$_���G�+������+\ŵ�T0�'��@^���&��@B�[��پ���U�C��&
��z�'f1��y {�S/ٽoEz�[�UP����;7N�bHI�6�,N'�,gM��ۥ� ��sM1O����׌)��<�J"��}�X�7OW��S1PQ6����Q���5J3�g��k�9�����]A��ۄ]&�Q���V���^]*��]�׀/�Y���H�Z�1W�Q��H)?]�)�xIN��d���*r´ʔ*R���H�<e6D��J9�ſ=�9�:��#V�#�f��Gc����V*��ޚmZhQ^y���^�e�D�������E `�m�焟��ϳ�u�;%��tl�\��_B@���I�P�>)�&�\�%5�F.T��Y�-��8
׻�Y. y"�J a�"mr�_�8	�ځ*�e�ȺoZ�t�����PO�/��y^��<g��4g������u��o�;��쟫X��|U��XA�A�Z
�$�ˮ�ҿ��OJu�N�� �fتo_�'��(�ġ7�����2ԓ6�"���,���j�B�8��gn\�/V�3V��<#���{U�o&rV���W���Ƞ�GNFC����	Ƶ�����>i����;���VԤ�Z��n����!���l���Iriq��lFjJ���nzr���ɳA):֐CO�1�����]ZY��)/��d/F�S�ZJ�*��{��i�v�U���������pZ�������3�#��Ly%����:�ς��:�ř~�3��a]��%o�@t��-M����-[�"Ԩ�9�A_�IҒ_����8�� (�׽��7{>E��԰���ߢ%?L���v/���X�q�#�=/��N�o���L=��[�m�dɢV��n�h{�φ 	d}oEnx}Ћ���ӏTWv�+��8�᜖�d䢋�[g��.{z�3�{��Y�u��Ɨ��ϥ"�|�琗���)L�\څ~���rV�k��G�$�ޏY�8c���}��2��2 ��}��mPḒ�G%a��w`N��+����� ����c�V�s�_O����tA�j��,ͽ#���7(맺G�~k��<:p~�an��%�뽘E�ZN֣�k8��d�m�>D͚�oF�h�P�a����\�5�?���֞'�$r�~9?ѓ�A�֟�p�B�krEA���nb$���SQcˉfS�>�����{��H�1nۿ��l�
���� IL8�b����aj���>+ �����0rs��%�eғE9Jq�C^9��^��I(	_+?WU�|��#g��T�@�� ƶ��Ǡr���v5#/�J妥eC{�J��zI�4O���k=b;�>��5��O�q�/�b�b��ߖ�sD^F�3��H,�c�çޜ Y2*٪��w����o]CZ@�9E۱0�'��n���m�_��	}Ժz�h�3���+X�ZHpT��%�I^��߭,�y�²�R�U�̖-�'	�8>�Ig/�Y}"�	���Z��aH�հF����!?47xmh-��P�����[:�߽��E�'���x�Ղh9�e~K��R2#-ަHY�PK$��zx�"g��|��@���<�ֶ�"�r�K��2�t%�JXƢz�0)��D#\�i<�1���0��}F���B��1!�+ Uz~�ɗ�F���x���/���U�����n��ͨ��`W#]-��2����a�����QT�X�����ˍAN9�s�ds�i�/�:-�g~���^�a��>�}~�U�s�}��}�g<�3F��?�~͘�d�s�!W��Ѥ�����Vkע�+���ĲuDb�v��c�b���<<��]jח���!B�4�b4[x�_�����O�:Yh�(2~L7~��n�,��3�MO�{��r�Z9�sn?E����y��۩s���gE�ӉiJ��K0E����ۋ��no�S=��O!��m��{;�k��`�}�;��_��K�[%���06�w�Ϗ@��<��qӝ��� Kpt�����2	{���"���y\:6wu~��������miӍ�=[�8	�dۚ�b�<�<:즲�ǡ3A�s�C�|v�vэ��`\��i�}�
�lZ3�8<9|{[)g�q�o�ĥ�� ��b�?�/���K���t��[�؂�u�/�.�[�ո!�%��c�{��_F��F
�n�\�F�|ӂ�8�`#=1 �����
`�M��m�9=����]��0��Y��
���/9j,�w�DO��cL����K����F�f�t�L<��>X�h�6 ��>ѹl53����0{��x\�:��/�2�+*:s�%y�K�\l�w�H>�+�F�I/�͖=�Ê:�"��=���+߅j�t�M1�"x/��g�>��6=8�S>�3��;�1A�O�Ae�S�u�[�j/AY���@ѧ����(g��Ec�%��:�Ѥx:V�o��� 77��&��.��h��� ٙ�5��$\�"u��H�?���F+0R�Wk���-h�:J/��G!@��9�.�GM��d����L;���Y�������+(<��cws���0���8��@Au-C����/p�B�/r7YCL���I�.T�����ҮQG�ɉ�5:�@�dL*�Ɉ�!�M����z�b���!�N�_@�Dwz��c@H�6Нd�<�<�{lt���O��y� s���� ��%��qq�X��\%jV"�`Tf�WD]��1&/�w.�S�Ef����T~�8a�>���=0���
���;��/�\]�����t6{�[�]V#�"��$��F�1�B�J*�>♤��Ѡ
�H�sY�H�"��r; {r��GQD$�:--���P��?_��u��Z������p��43� ,M���r�d1��8C1D�-f�O�����<��8�S\|v����%Udo���8�XJt&ړ�#�¬dmtՎD��o��3���8!��|޻ȥ�c#�\�d;.�ݱ���UC��n&�ͦ�义�3��D��c�p��VZi{V�3���|�s������6��>�kGd��6�n�0�$^vlj��e/lj568j�ԓ�,���lM��У�ǒ���|��/����?E�z+,"�qTo�B�ƻIqD{=x�)�Zo-�n�}�ε����������p��SBD�8��y ��=�GÒ����%l�b�rE����4D���+9U�<�P�t�����������=_h�a���ϹQ�:a���(?�h��U	� �G�+���| �T�%m��N͕�R�FyY1eO�C%��}c�� �e�(��c�J3�e9�P�kwX���qh�-RvO�ϩ!��뫶ڗ�@n<>9AOּDD�E�3��-�Sa��(ϕ�q�)(P��q�Av����^pٖN�|9&>>���;�:�����0(�a_L9z��ʣztF����.5)��9?/q]�m^i������^�5��ZAK0N������R���ذ�qq��\_��G�G����*�c�{A�� �xB��u�[�-o"0T���� ��!3�ިԎ�G�T��)�56��h��o�2f���f����p�~��zJ���^���[�Fl��� ���ʉa��a���w䜰�ص�����!��>N��c��J�j8.��OS�x2ε�u\NJH�?p?ST'�\��|�Sb�_��)�~=��~�����m�����-	K������VU�1�)���a����@�U�US�)��D�)���i�sɛ��hC�Op�JR����u�0>��yR|�=��6pg�ל%J�T�;�"D�[�F�d�4$?v@�O[y T,�f$!R߾���e���&��$)�5�/�K���0��?�����_-����82���ح;>�sm��g�SТ��o��G�[$�& �w����J�.�O���GI,h��8ž
?��Z�� g����Xh�G��
�z�O�[A��ڼt+]�uyd�QxL���k��I5yt�|���F�[��4�D�gC�؜o�xX�+7^��^���$r����l��c���߻�3M��HI"nP��Ǒ����+��������b�H@5/�RUU�2l�mh�.���1�FK�$��?�¶�L �Ѡ�M�u����A%�e�-7Ä�ֿS˗�ϕ,qf5l�ʗ,0Um@ K��B�����q`��9�����Wc�ֵ��yc��\yeL��j����.C�^�	aD��*C9}[s^�������Q�f4����{x|���u0R4=�ť��DW���va8��U��U���zrG��� ��h�\�mj^�ɩ����f�w�>)d<��n:L$��	?�&>��n�ZŮus�j!;��g��M������zp'�g���R^�d���&]�_����.��+�#K'<3� ��wnm��'R���������\

���x̺ �R��jg�_�#��+���=�Q�W��Pل�T#;���Z�b�@�]��F�M�I5�Iq����?)L��͔�Q ���x]�W�V^+�	���I�D ����`�s'ޔ�h�F��g�Pé=;�=g��hc�_�_�(AkYo�5ϒd�����%���m  ��g%��o�ߦP�,Ly����^J"7ҜEG�9��s��\?�p�?%��V����[�ɓ�(F�h�<� [u�q�J����y�&J�ǎ|ߢ�j%�a�3�1����K	T] D�^��C� 8�>6�j�b և�V���CR���-4�	����'SO��L֥�쵄��0R�R~���¯���0�ny9��
���5�x�B���&W����܄�67�0�H��L�6�k�%KSИa�-����-�B<���P@I=g`����â(Ʉ���KE��>4���L(�o�ς�:72�sr�l4��F[�9��×4'�3-� ��	�lw^����b��?�(-�n�بdK\>����j%�t�2lh�\2������ߧ�M|��dh��:�v��dqi{���4��c�OӁsJ9?{������7F��kC��i'��eͷ(e����w��n��oM�c7G^�㯟�y�y�=�[S��y]�_�����������t���jR7�̉�� �ٳ�q�G1lw���_�#�#�|w��ͼl3/�l�,+� � �{��G0�$`��O����<�vlh%�����ſK���Y��D�a�b�1����ﭺ nA6oU������>a��䁧�G	�N��dU�Nl?�G|���H�,�͹K�ƚc�5�YC�Q��PU�{���|1x�w��P�Z�m�}f�P��_N��b1�Os/�i^P2R�8Y TI0(}����Q�.Z| xv;��KA�i7��`���$�U|��OI:�C��މ���Y���K�o���K,7�#20AFz�qiv��JLQhC6�n2�uԣ��l� _��r3_^z���z��/m�'�(y��.���U�L�_��)�TЁ:���g�ۤ.�$|�jAްȹf�/�d�R���������7��W��m�|�M���2�:0�G�' �|�>�Gf|g�4�u�E�K%%!�6L�'Ch�{P��0k�yPQ�r ���ї ����Pfy�[�S���=�)�+������6��'���o"�hS�^�/�ߦ��nD���~#��j< >�f�=�hv�����:t�vd.!�>:�$/ٽ�{l6S�E�yQ��{Ń��J���|U��y\���I�/����o�W#�A�k�F�����Y}��n�J��	ܬ���du�3�;�~�z߂�W���.^*!��r{�����aj/K�����&a+;� ��З��JmD�{����g��߹��N�������z�`�� ����z�@{t!�������H�Ȟ��Ӥ߀��9�9;�pK�_�4��:c���M�w Wh��@���$Kp)|�<�?�{U�� ��ϭ^I�ꙻ�\����s��:4J6�*���Z��R�4q�u���O����lA+�gG�c� �����1���|�b�Bu��O}(��"�L׍Qm��7xR|�8����b���=���T���o�g@!����z	Z=����HiX�r%�/��X`�`����$�������{�\�u�/�-H	~?�"��H��c���ﹽ
|E����Gm�t��8���ށH����yT��X���\��_i(�%R�S\���p�Vß����Q}Q�H������ʿZ��V�]\�F�g�nAx��#��o���r��\�[��{�q~̷M5S9[�;�+y���8*+Ń�����i3\���
��k�+�Ò�$���g�d�ä�j�1��J 嵽�Gk�T��\��Τ<h�4��5�{��V�yL�0G��|�3�2蕯5��/��8
;V�҈P���] �ՓC���
��J�0�IR��dĶj�ˡ�6	u������3��P�\�۟����Owj�Q	���C	ܵ��v[u���҂~�h���@|.��p	Aٞ�l$R������5¥��7W<)�|`�^p�:�d4��`�+𷇼�%��oB%��M9����3<�h�	�� m��ͺ6&^	L��n*R�&��!ܫ�?����xx��x��C�!we5����k���%tQ$>�G�N:$*�J�;>��[y7� ��&�-	v�J���b�@��6i������S��1�Dr�_�x�`J��o�G�A)�йp^<�@��)�;�v�'!���<=��o�](���g@;����
E
�$�Z��ZwOѼKɛ�;+$&-Ag���Jm~=뵧ѿ!U.}�B�������Q�  wR=��c���w��?���*��Ra�̵�;�ʨ/���j��Jn4áj��^Ub��aϞyӡWޏx1�>X��F�b����tn��C�X��w�+%GsE����n�~�m�gH�;�X.W1�_�hD��/-F�<�fl�2��0q-<f�V��3��e�}��K[��U���
��B�N���V���̱{g~	*̹�T�j�@�.�y�;�'�j�޻����Ѕ���)}���se킒7@�PW��:�'�U�o���x�s�v�ˊz�.'H>��Mv�*��G�g���{{�z�?]���S���j�J˷�����ڣu2�t���V�h���{�<��k��|�\+E��Tk���X�i��j��(~�!W�iW��K׻�=����zO_�:����m��o*��ܖ�0�_��_^'��9�D㙭��S�բ'/�>h�湬�cLj$���\+�"Uʥo����цI�Ԉ�"�L
�3�˴e+��Г�PöK�a,8�o��vpC�xKE��@�0��n*z��x�_?3��:=��Q�7��n+c.vy��jY���z�&���@�B�}�]���38_pI��&�b��7bx .�G�"�8s�� �$�J��A�2O7*�7��L�T���ˡ�l޼����p3�Y��y�`"��p;AL,/}���\����;�����ci��`��nbO	�����u���z ��N_a�����\:��M\���7wO��g��ö?�v�ҟ��F���i��H�>�)���Tm4�Q#HJ�R��;�י���|^��g��$R��l�� ���M����d�� Id�AV���=�>p=�`�G eQ+�p�3�37��H����~wB�@Q[\?|�
?���"~E J��wts�ia�0A�d��8����uz�'(>=���撻p|V� ����	a��u���F8>�����K("Ih_�&�E���͚U�$���%myy���,�BP�;J "�G奘$��ѳ��Q���w��[Dq��&����{�iGLYg��.�$����P�Y�wB=?�^#�G�K�F�ߛKP������Y�=?��~��3`���'7�BoG��b?ˁ�E~�ߏ�A��i���mt��FV3Eբ��)�}[�����=��|���_5�+��j����}�����4�^���	���3����c��{4��4��$���s�����=�:�᭳�ѐg�M��C�ޠ�x� ��b��T���lɳ	��C��:���P�=�v��(*�Ճ�8��3�t�7~�p5[Qg#�<� ����81/�5^��'���BoMm~��L�:�(�nƠd"Y4�Mb7j�"�|nυZR�No���W�NO�	Q�������pa�T�d�9c�OR��$v�%���T����9*�]YOC?~@i��Q'��:=FD%����_xgj�\ZjK�]8~«\��ד���ڳ\�]���+��Z[W���6�}X���3�^	=m٩������.|�l��ʪ��$�����'��C��a��}IN!\ރ����Vyy����+�*�Eut�?���R{��/����1it��-eL ��pץC��Z�ʩ�g�S@2��p� ��9u��Y'�G�]�n���hG����~��f�ݦ���V�8�U��a*^�zyUay����Ӿ���fO��%��:=$���t%��J#�y�o��(�>�lH5�C��Y"��@��_�C[���J�� �)���h/��3���ŷ�n9F!h���+Ŷo�v �)�ȫ&Z�������=�u�u
��ĿR[^�:>.@no�F�`��
_��'A�*��<��T�"��
����
����P�U/]3c�m��'�����o�'��"�� �9���r��a��xx�n�n���c}���Ml-wx��ъ�Z�������b����4���A���������pѾ��~�s��uM-_�H-���������vk<H�]�Q	��"��ſj&(�I�,����̏}4����Gr�!G���oL��H]�Ǐ�Y(�CI��c+	��[���%�	x7�;�%��x7�{=�ŕ����{�ŗ�o����)p?&z�/	{<=}3K���v�Y�6��G��=����H>H��ܞ�l��l�9�"�M��AE�Ї]?���*�-�Mp��<�WY�;_7�r����~U2*�aє��儅��}�N���0E	�����"��/���եXȟEHYf���d� ����%�o�6�]^�g&,d�����e�J���44��
�u�֋
��-��yU�4��+�/���������{����6֔�]Ϗo���y"ڧzfY)T�[�B��Q�	Mr�C�=�X�t�xw_D�݆�*oS��5�Jd]L�w���}���<_��{��d=N�`[ˍN)k�y���=0��Wo���Q!eF�,�p���գ���F� v�8gP���y^��ZY�"w����=�Bǅ�fK�3��}�ϗ�
����@��s�C�ml�?+��C���y�����.Yh{�^Z�b����1Ե܅i 6a>ye��j�y���^Z�=�H3k�����&��ku9��8��h�tg\�0[(L1R'ڌ�����p�8���aZ�q���n��t�?�Q��� 	\F��E��[��Ó\���,��j�62G��,���=1-��� �r$A�3�A5���x��=�Jx�Mz����Q���]���C�\v8*:�r᳻j-�c�<�[���IK�jџ 1�����P��F��L��f��w0�l�E�O���vD�3)45v�Y]��{�´xy�3-�dK�L5>�i`Z����@�Yo9���ӥi��C��x��N�cM���8�0���8q�~�{l���n?.O�
����ݍܦ3z��,����<Q&}'�'��u�����UM����~@��ՔK[��$�'	l��a�Y��c�	��7�M�1�(�G.E����,���J��9 I �!L��.��%$h�Ņ��\������M��Ugߝ�����?h���,�S�޺�4���ާ��Х���L�J�0�ܔ�
6r��.�.Y��0�ڳ�<?�=��3�s}�~ �4��h����NG {�;��� Ml�5����K���O��t�9��=:��h�$�_�1@�:��Qvz"�u`�k�4���+dg}�� q�
{��~D�:M�<4W�{���}�%��4�g�Gc��t��A�|��`?=F��x���-ri�������t��������჻�>\C�~��L/�1=����瀍�{���v>��p,�p��u�� �����T���l����/P2GŶ���MV9۪{%���# ١�3�u�W
���]Ӧ�G�&p�`:�u�l���� �/�Ѵ�"�`Eg�@��m�Ӵ��ezw��K�|X8�ŧ���{$����b��k"�G�tB3��=8�7��6�F�	FKs
���
���⢔+g[+>=���\Ȼ����u�[���5�+\B����S� ����he�[��O��y� ��x|�Ŀ��G��_��'���qy`=U��?� �~4�uʼ��ss�ri_�ܭ��$�ݣ�?��`Pw���
�C[d��ԍ��s�!-�F�h|pM8�_^_rn^�h�Z� ~���L���:N}�>�!�E��}�δ�P" �nb}��*�ʧ1�d1�'���x�n�a�d3��+JJpWR����캘/�-N����bbl��qz��":�@�mz�I`"�/D�1��	��a�܄[f�J.�}n;<�6��R^�wM7��驌2>M�����E�Pո��}M��q��l<k��ce��&�c���M�?,��� 9���$��m�/8���b�5kᡦH6/��N.�QhL%'�8*���I�l��'�WOS�ޕ�$�����Ŭ�b��q��[}�9Vo\L×���nlb��Q��z޿�Y��λ(���*�6���%z8��5�]�#LD:֌�����38��{��fpiǿُfPz�"@�3��F{�[t��h��v�_��e�e3α��D�|��}�M���:x����}�!�cp}����g����l=}��\�O�_��~�VG�c�	��c�~:<K7b��dg���Hv���]I�'n�i�C�W^�OyM���q�Ği������Pb ���Z+�>9Q|�p�ƦcHƚ�p8����������$R[�Aj���q&���������=%繰�x�]��Q��r��Ln��3�[���k����!gy�$�5��dr�Ɖ�����Է�M�{���L9׭0��&�����l�on�R�WL܋Sg�i������0�E��w�mS�R]Η��I��9��[#j�T��9}�nR /�f����O>w1#5�f��<Rz��e(���� �i0/S6�Xr	m��s��~�O��e(�P��S��>q» �e�z��j�m&� ��ʹ�B����F�a�H��x����,g�h�L����fn���3�u�Z��u3����I`�ڳ|���˫5t���؏ _��Щ�H��?._�-C[����*(��6~:M]:�{��Ll/����U{?
�D�S&[O(B�h%*;>A)o~��d���n�m;��몦?�i�x�������~���O{J��{΃>��]��|[v�T�<���Z�b����*����_J:l���*��>� L�8=�M�����x��og~�t�X�["S�XHH�8du�(��}a��E~
s�~� ҁ�X���J�ǃ́�')�F����t�텻i�풅�P��7�-<�w��������Z	#�Zdg#�+����]��-��u��q���]T�n�;��ǉ�nGL1M\q_^U����eTo]奇8VK���Vo�ϻ;{/W9��U����d|���$��W�����߆b�'�~�s:��s|���x�Ì���߅�<���vG��V��釿n��K�!Y�+>L��\��)��E<��Q�[��U�O ��U4̡P)��姯���t��|B��5M���뇯VO�"�=�=�<��.��C&ڿ�2^��Y1����t �����8�����	�@k?�y�p��[�)�X;���$4�ѹ1�������ck��b��������������z�~=>�_���Aq��rVq�'�?.��;}��[b��+�k��Fqm�Ԏ�]�k���������T��ڽ�����F=q,�����*�|�1����4�٩��g������E�Ɖ���~�j,�n����'��Zq���� ���g�x��Q�/績,�o�������q]a���ӵ꿼������tw�v�~���;];��� ���[�1��O\�<��Xwc]6��}~Y��'�cu��bsh������WqR��X�LՍS/���11-W�/�̊�&�u���`�ύ����r�̽C	��-�a�'y����HU�{R�$6�4�{,2����FL萉���<]����_İ5�/�K	�.��F���[A�x��g�5M���{�~�)�6���׆�3��S�vpb��R�w
��&f��5A3���ދ1��%�/�x��̿L��쫱�����QO��h�7����,�aok��<��8L�A`-@3_2n�S��=W^�<��l���fr���{(U{$ݥn	ݬh����'�)�| ɡ9����}vߞ��6�u{��H�>�;^_���դ�����_�
�a2�A3��m�]�F�gj	E3s���dÓ�'R�.�N�߹�ֻQ�F�5�-��S(#yyE�<�r�;�Ly�+� ^��!^.�99�q�v��hc��eG�Fʅ�ь���K�	z#�&k��5?�"_݊�fs�§�֙���G�:ȓ��_'}X��!3?p�5�w�S�5���e���F�����`�[�b4y2[��Lp ��5jr%g̔qwB����mh��š��6��S�/qN���$�x�;P�Y�����A�PTo܌����5�F�A�X`�<T(�[ݪkމ���;�Z�Q�Yk���>W�$�z�Gw c:��	r� �|����ɜ��<=�ڠ�{G��o�[$��zt-Iv����r��w�J�Rw��o�"��S���A�}<̠��(!��9�F��??밣�_��$g�_�T�L�9�ЩuA[�{��)�V0l���t�*�,��|�t��k�Y"<z2o�oO�0����y���''����_���O�s��l�t�on�S\0L�7*�mL)�h�S�� ���뵔�yL�!�� n�\D�icߝl����޴6�V�M�a����VA��	��F� ; S�Gޤ��Y�l��J_b��R���嗎��޻�7UeçP�4UQq������6)	����%M�6�&!9��(Ղ��㫎���̨���e�BAn:���2�Τ��K9�Z{�srr��|�����|��u����}[{���gȼ퍔�5]&:=�>ض/���.�m5<;��Ҵ�ˠ6 AGs���o�!��A+���*;�`�6�4�|��1*�*���Ek����N4�m�fop���tN�_�߾ۣ�pvrD�w��D�����-���X{T~���.yvؔ���HQv�S�����a8��vˎ�YV����å���}�+�h;��2�˨H&�W,;�i��7,�nˢn?��|0�F1g����a)����c���}��au{�U �-�3av�⸨=�:�(�,"�"i������;�����3��"K�)�{Y\:�3�aL� Y��P�f'���Fo����9��^����M���S��.��h��)����P�X�'��?�E�D> aR����̊�.2��0��U~��m�.7�?�Fmۙa:�CSA��O�"Uie ���#�ٶ�[���9�d������vTF��)�v���_Z�=�M>��	�hW�<�OOCy?�dx�x���fd���0��o� �1�_�N6��W�����ḋ�~��OQ ttce~�9���ۆ-s�(�a�/����d �l�m��D�i�޲����-�����L�zӀ4�f��W�l���ٳקδD
wX�/q[
��]Z�D��5��[S�YޔJ�\f��s���I|�r�	e�)|��Ͼ��{:���:��0��e�u�M)���N#�.��g}�c�ˆ-l��[Rv?�0�Le4����L��U?8u27� ��y��o�����m8[q�b�<����[[�]Y�
m�k��ρ���8�~����h���`��^:�4q?[a����ZvlC�<�c�5g�m�,�@�-���V`&[N��xC~yvd�x�ֶ=i�?�}�Ț��s��m���7d�X��gOV��{����Sq��"V�(#O�#�����Ͱ�;L��a�_����.P���"������Í�=��X���� [W����Y��h���(pֶk��s1��=�� ))���X�'xf٢���a�x�����}��NR��,�b'�"��[�<�g#9~�m�<���L�ՊP�c���mf'�
� e���7
�ɖ�݆��[ɛ����u<��L��f�=�Zd�J�(�:Lt�4$��K�	��k�̪�D*����E�zf��&��ֲ�͆-�\cx�6v ̐m�{��;/5GR4����}�AcJ�(�G�!�1�.�d�x��`X��f�u%\��(p�]�5̴�����H]�TJכ�D��=�4���mWR�gm�J	�	MǳTk�f!�%����ɘ+����g)�>_��ىF&�5��1`e��d䑫�ā	��۪�w�s�Y��8�1��%��Y�)i�+O��aa�9�*���[��l����x�U0=|���)=����x��S)�1^T>�����u�\��'V�r�d6�B� _S�R��fj��[{d�� h�J�2���6�i�����Yo�T�v��=�mw��#C�|��,�=~�{�a����G�jX�*h�nIB���w/�O���+�v�r�0�0��Ȱ���y�,�pTlؾ/�0&ʩ5���&�d���W>�
�isS�k<&�	���8��y��z���	�AA�k'�oǠ]�X�<���c�qKy�zc��le�zwb���y�-��퐋Ar�5�j[#v�K	X۶��f�ƁR&
�l���m�d|��SI���En�;'�v�@�<k��v����`�1�5"�:��i۝4 �B��m��vy-X"�= sMz�����]�Td~��-��J'1m�Z�B��F}L�OX�MIĞ�~���Έ�N�����fMd_˪��\�v�0�ŋ� �q4�mj
�q�����>�D���d{E�l[_�;��C�9��#��aW��B��~z��g{dy�ZK����J����h�[����߮G9%(^v<��"l�,��si�121��7��/��eЊi�9����&��њ/{��A`נ�ݶ� 4����� ���XT�|Ra��G�vp��.@/��������<�?�j�Q���c��"k[�h,��Aض��<�7vp�c��\A���w�ළ�kT	6Rm���Zr��b�b���ݱm�@��!mdV�n'��$��Rx0��0:ԻO/<�����8ǚ�[�r,�d���8�����l,�5հa>�����h*B���!��F+~�+|0_��_*vBV�B0)�EIt�署�`e��ύ��(��`	?�Ĉ��\��w��@'&Q8����RϚ����RА����e�*��'��Q����<�3t�lБ����Ȗ���.#�����d���7t��v�W��)��-�q�f��`� ���uy���-���K=.w�\��.�ó%�:S�o-;=Ӽ>u�6?+��Y���)&�n����J�?�������e�E����m��������j�=㿢�ʾ�_,�&���)�5��P-��{�5�]dBه���sa�C��!��d>��W���B0�Ҹ� ����1m�d�g���i���8eQ
��5~��MY4~%C�nkx�t�1��R����(fV��ݞgFX�ƾ�j�чV�� e4�zh�*#e�����#�]s������lÆhG�ֆ���겎ש ���/�U��T�T���X�o8�T��g㸽�� ��Xû"�-������C�wH�+�[r�� ���ќ�)��X�������-1�]���B�F~7*�2����.�d�@q�Sv�����k;г����:��:F�%J?�l�چ�H�߰}/뛿v�+j	�6En��^x�Z�aJ�л�n�ÊZU�0VQ��'������X��S�xM]���xz}2"�F�AT>���Om��}��l(��DT���3\�y���Gal����������J}ph0�+�e���M=�ǲpT9԰��h�^��u�u���)���=�4�p>����ӟg����cJ�G��� u�XX�֜��P@xb�b�}��"�]8��F��þ(���Z��3��֛+�֖A:���	�-���Ϸ���Ca�S�X͢3�����:��(s#[n�,m�7�+Gܚ1��W�K'�)Gc�)slJêa[�n2���*<x�J3�uV��1��u ^5}�p)�T�_X��c7N�M�HH��8I����_�$(�:v�7�W��'c��Y���5He0e�;7:��0�@-+�+���QK�ͱ����NaY�ɰ柶�S��P:�v2`h���T��w:���[_���I *�k�KG��s�S�|4iZ��m�#�oE?o�C4N2W�'�]��Ԋ��:���hA�1��P`"[V��jl�OF��y��o3��}��Gd�]����l��@�n���ɏ��V���K��Pظ:'�%�p֓x���f���4]J�i!�-�=chn�D/���S�[k=tn��ȶ��L܍,� �C�P�a��Bc��Ciƽ������؊�&����͎�$�%R��}�u���y&\���Hjj�MX�ȅ��4<x���Qpc��{!��5F)�ba������1�G��J�ChOI��;��yD�� ��4�Ѳ�#�"���(���>�T���s%�5r/�޲L�Y"w�`w�US�a��Z�����z�� �ϛjX}��p������p���MG�o��Ѱ$�yƳ��ϰ,|_�d���������	�W{:���5����"�u���Ͼ�},p�)X�\!t)�O��η����!��[E`<G
gӍ�M-�/ˡs�dS�b��8�[Wd��c�3$q��8��5~{Wf}�`�%\	l� #�*Õy�Ҷ��J���F���e�>P�I�!���lxg�H7� �.���4�B��˝��a��!~Pis(�_��3y�R֊���΍g�=�#Rb����vX���5|tE?X�:}8�t|!�sr��/#�[�ȁPX�l�Ľ�-�.u�y�]����>�z�6V��ۖ�e�G�P LoZ"ې�����2�`)�<�M�ox諎_�bL���p���{��.�;3�i��mX�CIž���v$����%{6�U@�\f�#gXU����S�A������$3G�����5��`���ƽ�K� rE�� c�a;|=_�c?+SY���}�ݠ�Ȭ̇��db��Z�K_�����@+��<�rmI�qͪL�$r�w��!a����(U��,�n����I�	�o>�aGt[P��rb
����(;����̰��*֑h�cGٗ�[9����~�}n�9B�J��"KĒ����f�!(��6fG���߽2�=�;�:�N���S�m��/��h��8W,���C+3���w���|J5�����<��_([;��ٰ�iȫ�+�z���Kd�ȗ@͆-_E�ƯXE�gs�5�'��a��fZ��O���5t�h���a�	G���}r�����)��f�V�W��}�����{8A*d�������=�����O���~�0���V<`����� o_ y�瘆�mC��E��G������WW�ȭW/ŹϖY�́���"����f��7�Og߅87��Ϗym��3��A����#r�%�>��b��A�4�Sײԑ9�̰g7�����?
�6�#-t��;�楅Kmx=<\:��Ll��;p��o*q.J�}�N����?-��G���>)).��/��bna�PDU��bq�5|�p�f�w��0�%x����f��zɿ�_���!�ߵ�N*��0����(ֶ��_m��u�[c�����	�PIF���T���+�ˠ�}-��}9P4�Rc�X)~�g\*�|:��"<��YS��v[/�f1������a��St-�*�d/����@H7�ǯ�n�y�l�#���F�=�"%5�4Nf0�V��?"��Kj��6�ah�Ȭ��WAj|���#ѧ�n+U<J���i�3~�Z?�D�2
:�5*й�T("+�YA�����Xvw|�'k��\�&�+���l�_�P\È�>��(O�!�#~��k�L�/��\��ܷ�f�P�πq�[0l�a�=����ӟu���Ꙙ!���q�WԈoPEگQ�(׸c��E����K���U�r�>�"���6�ze���bZ�F!�E�e��ti	���B����H�S���Hs�&vNk�������S����<�N��$2t@�㫲E_�!�v&��x�xZyd"�|'Et�T��a�-���S�<�8��/�"�hх��b�LQyHc%6:ڃ>�#0�m[�U�����W=w�*�q���j��0:��GV;�ie�Uo	�S,�E�,�����v�6�Eɋc�,�Tй(VAE�I(�xX��U���yR�W�c���gV���6�̐A��a�>��$��Λ�uޭ���MX�%��0s�t���i��
�̎�d3#L�����]ΜI�ls�����`��lj��G�L|r������PSyOA���af���q��/d.���}m%�0��_'m��L:*C�	k�|�ٰ�i�+sM���.�Ma]���c
��Et͢�ʹ�{�RhZ�k�WO�0U�ʾ�
���,
H�"�q��*����:��j�W�ic��H�k��{ڪ�P[���ua\�.su�[��*͜p�U�3�o�����~v�-�2ղ���Zs﷏�M�0��g��O�~�3��)�������5@�b�}���W��|�4��5g[|�w��I��S�[��~��<��,�qx��{�j���*��ZmT������K��oG�m�;���7�I	e���}V�܁$[_`�i(]������K;�WGR͝���k��6��}iP�lyM&0�(��6�[�����k\c����\�����Y�%_S����~s{������Y�c�ù�;*"/�$��`5���p_�L�"��u���Ց.���Tu�ٷc�?E�;.?�/PG~KG�ȩv04�W���>�v2X¯�]Ƕ,���%�F*hf�]��.��e��ϗ*�֘2o�����@�K��ʧÿH5��6�����ٰ([�EOO.� �0�0}������=l�-w*�9�7��i�ez��Rsn
I�#�8�F���Ȱ�qðd��'�c���{�ۻ�ǦIC�ԸpG��AY>s�a{�LS�V$,��to��6�oL1�7N1���k7�h�{��)m'di�����+s�1�y��C��������O�²����8&[e��9|�Tе�E?�*����"���ƭ���x�� a���V|��>Y����1�MY{�U�#kO��~���f�RY��K2�ךn.� ��g����GbI����+�+2��4��y�F�/wD<�c�sll'/�,y,��.�A�M�FB{�nNX���'�F�ǸMU�:����a,��k<����f�Pc31��+h.E擥t�56�0�+\��w
�2�/������ ��vkVe�=��/Weށ��L��� u�
�k��R���f�v�L)�,�4�3�,�$�lu�4ĸ���m�Λ���l�#SX�tCd����w���)S2�wᮤ�j4��g0���J�e8+Ͱ�%��)L������:�����6yP�,K[KL�h�v�l�H���&�V�l�9�M(�n�S�qa��Vyٶ��Z��i���`ڹ�hD�52+�,2ز��'���b�͋nyW����7x�|A]CWwqb����_�V�C�Uq�Œ��Pd8𹲱9zH�N+b����^,��z�����'�{eZ�.�L�.-�liۓg�w�
:�a������U����]4F4��N`�hIi����f>�pq�a�*����5����'Y���Y�'�;�9(���|���g (�-�1;2,/��Y��v"5�3���֝�h5Բs:>W�奕�~%4�,b`_�n;1hL�4l;�hd��4�����޽���d{>/}��{� *�n؀�a>�2�s�{ ��\b�} �T�@2P����͒�[d�γ[>d{x�z���G� ��3�3�^�&ܮ��b.Wo-�>yM�nl��FY���3:��V^�����R�^����@%�m��a��z��;�A7fS)������%}��֛jX5"Wn�M�e(��AҨ��`�s7�l|K�5�S�wƦJ�U��mM(�l�b�q�k�9��D�/�s &��E���-(_���E��Ċ?6i�yO��B���p
�~���oXQ��(�86S��͎��Tq�˭m+3Fj�CԴb��@FX����,w^���=����T����_�y�����@���v/7��'���=D0�T���/zdHY����6_`ഠ!��+\�����!�9BCW�5ڵ��!���m���X��gU�jAPL��\�Cs{ �1��)�B�	�#�Xx�Cǭ�H�n�C�~x�bh8�ۑ�)�RO�S^)l07��҂��$��R���̂�}Ӣg����l+�2q��3_��Q��C�j���Ml�?;�VI��m�J��˅�M�(*��d��U�d؞0�noI7⊠�`ghx��ᏥV:�v�95�:;�Zo�N	�6�����Ĺ�f|�/]ó�Ƃ#+e����U�|�_D���(2���C�Y�h�+��閭'B�Tѓ��0н[�3��<4�����t��_ܐ@�0�
�\�pt�0P3禛"����<��v<��@��t��ǖE�����E^���V�[�.8���4\������d�����zV��-ڃ�rc~F}�b���fb��n�<�E0�
R&�3ه�8��zUVEp�p�d������f+z!#i�%�Hjm~{����`�n2����7�w���Q֧^�*�����Yd�^P�yv�c
�Ejt��"�L��^�{�D�ױz|#��0�bɼ��Bփa�)F2h���e
?��k�'�0+`0�պ7���k�ӁMle/�)�k�n���Xz~d^��}
x�:���M��S/Q��p�j*x�`{�5���9%�斨��7 ��Ըa+
� ��~�����U��c=��SV��߁�����Д��J���S����?���K��Y/`��,�`�+�q��2Q��]#����l�^3q��fN' �v�?�i�OM��F��G�R����ےf��#q�Ϗ�l+9�A������l@�h�g)|��-�!��X�@V��lۤeX���Ɍ�}�넗��4�;�/�x5(3�\�Q�՛~; �cNK���m����T6ʲ���t������ߠ�S�v^3����3xh�̴�����}��}fř�����w��L��?��I�φ�Y;��![��3$�ֳ�g�����MgO5X��Vã�}����3n�X��xƾ�=Sϱ��r�}��<�e����_z����.J뺤�Ʈ��^���J;rّ�#MG��z�#Ǐ����o^����oo���o�����,�]�]�w������ڿ��]���}?�����G:��v���of��.$x��>C�u�Q�yY�	n%%X{%��E��Hp?�����<�5���{<D��9��}�Fs�D�Q�ï"<�����TN��>1�×	����L/�0���)��܃��[!|�D�ߟ����d?������Rtm���ãV>��f�߿����������o�x���.��3��&$��lZ8���{�s~��7'��AxQG�.�O��"|��8�-:��������V����u��7���'��YW'Ə$�_Gg�[t�b·��s�F�_@��:�b�ߧ÷~��K�?��?J��:��ߪog·��~������'@�RDrU����Q>��]:���������o |��&|�����u�U�u�����?H�<������?M�"��[t�}�����$|��	���_�I�?Jx��j$����&|�!����#	�Q��#�}:�����K�Gux�7���o��o#|��x���o��/�������u�g@��E�C:��Gu�ό�������i���'���oM��1	��$�[���'����/е'��t�������KB��I��%���'��&�p]���G]Fj|�4S<������
��rc:�V�\�(�F�\("XIP���&�����ۛ9�S�w<yr}E)�	�vq��a�O�pQ���L���79�XD�#��jJ�^���8��Ϸ�~�7�|[	n��ҿ�ӉT����������+�V�����<�ƇI|������Fj�OO��o��4����=��+	��N��3>6��n�o<D0��������`�	No�A���}�	~J����Y4�Ί�G#�{	.!���
�+	�Np-�ݓ8��Y�M��Ƙ��'����=u	���1��I�KIB_|hAB:��I�GIϿ�Q�S�<������� ���?��7%=#	��<>���p��(~�唾��j�k�'�����N*_
Uh�O[��6�W��0J����5�q��~�D���'d�������ŷ�gt?��Ѥo��.埦T�O���8��Ϥ�\L��t?�W����4����Z�J��D�g���q�҄5����W�x�c�{lç��C����l��)���K�Ϡ��5�z���9o��:�����yT��Ś����P��?��/����)�
]��?���.�k����g��	¼����;�~�ж8ƿH"��S�һ4遜�[��ſG�{1�?M�(�K�.���(�2��H���{���I�G��.My�ǟ����{�� ����M�/3<�*�n"����H,R��N��@��M�xyď���U��u�|�NR�d?��(=��������l~���	�3��ޏ��5���t.:M��濌����8M�5��#���L�H��`-AA/� ��m7���CG��$����o|�����"�=�^�$�/f<��e� �Mp,����&XM�:�N��	.!x;��7������#�Hp+���B�m��'�.�'�<&�Ip�I�-+�#��`=�f�K� ��`���%���#�'�O|���|�`;��� ��Ov��`7A��K�^Hp�l�y�,&XI�z��o"�'�B��k�'x��$��!��]_%���{?!�9�.��	�-�p��"8���`���	6\N���Z�w���&��#����_%�6�	~N���	
-4�	'x�+	��Hp&�Ym�L�����	�	�����r�����8�lᰈ�~�o$Xt=�˴�RI����zN�s3��e<�M�ɞ�5��6����V�?\A��<+3	R9[��t�.$����A?A���
Tn�`;�l���p�u���н��[Btn �oy�3�0�t���HP��_��;�!��y�����T��?��ۧ����c����� �g������ԏJ�#�~�Ͽ��'�|ە�aQ7/���]Do?�w{�s����R�=���17G�Q ���1���#�AP8A�q+����a?峕����[�3�S�l�������!��~j�ͤ�?���[�8�Hp�h*�P�7�?A�t7�M
�<J�Fi�o9<t��G�����9��-��+K�oF|Ѫ��c��Ԏ">T��ߴZIp3���=�A��.�~�H���_�^%�/��C>�[j�C�t���A�۽��!j���_~��h���R��"ɕM��p!�W*����8������|�����4���N�A7�S����������">�h&�%ɇ� =G��x��`ѥT.���T�M['S�̈́���t��Y*�#T����f�ۭ�D�n��;�?&R������4NQ�)��C���z�<4�ħy>`�q����>X�,�|7�'���g���N�)��ߥ��g��������ґ�i��_�.a�s���A�KH'�/�aD�ɞk�����(���O�z]p�z��mE��(�JFG_��tnK�έ��'�CcB:yI���|���*1���K';1��I�����rb:3�Yw����I��}���oLL��,ϡo�ϦӤ�jO\�GN��O�N��%���O���Q��l>M:�~[��~":�?���ȍdt�ի����=y��Vy^N^���C����9-:o�D��$y�'Ķ�.�:��˓�NQ:���O��}���ӣ�������i�)JB��9���eI�$����9M:B�z��&�����sC:��p�w��Mԟ&��I�H�I�=	�I�$���M�>kO��7~����:M:�}I�����ӥ�Ln���y���������8���N+�y&9���P=�Ap��fy~*:"ͫ��r:/%�����Y�>ҭkfd%�7�JFg������Z:":�/��zibzM�NI����t�=M:�U��|p�t�$t>=M:��t���Y�y>I�9M:�����i���[g�|z�u���Υ�Ig����'��lkO�ϳ��Q~��%����J���	3ȿ�S����l�c^<��(}��>K��h�L~���.��ɿ�Jp#�M�����?p����к�_�A�9��ȿ���o��Ѻ�Z�{*�k���/��F~܏��T�<��ܒ�������!��龋���'��,=�	����J�y���hW	o��3V)둴nt���/����_���8<t�Gd��.�o�O��p(�N�u'՗ʝA��7��)]�>Iܟ�O��)p�ϩ���ݴ�1ѡ{��6�|B~������>�����~`
�oW�yO�L������۩�`׍��֣6˴���ֻ�����wr�Y��R?,���B
����!ON�W�k���g+�.��k	n$�NPs85|r��H�޶��W������"ᗄ�~����8��$��tt����ԗ�k�_�/�W��~�Y��җ���N��a����vr�S�|���-z��ߦ��A���~��_�������'��z����GO������x��s�{z���Hמy����t�����җ������[~��ߣOO�*�r;���qS�Ɨs��~��g�������y��/������W���wǏ��7�������O��7�������x��E�o��/�mz���5I�h_Mʷ�����>c0���S��38t&��H��$�E�?�PZ�eYߺ���n���#������J���u������?����*����[�$?�#ۚ3O�����!�v�}�}���mW-����;[���^���=!�`�Ơ�u5�%��w�/$��1 O�����%�WB^���y�Ot��q*���`�1�����c%��{ܒk��p�+g9���:���A�l$W�$�J]�5��{\BvN����_	!�"�o�Wt�����Fxd��R���=�h,��R-���*�or9����� 5&KVJmD��	p���� �&4����8�2���`��>�
,�n0�vO�ew.}~�W���㫧���3���.13g��ʀ�ٍ�1�e%�v�=��+�����P�Lr�E�v��q%�z��.��렣�Ihj�	"��K�K`�?�N�^��_��O�0e|ބ�S'M�2e��<A�]�-B����� �� (\B!�����<�\%@׺��j-����!����/`,\^��j�{�0���| L|�C���
��	��0��3w�f9>�	���j�ud�&/Ҙ�)c�O�'L�X0mb�X?��>~�}���k�)�ɓ����]'L�o�+(p��O)p'���%�B����\'�n��%	����K

>����%9����y��|��k6CxP�j�:+ ��yT�Hj �g �C��%�%x���b��T'0 TX��4�兀�f��" -��C��yX�r1�4 ��*!�����|���q���� �p݅y�9���K� �5ׁ��¶<U����P��	�^�H�3�%�XUa�K�~w;��U�O~Gp�j��A���8]�s�\>���1F��\��v�h���rT��#ç���[N�\�4� ��`���>��O54ӵ:�l�/g.�����n�_'%}�
)�qM��ϟ��X���G圗��/Bؿ�<aw,<�3A��ѣrS�Qy�G!�0�ˣ�V�u�������Q9��_�������_q��(����5�&����A) ����Fa���/Aa�)�#`��x�8��E�ǷT��@KA��Đt���T\1��ٶ��D��Pt'�M�p��+
c�1Vo�p���]>�f��Pn/�@�J^g�)�^�#_!mv�<�`�p��a�5M���o���AE�w�9��G~���;�:pO\���٬����ŎUZ"a�E��B	���r�(�AP�<˦��H���`.g�X��)z} >\�=���&W���nr;��Љ��c	�V���B�lF�@�U�r'-�f�"uh��`>����֊r�펊TU���F0ז�+kx�0��Z>K�1�U��cj��fQJ*�*+����s暫��j1�ɨ�
�,�V��+�bA��zO�R:�= Z���E1����CR�/ s�SP/b�ݣ�� B~h(�6��A���+1�Fa@E��1��5�S��b�:�`@�CAkk�3��Q{��D)�r�� 3�1�.1����n5CW��&�x�1���	�9]-:�P�ݻL�\��Qb�"t1d(YB`|��#��M���)ֻ࿴�������M#Ϊ��[#�%���0@r��K��A
U&ВYz����	��X�{��i(����g@v��#�3��B�7����dKS�e���z������l���c�<��Uز��j���쓑�~y$��{�ve���W�`M����,;�9�H�SV�Mف����p `�٠����`�4�끿���X�-x���n�
*y2c��Z*�<�Զfw;���S���CjAb7t%�]*�,��Nr�3�[�Ufj)֤A�"'��f4ơ>�"�����9�sxg#ڹȲ{%�'���.��{�F2X�`����g?��Ǝf�Ɣ�i���/�`:�1�Rp�zB�P��+�v��K��\r�a0�����^f����;�sN`F�q�g`_c}��r�s7z�E.0��`�Ap5�z�u ��\
)-l2 �%�jD��e���/rl�g8+S�N��O���Ȭ��~9��^7�����j`��b��:0q�2�	]ֺ�;w�=��l�\�r����[��_^c�ۖbWP�2���P��<���fD0�لK�ܨ����l��%A��R��!o0�������&�sV7�&+���*�,Kc�R�PĊ�0S��+��1�I�+�T��Z=(�2��N���np��8�fb�e�����b\B���K� ���ƪk�|c�w�迥#�nA�����N^�����b �8��1���0�`�N2�@bg��q;p�η�X�yQ�1R0ٛ����k��j��>0�J,Bu��\�fzȌ�s�j��L�`ׅ�r�8k��\�ٔT���c�[SQf�����q��c��ƪ�ѦOTYe-���b�rs-δb���f�Dc5���X~-Suf
�B� rU�R���(��U5s!CN��뜆��c~@��� -%�%�(�U�ȹ>kl~^p�#e���R.qR��AG�8��Df=D�7I�֫ L�.�qĩ�Q;�5��d��v���$; %�I�@cT9��I�J+S�ťnԸ���!�^'�����vd#��I�ۡĬ��C"wp
�tXZ9�K���\J9 -+	�-0��`� �Z�~��}̦���W�2Nv�>\� �46��|�/s�
R�W(�q�&;3�-`hJ���<�Zd��?��x�G���=�������	��� <a3��A�`���� �˫Qlt��X���XM=�p4
5�+Iw�u�C�E����Z^RS�E��,B��2�c>8���iG�
d���
��nq�}�&!$9PY9A(в6+	�>��$,s�0��	0_`�xC���"(�k��d�������y'�k��=Wqx��c`7���f$���P����U8hi1�
t6�٬טq��e�(VBc��\8�{\-J:3�(�f`�l�i�Ahk� ���+�*�ftىy-Y���=!��/X���� sǒQ�-��L��+�hx5��l���Ώ���p�V��N@ĔBT5:��z�ב�\�������k !a�koX��7���aK<� {�LS�2M�JCO�]j�9;_��b�1�Ӂ�7DK�� L�����r"�+�����QY^[��,����ӨO�g���_��W8�� g�0Bs����ߟA����O�Di��ia(NB/��o��<1�����4����V�g�� ��0���s	�j�U&��^��2��CZ�@3̜����k�[�ǷF_�ڭl�Rl*�l�h3(�� ��x�h�ܜ�E`�0�7�����Ҋ9�F�B$�"��[�b�3A6n n����%4z� ��iЬ��(N��0�|n��i������G��.\���(�}(k�`G�8��=���@���=��O`��1�C���nxt6()(\K�BC�î=��A�%1�vnv��:�dw@�� 1(O��*�z\������bRЙ6�͑cr>�����j��O��6�s3!��:&�����p�=*���~J{+��wǧ{�=
!�+>�Q6@�X��5�~7��Թ���i�� ���ƜP��꘡֯V����pzlF��W4��FV
�T�`�:4��ǣ�ϙ遊$��.�Us�rb���(�c��#qz�c�a��3���P���N ��вY ��%�:���`;�3���60p΀�~ɇױ��j�#�t��4�6���*@����JZF�%`$��.U�EC���S�W�������O��C8�=&o������8&�BX�����c���v<�N�)�q|��oՄ�= �_
��� ��9FD�H�XO.��,gn�3Gl�I�5��q��m���Sqۋ�5Dd�4Ɓ��*`]U�����U!&�#�%]%�����(�CA�I�r:N��@S�:��)�X�.��&�� �>e':\`Y��*�2`=�������8�����Z?}�s�X�i��Dk�Z�5R��u����[�J�*ό/#�]�����+��
.NC��C[mR�+���Ҁ�Y��`����
$�mك�ȱ�-Ea�h�	cns�6��*���C����|��ꖚ�D��1�9 �F��?;z����8e��y�T�OP�����C�8t߈��W_P/؏9WU��|�����N�@�!;s����{5�sP��f��EZDX$�5m3V	%UUf���ls��dnO�@J��F6�2��;���Se�V���sw�3V�R�5��a��f��cz�1c{e��X��c�k���%
c��ǭK�Ӈ��yX7�W>�,����!w\�}�T��찮������n�{�2�ϯ�7tB�����D���?���%�gI�<��+�Q�+g����y����N���5q�N�0m�,s3-*1=���3�!��c����խ�)�#����� ��r(w���F[����&�z_�׬+�*�R�\���Q�A��'��n/��3��F��'M�J���[|��MZ㊇3�9cnN���.�&����B~>�D)
W��׭g��|2���7h��r�։�vS\M)�d�1�Xb1DEKC�V��¦g��!��c�o�e�����B�lr�X�C���+H��7�� �Z�:	t9���@jǖJ��X�(=w��5�I[( e�f?Y���h%K�5��F)��(\Xbw�B�u���j��+d�EE��Z���1�
9�k�-��A�W�ǈ�slZ�_e#��ejr�6��g�m��H��G�p'}Po�7��B���C�4��r�w|*/�"X3biUE�8*k�(\n��l�	����E�ݍJ�d���M��O%_2`z�?�&�r�__����&@���/E*���Uà�����B�Q�yn��d�ܲS�hJw����Ug�c86�,���v����R��<�Z>]i�Q%UfPgH�=5J\����3� 7b�(���E�A{�P�G؏#f����R�(����tB�+[�����yZ>P��U�S�+i��{�C9�\�(Q���r+�o��n|�I��_~qd�Fi�g-�6�bk-����8�\�؂9x;JQ`G�юN�p��X�d�$��~2����OQ�����m�_ En�϶ߏ.`�N��K\�x:�j�@���S6�饟�o	zU�}��6
7�6����R%�y91�W�Չ���cDa�*�G	�]n�FwA�(���تL��_�D���ʏ��C(O9.?���P��������=����3��>._>�|�$H#A4�l��函�ďz����s �|
�.�N��A܈/z�
+!͛V�+�A��I���|�+��+����!D!�9�+/��B��r��^�����%�@���?a���򌃠/S��[8�+�~�W>�M�<����Pq���<��� �([#�Yu},I8��|B	���^�6��^�Ewt���a�W���_��!��C�j���zi�<�!�8�k����y��!��'SX~�q��p\A������ ,���.:.�.<.��	x�}�� �1��~� �������!��pp� �C���gC8�2���	�k�W6 _Ӂ>�ѻ �<��?��T�qy'�� �Bx�����ld�ap���5v|�/�x0�gwZ�A��bzCJ\��4B}�PF;�����PO�i|�y�-C'_'�@亝-���֜�q��	����f�����|R�VⲅR��d�� &���Q�o����t꘢{*��q[��yQg�Ķ�VWȻ8F�<�l�S_us�����P� WJ4�J��)R�ʂNR����*��~���p1�R��:A4�q���e�VCO��=���,c�X�!K��W�l0k��=�?�;
џI{e��.����c���}�� �E�<i҄I��`��fn��Ʒ�)���.hҊr�Y��.n�-�,]�OjhLk��ki��Py�e
�,l�"Tq��[R���H�蓇Q�ׁ�c���A��A[�m�����߷���1N�÷�b����LXSe���� 	��ƭ3���Y?�ˮ�}����c='և$M�.E��A���'�n���t��c��������`�ְ�J��d.5ε�%����,T���&%5By�h,�a��kJ�
c�j�0|=�wP	8��U9�U�k��+������	y��o�:�)�y��R���p�_:q�� eo��g��-A�����!+��s�aI�d+3�Ҁ�7n,%\���国�%���ݼ��Z�u�N��(s�0�;�={{������K��E���>���&�.@.��П��7:<�"�2��%��6 �}[p!rCQ@w����"^Q�W��1=��6,�ĸ�[hķz�=��U=�X$�=Z��WT:{��<���c9s�B���wcxiiiɭ�\ڦ}����c�"}�e��s$���f?tx���uDVD׎ �f��	�6|��S ��Y+�p�/m�k��\�T��&�$���}���}�5�2���������&���^�'�_�'��'�@x"�O�p\��p�\�'?y~��If��sY��ݥ}rå�FxT���}�������CXᖟ��w�s���� L���9@�_�٘���+�I�����q
a	U.6�[�XZc��=��Sf�ԗ���.oMZ��'�#W��W#�X��*{���idV�0�$�>��� ({����T��4p5��jP���ї�3���b�}^;��~o�T��8�كA�Í������RS�EW�w�9W��߯�qAkׂ�z��}&f?q���<
i�N�!wQ�T��5�M�����̮<����B�m�7�B.�&���	.[�Y�o��A�4IQ!R4>X�5f�	��4�)�U,�����r�8��d�1�2������T�4o��q7�����<'�=�#�r�Q,��Qi�$�U��#T&�q׫���p�_(�-ow:��7l$�6e��&z�@y��?v��Py�4�ɹ�ָ��!�g�������X����hM����	������YN�z$�����{����>�����&�.�0������pp�C�F��$Jw��O>a#�[ ,�0�7�ʇp�1z-蓷C�3��@� a�X����b�wC�ڳ V.+>qW�{��8<������ ����c�WõUꓗ���
 ��D�?��
0i L����8��M}����6��s!s��PS�<BA#��t�p���i�����/��h�g6�p��O�����/���!ThTA�$�!�[���# ���-~�羄�1=����7�@X�v�p��������u��
!L��j a�)B=�i^��>��
�Ū>��s��)��gsb��`e�zqm�����}��������R�,�ύ���6Zi=A��scm����^���0�(\!�e}�N�)�_�B#�9Z�'O�{���7�<�W?��a�k@׹�?�����v[��	�]3�~�-��-!T��u)�|? 򨭈�T证�9�'�B�Q�J��7�bi�����$�}A����������>�=�ت�@��j�����\��J��s�zHK6�]��R8Wt�\!�}�ӹ"���-V��\��������=E)8�jѾ.ݸ�]����I��x�|u3w�~_����#h�A�U%SX�����@��A{Pu��=�S^A�u�1��f�p�Q�&�4MU�T���UGE�S�ͳ��k�ћ"��x"�K�ÉW�N��i�Ag��l#b�q�TD��c篳����a^���4��]M�0��@|��~.���<��YA�z�h`!�$��e������+�7���(K*�Km֒ճs�pJ���_�ծ��~�o�g�ޜ�5�_���L�g�S����)/{�K���J`��W��w��ouT��Zˡle��l?�a,��ٽ�^�Ȥ���!7]���tE|M�bn��Rx���!�m����5G�P��\z��8�M����\-���g�š��y|��[%˅;�E5���Ҏ,���\���6:X��|�$N��U׬G��Q9�N�P�ׯr�k)�"N��$���&��Xy�-�&��������g(��0{ �:�ak�"v�UnOO�ߜ
��E]��5��υ�lr̶j�>	�k�$��y,]�g�.(�l9g��|%\/~���m�p��ul�h��f9�ʟ
e�Z����	�}I��jB�8���D�+��VJ��v
�Hۏ�I�"j�h�$vO�O��?1')K�;K���o-�;9�	q������W�K�vy��Z�����<�q�#$xi�P�t��
��N��z�={�������J~�؟u0Ɵt/�:��/r���_N�"8/� N4�q���Nů����y5>oc"�	(ױ����(m�P_~`(��a�k��5�ل�����|��$y&���N�`�H�;�0
J�K����TFU��M=��5�A�v��$ʛ�K�N9�U��N[e��K��W!\Vv,r�t�.r����\�"h�[�a�-=ݯP�8+F���s�r�򫹪�r�|qm��u,�\|?c�+X6���\"��&�-C";��.�bs�|3����լy,)��#��!�nG�����v�8���b�$g�ٞt���&�3��Sq����@'_� J���@��������1��G(��E��M������Y�������זT��E~z�����������(	�X���rWO��I�^*�Μq�T�Ŭ,��A���y����P(�'�=�� .�c���EuK�)�6���Bl����s��b���H)�����j�˯�������jr��	\��&�?�ǌl�>��Z��N��p�z��H�|.���UbbV��q.o�;��O.���*y��jK���rc�s{��m~4�xBc���/�W���-�ە�:f�Zc���!��>p�e(�*���}'E5e)k�K}q�k�/�D��j�8�
�R"wI.	�b[Eq3L4�@�OIU
O�.� �2�"nO�NUOE�)��g��`�� ��>'�!�������9=Arn��%�؄0��ϰ#�+��)?ۂ�lz�N2aO!�O>%�H�q�Pk��]��C�Ue�_(��9v���q�3���������a�?�d�o���p>��7}�������1��~�t���J&�ו�$��h��.����6JM�8�r4&clD^���@���x�xdV��dٔ:�8Ĝh&&������D<�dt��OZ�SĨiS][��ƍv�yN��l?l�3ѪWY^���^����_����F�ݙ�W�TēPW�K;n����!4H�	��G�q�L�ڃ��h��7���s%#�)��,��2w�����ĸ�"�)�Y�얱�YN�����-H�{�s\V�������QN-�<ky�H��5e�w�j��T��o2�81�p����$tPޓ6L4PP������+�1L���j
��}rr�����<���us�ADuD�1���X|]1�L1�N���s�-?h � �[�e�8�TYLU�y	xJ3r!��O�H=!gC8�OȷCX��ՀӾ�����m�}�l\N�S��KA)g���A�]��*�[�
᠎���×�����R��E)��Iq�bVPe\����w�$��iA��C.�yB�C�AN;yxq�̝��>=�3H���i�]��z>R��4��i�S]�$ꯢгY����� h�^��b�g�G�Sh4 -~z��T���9��9�.�=Đ��W�5�#
~z�|����O���̕ .D6�TA��Z��}��C�t��8�>�= ��=B�Ur{����m	÷7��Kf���t��a'�$�gq�1�\R��ٯ� ���������������"з�65+�j~	���Ϗ]��]N�~,�zBn�PFa?�C����O��k��u BUHf��"6�~�� %�㳳h4oqӎ��dƃH�x���|�*����t��L�D�G���/��:���XТg�d�+]�0v���|�ت���6�����\c�֨�A"L�^�U��j,�jk���UMu��sy5n�'lޯ�p����yꘗI�����\VWf��*J��U�jc�y������R}�QE������7 �O`��f��	~�����پ��N00u����L2����{ް�/�p�E?���K/�\1�̬+Ge猾*w��qy��'L�4y�Ԃi�g̼��^�p���7-�4{}�Ł�Z��e���oXpc����7���֕���޶j�w�	���[��q������_���?���ͦ�|�����~��c���?��ϛ�|��g���٭�m{��_�޾c�˻v�ٻ�W����o�m��o��λ���~��'���g�����+��e�᯾�wבo�����=�~�=�wB6\xȥ���鄒&{��[�
�g�s���K<;�b�:qGs���4��5� �0��QJ����j�/��;9���|�ָ�]5>���j��l�4GzB�&�)�s�J�[re0k��e���0�m��4�_	?4�2���ɬNę��E���ow =f>bX�%)இ���Q	R�[T$;v��8�r��F=������NH���|�ӉK͛����R�X����j������U�۱��x3���R0������oĳ���Ovi+�[Ʈ���E�+��U/�_Ny���sH��8u�Q{3_�L���Vv&�ran���2Y��"�y]��$���n�yX����U���I������ieU�$��I�yсB������]������8����~��1�,����;I�������Jl��6�6��E4���k(��(����QH��a�WC���~���y�ޯ��s�|��>�n����<���y�_�����] G3-�pc����LG,%�;{T�j���t�=-֛j��9�Bm�s2s��c�g��f�WadslA	�-���Y^��V�?6������

�ZA�{M��9ukI�Q+��Nѻ���ޝxT�=��`vq�3�C�n��sj�.�V��7��U	�����B���K����
��#v�w͇wG��8��C����(7Bd���\$�_�Bq늜-n=���6�C��H~$�
;���1�E��2�/�4�<g�qZK2��0Rk(�^��D|�D�DIC1ibك��@���u��ϑ�ɠ�C����8��y	2!A��zt�?U/&(`������{	�7l��3�J9jt��cƦ�΄����!�����{����=��3�����;�=�����kǕ�Ʈ��ˠ��w1ʬ÷3i��M��?��X������}��W����&铡8���~�Б�ǆZ�=ᘯ��OX:�B�OY��	�'�z���{W3.�ዜ59v%�]G��t8u/�s��^�O��(��d�����*��(�ݱy���{�k�����s:-�_|U��w��� ~���@O>�O-�_p~j�Ɋ����ɮw�z��B-.��܏�Y*� �Ë�	�r�r�}�a�υ�-����#��κ���Z/gr�4��ux���":�˰S��=INo8��t������"���q�2�8��Ȧ������>SN##E:��H���.��"�en�D�����$9B&M}@V�Lo.��^1��"Cd��/>-���+Y-u3$�3'�lxrۧ&�2/��]�DΏ;�Pڋ�(�&J�3����>7��&��DD��N���S׍�a�>_��:u�u�N�i~�珈�E0���u���Gԏ��2��)$�d��o`��k\�IL>�"}�����qB-`"�eC��f#-N�����"	�Kz��2@8d�9�:���钡6��2�-r�,��%(w�=��*��\���B^����w�}�H��jo�^~�_�W���ö:ڴ3q���aN3L�fR���s��b��\�o��Ef���\i�6�f��͔���!�����n�4o��̇���g�0��9d��c���6��ڀ�p���c��w��|?�{�Q��Ѝ�#������	�)�·����A��~=���X&��}ct4el��oc8����?-�{�!)�Ǝ�Y��[��+�B��Pp�h�c�Qi����ɏ3h��Х�c&�/�N���ӻ�A�{�SL���QD2n���nit���=����z������}O�,zn���m7b�����km��v5(e���o5�G�I����O�n��U�;.�nƻ�6tiɠQ�[珹䛢��N�C7��^?d��ck��6bd�شA#�����?����k���_��ˆ��G1V+�}_�E�{j�@cF��]��=`!�X0�J}Ĩ������ٟ�]�)->��Iv���v����s��\[����gL��iu�5�3 w�}z�p°�N��S�+Y8�7�ߙ#����ޡ���鍓;G.�����8o�e�\�����Y4:���u�$'O��Qx��S��o�ri�)��(�d`bBqm�å	w�����VN��]:;]մ�~����C�?1t����jW7<_���@�L�r���CZu1VNJ
M�rںg����D��j���%�Yd���RZ��m?�e�����n�f�f�����0���d���/�/�fړ5�t�|���ie�c��,6�:e�-;��@�d [��r�����O���e�lߑ!�b7���j����6����O-��e��/����fӼ�W�y��e�Y.�e��i&:�S����\R�+�ڬ0Wّ�2��������w繃}���m��i��=�^얾Z}�>���������q�a�ڽܽ½�-!�wܷݏ>�6
�n�ih��y��ﴢ��s��#�uv�\!��Y�y��,e�5M>�/k�w��/�g��ݥ�K�����w�;�}�=���ns�t��n�������u�rsW�#ݮ�e�-�En����.q��^��&��	�,w���Ns��I��n�;�Mv�����>n/��{���������|��p>�%�9N{��V�G���V{�j��(��^l���K�bS�^m���1�X~�y�����	힯�[f1�#�w;��yanAu���ؑ�~�A'��������tt:9�N���Lwf8L?��Lp��i���a�?��u�r�tR��^��������s�I�Dg������	���am!��Y��������O����w�w�O��0��ģ��v�m����;�3�cNC��:��1��644t�dL�4Tǖ97y�ﴵ*v>�:��܋���VN�S+��e�ؙ�P�Z�tpN�D+�n{Ò�����n�O������־?Zl�������n=f�F��Qk�.��ǔ�=:���y^���3�A�_FJ��5����<�<�<�<�lpwuqv�9k���e�B�*�Jg�s�s�S�\�,p�;ݜ.Ng�[�ʹȩ�_�����dOU����v�t�p�;�9�8�:=�
쳅΅�K�w��,qJ���uNۮ��r�®���=l>�����~`ߵ�۵v�}�n�����������l��ٗ���9����o�wz�>k��_���g����d9Oٍv���Lq�9�۟����u�����i�4w�:}��N=��N3����i��qjl����4r�:��}ν�Jg�s�3�y����u�;s��N���d;Ü$�����Y�\�<f�ۇm�Mw&;iN�s�3�9�Iu;��@��C����=����O��q{����cog���ٛ�R{����`K���}�m�u�Z{���^a�o>M��cL�Z�����}��Y�bc������
�s�w*GOk���QA�b3�L���i�sF7�ޣ�E����꣏�cZŶ<&�G'���~'���#sJ�,��y�Mgt��*�Ulzl��/~t�`��+%�X����̜�<��;�O�^�\�h�{�����Չ箼wA��S�;}ѕWEǜ:���]�,���1��Jl彭b?���s�64����)-3�?Y��V���r���G/]vjL��%.g��1+No�2s����ړfn=qR�7��u�͌�i��r��I,�ؖ�*&X���`0�)CW�c�W���k��k�=��{�k\�����������.'��$}tb/<�xL���Z>���},�`�-����`>�u��=��b�c�)^���u�׮;&��G'�B��O�V�	�!������g�i�A���w��J�%����f�\��q��ite��[��v]�e0|-��	�8 ~:�m�vݑ!F�m:~b���̓Y٭H�ɴ��3���;o��w����t�^d�2&&�e˖�/�񦿛%�e�<V�����k���	��CN3�|��x���k�=[|�bEp�
<�,/�6��7�]w(H���A�i<n.�6E?߽G�C�3������c޻h����ז͂�1��[Ů]WݴY����݊����/�#M�~�`̊�=Hu��uɧ�]W۸�ѽ�<�u������/�ddN�f�2}�#���Z�f��k�4m�l�����׮�qF��H�Ѿ%���Ŏ}�Ń�6K�6Q�.i{q���+b����؈U�Y���Tׯ������nipK��ܽ��{nM��䕦�F_��2������I��~ͣ���h�E3����;���.�<�&�L���.þ*//��S~��G�8�������+�w��&�W��|���;�;�m�ݵ�����]��:���7��ˏ<�q�K��v�����`p��>��>/}�-�"|�"�v����~�V��`�M�m8Ja0�%X�T�������������HX�t���?��ѝ��r��B��S�ɦ�� �A��
�Ҽa��i���\l/���������?J֛qv�L�T�`ϱ��L�v�5Ǚ�;e926�8��r\d����ۑs�yf�i,�����Cs��1cd����9�[�w��d��gw3Ǝ���p3��5?��Ԗc���\���T#�rV6�>�R���:�d/���\j�K�S���c:ۺ�l{6��5)�f��,�4�ҺQ����H�|l�P��bN���\瘩v�mo7�|�a�d:%�|h2���Qs��+��7��n��T�j�����,��{����?�V;�����,�3�\7�T{�̕�e���D�迩�������Ԟ��q[-��w�+���b+e�il{ڇ�V���Zce��+̩^���[�.�S��!��\;����lt�Т�i�Ti�7}�w�%j��v���\f���6�D󦴱+YC.7?��I5�b��ڌ&�4�J���6.��l1c�xӓ��$���2���k�\�7K&x��<K�7�����\iV3���z���f5e)!�43�n��6��t�%{���<bn�������Iv2qw�>v�m)9VKw���~�6bg�`[Ƕ4��M�����e��Y)!���3y�
J��e���.�z%�j/�%vdx�n��W��d-��f�����i���-Y3bn�����R�f�����,W��� �i���uŝf�I;�������(e��([Iin���J���A#lo��gG�^~8��G���!�K�|r��L����fB���uCE�P�1�U�f/����ds�2��YΥ��B�'�f�m7��u1ߙ�R�^f-S:�W��6��7FS�\V��I��\m��V�1s*}�Ns����&����r�%�As�%�Kr9E�٦����4�/��J7�E.q��2���,��3{���c��; �t��:��X�����ٓi�,�?���������{2þF.u�n��T����)����0w�GG9ݼ+5��\Rd�92�y����Y��A��r�qd��-�כ�ڜd�V[�n{x����Xz�[���M�<{���2�`�1�6����9���ڡ�(�)��C9�N��^dFș�D�]�u�Y�ߜ���S:�\J��S&�k��O��d�W�Ǩ�4�F�B�e��<��2	m��m#j1��H�F>7�噣�|j��j��!y�Z��+e��kN���H.��~�ud��A*̓^[\"�V�H�19�j�E���m�eM1Ų�̗^�~ P֞��]�f�-��6B���ig^�Y�e�b���f0y��v���d���Ws����'�l��,�~�]N+U�r�}]���%�|$�K#��63'�8e�z��2���k��2��7i`�ڟ�J�d���'ML}���W�����f�������.yX>1W�D�ɜb��6�h���s����d��d�2%�ϼb��B�T��Y%O�/�j���	�o����fO2�M�-���KC�����/1��F��;��> 3����>r�YeZ�L�ڜh��~6��[���m���I��=h"��&�|#�{��1�d�^VL��*��	���c�3?J�9 o���~�\�I�ia^�����؟͙&����|S�Ƙ��O��nì���O����{G7:7�M�&g�Y�����-�f�����p��U��̷�����)w:w�;�v����ǖ9ef�s/KZ��D����������YeW�C���ow=�<���݇�C,�G�����qG�',K�	���� �{��m�t�4�c>e��?�c���<�ZS�<#��g�����s�,r��̬���f�E�"G+[�l1����^��_�7��U��uߴo��~Y^���O;�:�%w���[�-�������m�m�����*�:{�=�a�:�W�g�l�;d����p�El�mvY�����e���̇���Yg�9k�?\�[kֆ\�:�:w��c�*Se5�:덻�>2�u������������W|b>a[��T:�fY���g�<�l�mr�%���&���ң���}Ь��|����u�K���g���J�r�������T;�ʷη��7>C�FR�X�|/����wB.���e�Z��ڱ��1�'�sPқv~1�ʯ��`_pE�����ײ���֨��BJ�sSͥ��]ͫ�^�����h~��8:N27������+�3g�����=�=N�����q:9�󓭴[��;�m}���|;َ���l�g[�X������7��ؒ]���˳k�2͛��o*O��|i���Υ�R{�s����\'��qR��Y�Nsg�����uZ9'8]��a6�:�K�^��}׾cw۷٦WpL��E�#��~v;�:�N����k�;����������Z���b|'���������s��/�H��������j���O���C�����{�[��+�s����~�~��~�o��o������ϸݗ��n��k���+�V�aw���{���}ս߽�}���]���r�s�q�t�w+ܠ{�{���]L~ԝ�s׺�+���M�n��̽ٽ޽ڝ���^��ӽ��s�s�,7��rS����%�n��׍s3�n?������sǺ��y�dw�{���~��s�pz�=����˥��0w�^}Y�/�s��+���a�U��Gj���n7������fվ�DG?E�6��~��wKLv���3�tz�S�����/�{��_�j9~�IG!zՓc�kA�'t�^Fjط�&N�D�ៈwa�u8bg����FE����㢎�DE9N=�#�I���(/ו(�&�qR=�7��9r+%�2^~6ʻ*3"��8|E��L'�I`Ը���JJ��N�?~fʏ�IZ]Ibkuȋ秈^���=�O��ԭ[�Nd�����|z��WP��M&3/<pP����H����F�qu}�����n����9���2�gf�eO+ΟM��7=赒��feN-�/*�̂����W�g��(=�}�Az�{�o�(���}x]z�ނ�WD�{/w��W�ެ���ȫ�5�i������g��b}��l��.z��1}N����W~�f?�-��ׁd��d�÷o��Ȟ_$zu���ЛC�k�~-����zt���1�Ծ�1�+�����е��jT$G��<�f/��#���F��׍��'��h���s����gN����q���43s^�wK�,GY�R�t�����{U�+rӽ[�g��E��_�~�����6J�v�,�n�����Ez���P��_X|l݋r
sg�H�EoQ�P&T��E,�����G����(�\���o��\k"%�m�$� !o�.��e�~�H��@��O�����ot~�TV�h���z��\�x&S�:F�/sj_���z/�g�x�6�v�	�Q/�Pb�.TH�0���.��N�(ɟEq2����!������Q���+�Ee�~���7�q�HO�mi���+�]�rӳ�el��Re+�oiK�Q�j��8�-����GL��v���Po\�YDg�ޘ3R�����Ee���K_����h���^FP�!�᫣%yV֑�Q��217;/K�g��(m���tFe��wB��c�{f��>f|��22N��/�/c��c��|L�\���f_(CÏ�H8�dPVֈ�3e�����d�������=.�/C�yJjv��|ދ�CΜ=�@F�E�#��z`��yGf���=�HB��6C��g�z�Մݘl�<}D�<�6�(����ܠ��zc���l�Ë�[Pc���ѫ�X�Eٳ��C7���U4N_-;6;{FJZ���
dq	?KY��Pʝ%���e 49����\�"s�x�SQ�-��Ȣ�P�KJ���mT,J}��-֤ ���ɝV��.)��x�b����S�VR�����͗��9�Y�dz�>D����
'��$uQ�:K��mt���u�Z�v)�ƒ�JjpV�|E�(�jh������gIu.��k�r<�¹��͓5�F�?����O���*6$/;�0T�P��;�����>-�0�L6�cC�H�Sik�|6w�T�_��.4�ڰ��)��z��"�P[:伾�^GJ�GPW�;tF��bCg��6)��ߑ�3Gf�cH�/�!{zhu�&&eO-�5��5#��ɠ���g$��P}	�����%y^A.Kɫ���&�g�k�Ƈ�|_�r��`|x�m�Ə�T�c9�?���ӧ�*�6G����!O郞}&����]�.�ֽ'�x��:��w�>L�@�;>�t����g)����e��5?��$�P\9Ct�%z�j}1?;��8ј0�ǍK[o\��>��������Xof�����!��đ�-�'��	Ь�i�7�spG�͜�o�ҭ�l�UV�څR��Pɡ7�N��;GY�=�����F�����a��uD�ȝV��;|���C����ြ��6|4:�L�^���St�gW�X��C/�=�Gj�=�>-̦�P��g ��v�~�.|ifhɜ3=t+�i�=�m���r�a����l�]`���;�3�78��i��<;��/��xT���[��z����x������E�|鱄5�W�Q�-Zt�ŁOd���FM/ydom|���Xp�gJ6�|Y��_�$W�0=Ӌ�(�\�ż�ʔ<��K���9��	�&�T�����v���/��:���9�\�$�@?u�ȿ�д��z)t�z���q?����{������;�$[>&��B�얆~�&t7&�4Nr�4��<Sl�3����Lws9'�W�xs5�^c:Y�s��&`�i:�Rgn`�&��,5]�ͦ���$� a��w���.�ה��}��YE��p\���M?�(y<a��oB[(��%�n�����-�;��h.2?���Ac�v�igM�~v�9���6��If~���$�X�l[����MvڛǸs8޾�ib;Q�����inop6^�4��<�^s\S�,1�;כ]΍�-���vL�jg�����������Dܟ������r�m�6d��ݵ��]�F��\Ӱ�5���;�E��R�`�*�����[/2w��0e�MFd��#���9"�E������_��h5���f��ͥvS���6Yfk��v�n��m3��_��c��	��m
�/m
�!�wl;�tj;�tn{��޶��huE[1����R⣻fċ�?�L��f��'���&bf|��?��ǧ���1��8�ѥ�lI���2޸�1�x��Rr�i�n�i�}�0�q/Y�b.]e�^�J�?V�iJ	+c��U�Mۚ�-����F%-%�u��t�8I���(�2LFK*k�6yE^��.oț�Kޒw�]yO�NFl\�Ν6M�=����v}���]{w9o�y��[�>��᠏W|��'-�=��5��\ZSRsy��5�5�k�y��񚊚-5/�l��VSY�qͿj����槚�5?ׄ�W�}���A�˯o�����3�u��:a�g7܏��t�=t��z�px=�/�'f}=�l��@��b���E�Idd��9Al�h1���Og��c8fh.�͛���\N�o!��b*Pj+i4�����{���X�CI�Ҫ"V�[K�5m�ݍ&�N^@���H�
|�b^[iUzG����^�l/���.�@�q;���(���ƞ,N����d���V��07�8q�;G�S�s
e8El�ɸۉ�$�`'qb;3�3�
�K���'�x�=�i�����J�(��v�yWq㺒wW��ޕ��'��n�w��w��adw�����L���LG�Q$g�{ދ�^�׋p�F��G"��3��Df�g+~K_�W�%�R'�4�9��O"*����K��ԯ�/1[ΐz=H����� i�w�4[�(q�X�ę�b�1�e�ԏ�2�r���H��R7q�G����$�y��Ys�8�'�o�d��ϣ�ϓ�*�7C�HgM��r��/ɒ��bٯ٨li\1Ml`���7]|�s�C9R7-WN,ɥ>��/�@"�.���I��<9)g��Z.͒��|q��Yi����=x!�l��H,��6Er�>�z����s�\(N1Z��>��R�H���ķ�].-K.���W��/��"ʶ�~�H�	�$b~)Z�V�L߷��]ɲ��v�R�_E��ROn�Q7�إ2�].O���v{H"�>*ΦG���(�}�>��|LF�<A�l`k�Q&�md;���gI�BZ*Ŀ�B��
qT�����������Y;^�6�UZ���F�e	��,'�mc{�
��l���>�7Z{�&��ڨM�Z��6Yq����֖��wZYfMs_f�,)��nTy7'��ƕ�X�w�mR��:U+l��J� �^ҹ׺r�m��>k筲W������&�o݂����~k������k���p� ���5p烶ޒu.d8��L��C3o�cV�w��~�؃[���R:����I���?;n�����i�r�9������zy�����8��5[9���m����O�p�$�]���k�fr[|{�jﲭpm�8�M�s��8���:���S\��xבD7�*v�T�In��I�+���n��C]��0���I�[q��%�i���ߏ��?Y����L����s$�o�s�&�Gi��f'���lB������~��V<受
VE��Q����[��7r7�%m��I���_��߹������������~�����l�GTl�ݳ��Lv�;�������o\��T����<�u���M� ��we��y�.���o��5{�r��/�=�S�f�H�jq��#�F%�Y��J4�����ч���ǣ��&:t���g��c?I�h���<'�_��S=&p̓���ɪ����u�~d:����IV��C��-���c��.�+_x�?�/��7��w�g����)��m;���ǂ�e9��Y��|}Ll�,aA�Y�=�ݛ��M��Br$+W�3�}��=�0[ύ3�8���n�D�4���o;������IP�d�+��yz�)�+(ʝ�g�����l��njvn�L���/��\��{���}C�kQ�9K���~��L��)(�ǄHAfV����T��:�}uQqV���;���3��ء�,�5�b}R��EƑ��o�����7��z�?��kJ8�.	4D[C���A$55��5��c9@��χ���ck����ӏ�����˶~y���?Zx㮑�U�xw�ܺtP(Zu���U!�qK���*+/���[���i�������s3�Ɯ\v���&��ڶNb8��a�_#�>><��gC���x����%��vxh�#i?�<�sgtߑ�ݪ�'6=���oI����O?���+W����QJWb�t�
O�*�π+�$�8)��kF�Û+�v����&����[P��;k��S���(�=K���3�0�_��᧵:Ծ��{�ϩE١c���z)?r�{�m��������n�u\�Tj�ƅT���(�����}�?����$ե�0ߔ���󏏊ߥ�{*���L����T)䬶�dy�M�T�_$jj����[7���>���>�KM| E��avݺ�G=��{�w]m�a�Ƅ�p�����<�9^�.������X�����J�0��ےcGu��[�|X�Ϟ��:߮YX;�_����)��@?ߜ��\��Ʀ���|�U��uor�G�0�T��\�����3m����7�]ߏ����?v�?}��}�1��A]���.9v���WO_8�β�~v���S������g�؎�x�*j�~�A +_R?E,.i��A#F�rd�>Qlv^��p�;bب�%@�Y��7�=d�v����M}�)���>�.����O�b�;����0.5e�ر^Ji�M�qb��E���@����G����Ӈ|M�)��P^�q�F%Ֆ�v?��4I�����,�;����}�v\����O	�
���d��+�ū~�9����&ţ��k�������O}V/媮+�pI�H|)��){*|5�L$�@	�rx�	"��	�:4\�oEӷ�UP����G��<�-cE���Tӄ��Ȟ_	�G�5>4�E�h:�e��:/�B[4�U�u��vk���W�¶T_A�-��T_}�;>
v@|����p8�ǧ�	(�sPO|����K�b�_
oG��2�
J�WO��A�W�4�+�d-'�՞<4}x1�������oG%�>|-�
�XӁ�h��?B�Zw8��B��uY�� ��� |m�y�%'�l�2�%h��ގ���A�W� [Ɖ��t�{� �
�a��~G^���O��Q3|���K����S�n�_g�ӆ^ԅv×��P1^/ |-�W��9�^�/�O��r��Z�/@k4M� m�4��h��ބ*4x7ڂ/�C��l�r�)h��/G�:/\�vj|�<ڍ��o�=Z/�	��W��^��>"��r��h?^�y��'�n耶'�jy���>��ɺ�=��+Q}|)������(���Y�X��c����f]���}X4M� �/��9�N��a{�	����e��Z��4>t9�(�t��h���'�<��0-�t�T�e����Z~��U��P�3� L@���DT�ih=>��6hن�tG[5\�*5}�g�i9�W�J�6���p�گ�pЙ,#M.A�^�tH���g�M>@��������l�9>ތb�e�����,A	x�7�?�vŶL�[P��s�H���J�j��(O��Ϧ��0-��7Q)�
�C����\ӇP��m��8�RӁ��X״<p	Z�e����~��h���q,-LC�5��*�<�F�S�v�2�'�^m���#�WM`�h�p5:�m7��Z�:�u����@y`���W|"�"�0��+�(|	l5�����=>Dq���u^X�t^x#�/�����
�ꏯ�ߡD��+�%i^�;��Ñ(E�	�TMބ�4}�$�����dM�M�nZf8�i:�vT���G�<��?�>�u���EZ��Yw�R|l��ZN�-��a�t��z8���J�_�g�O�^��[4>܁*��]�S�gL�?h:�7�G�3Ud��rh��6�b��r¦�Z�	��Zw��>f�G�Þ�,w|"\�b5���2�'�R���AIx��.M�π#9�§�� �,�I�K`/N�k^p'Z���3��7i|؎C�J�NA{5�}���i�~M�C��p���D|�b6��෨��wـb���E�/�Q�9��a�O��Q">EI�T8�g�R��W.C�ep%��/��Q���\L[i�p;��W±臚&��k]�Gh	�f^Bj8���p�y)�z���39�ܣ���_�ۗ�7��p%:���1y�r��P}|%���m> �X|)܂�5�����,O�_Ӂï��pJ��з�i�(�s}	_ w�|����/�@ӿ��뼰)��e�����	��k(�ƿVď�j|x"
j|x-Z�u�������h�-ڤ�,���vMnD;��p�?X5��z��:�~�����,t@�NB��StH�}Ji矉�G��r�:��W��QO��@�A}����/�_���j�;J��7R�e�O|l|3���Q��C�4|�O�A�:>
vDK�	p"
j`.Z�e�ע2|)lv+yh^�m��a���?j�p!�ė��n�=5}��px�r�J=������4�P�O����x�I��2�!��t7m�/��(U��Y��&:/�e�K�+h�ǯ��[����|�(������?N\M�Q�G;��5l�4>�}-u����h�_��U�6�
w���JX�aʏ��{P*�
�x�2��+�@�×���᧏�������Y.��	O���`Z���m�8��$�i��q�_?�r�r����~�/�_�f�jX���
_�?MƧϰ}�p�J�W��h2^��e�K�T����P	�����Z��V��������ײ��ʹ���B�5B�:���^ ?-'��"AZNx�K�U|܁vk`筴��ë�~-3t^�>�(�$��(?���m,� V���B�'��Q�nB�5�
%�a�v�> �M������>n@�5x-��k�sQ���5^ɹ��g�3_'�
׼�z�/����*�;:��)r��)?L�I}���]���x�×�gQ<��~���O�%(�q7�\��w�'�&|�鼰��l��QpZ�/����4&��>|
��yỨ_�������	h+^y6��2�+�n�/�U��}ʉ�ix	�ֺ���A���3YS�c@���9�9�>���+��(_#>��t^���'�,�_ ;TQg||��+�hCMވr�ep���'|9l�	�-����G���{�K�����G�ZN��s�Հ8�/X��lp2ډπ��n��|�z�y���~M6ޯ_֓ <{�^�[O2`�����nՔ�����/�W}G�������x5��p�ei|���+�g� _{`=��a&Z�����bM.;���8����N��Q���'�U����h9�ꀞ�j�0�����P��.A�5��\������n�('l�#�S��A�5����>��p7گ�0��^$I]�(Ґ&�E���W���_��(��W�� ����R��7�������.�3� 1��O�}#%��pħB���rM�C�:/�����	F6��j�E�a=���:/\��k8lX�H��ß�^��3r:�q��ȵ,#]�H$> w�(|%��⥁�A���Z�/�o���*ة��������a�(#)�D�M���/P��hl$G� �b�>�J4x-��41�����0*�8��fFVk^p`����h����ka5کe��b���g�I͍T�����nIj��(�!����%���Cc�$�S�t�_ �@��
�1J�W�>'�e���dM�њ��p� *ƗC��D��&l��A�>LoK��3�F�U��]��3�*��$#{���e�W� kO;h|�ҁ���s��Rwx=��/��P3|�5ח1u4bQ �@�5<�d�� �P>>�z�+�	qF�����i|x1��2���<|9<����D�Z���-:Y����x�
�
�U:/lօ�N��{�v������f�}�x��2���6J��4><��Q/x{7����C(/��ۨ/� >����`ہ��E(_�����S�V������M���d��q`	*�y�T�qzy�톯�M�җ���4�
�w���><��(�Uh�����z���S��VZ�"گ�§Ϡ�Z/�y ��r�W� �Hd;�O�m��41��O�Τ��(x�Y�__I1�_	�d��q�h�T�cP��F�Ɨ���نh�0�����&|\;�H���ǲ�����X_4Mx��80bm�e�c�!��"��v�w�(|%�5��9̋�x/��y�(A�L`����/�?��>�p���Ṵ!>
�@�9���O�Q��G%�jX�<��0/����K`���3�8>�v�r«3hO�~�6i:��L�P��S�?�2X����VY�%| &e��i��
tP��BI���i�_�
;�p.j�/�5(/9�gsY��0���O�A;�`�L���7�%�>�x}Fӄ�_hd>6+$�Ƈ��f��q`��|*|�Ǘ�+��O���yԥu��\DZ�X�����S~| F_B���']ʾ� _A9�J��2�k|"�-���c������Z���+�� ~�6h|��틦��N-<�J�MD�x���-:�i��W�\��Ӈ�Qp�5�_�kY�|	�M��uF�C9��K(�z�
���a����x
�Ka��iG|�A+���?��k���7�5>܎v�+aϛX�5췔:��{�ԣ}`�e���85���Q _��x|%��̶SP>>����>���i4_/�?�%й�m��w��*��m�����N[k:��N�5^�r렆�;P����v⥌2�*�磽�/lp7�����'/���]�R�;
�e�C��T�2��ᝫ��/�����*�b5�	_�F4��O�,G��z�e�O����/|�x��"ڠ�©kX��x�Z�e���Q_��~�:j^�G�c����&��Ǩ����0�	���8o���P��C��jx��Q����b�l�����(%
j�h���>E}�����`�Ml�t^X��꼰��,_�/EU�/l�,e�'��萖n�`�mH��o(/��Q{|,B	��
ꉯ��D������&�28p�5>6{�}> �G9�r�9������,w|���j����� ?D�5/�&�i��;��<m�g�m�R�	�A{4/8pm���-h��6z���e���!�K�ۨ��Q������mʋ�2��M[�������ߣ��8����h��{h+�&���
T�/���yZhߧ|vB��	�LT�O����ע2�nC+5������ҶZ_�ڤu�bۈ�hy�8��g�J���N���Glc�<p�����>M�c�-tP���H�Hv���->������N����K?���e0�3��u^��_��Ƈ;Q�ƇK��V�}N�h|���D�Ý�\�å_ү4>L�O5>l�u��p'���p�ה�1�a�7�|lVM���N����K����}G�5>|ehx��������?R|*,B%���'������u^��������h�Ƈ?�x��6F�-��2ڎ���j(7�6+{5/X���l����ó�`
�lB9�*�/���X|5̳V��p5�q�$�J">���T|��Y���i������-���|,�����㷲Rӄ���?B[�lpR��J-\��h���V�i9a�V�)e�3�Zi�/�C�Y�ǧ��'X鋯����o��KX93����������P�Ɓ���}���V��R|����C����O�J|lކe����ZӁW�ė�oPd3���JL[ʏ�d��
ע��rx�����d�n4\�a�i,#|,G9�@��*x�,#�;�L��3I�_�&��Z�U�+a�P+U���0�T�0���HN�.�gT/#h[��
�E�5�L����ᰳ���8�	�����SX.'�y���FRMދ����@�e�<���GAM?D��e�YFށ*5�0�~���c����i�+���.�Q|�z>�ޕc%	_�ie2^f��Q���Y�pT��
��YNx�F�I����l�px�%Vv��a�KY�5�\H�bH�(�l� �z��@��_X�
��W�>�hg|"<�J�Y=̹�J���_l� _
�@��U��5���GA|�{��2|	��'m�e�#�|*���kx?ډ/��o���Qp��Vh���M�����J����'�ꛩ^�����̃π�n��k|8a9u�px����2xb}^煷�M��p��2k8�v�Sa�Jʉ����|<�^��-('�DQ�x�j�������'�(�%�+a�)'>^�rZ�1���kh| ��}�
ǡ��85>l����t�T�q��h�nA�/l��rh�p!ک��ўzN���^i��a�_�=�vG��x��ג�a�,#| .E��e�t=��8���+kP"^���p�NA��X�&��9��R��I�q�
��Q1>���ix�lt^X�J5��@��	p$Z��ºO��G��h=�Fl��4�y�v�g�s7�>���=�z����>�m����-�V�	\������||�E�_c��&� ��eꎯ�/n���J�p;�&����~�*y�a��_Ӂ_��wTRfM���Y���r������9�
�������?d��π;>�����+��x_���t5M��{�� �`���߹�_h�>�}_7�D?T����2�7P䉔�Gb��pgGzj8���#)�j��:Q�q�.��G��(�g�|*�-�����k|�dG��+�Y�~�6h^��F�l���V-<!ʑJ�����3`�Ǝ��p8�DG�K�3(�5��EmI���[�Ǘ�K�:��/����zl�Țv����_�%�j��$���WPYk����Bk4��ޑ��D8m����h���E[�<0��#��Q0�#� �_�}�&��dGjy`�8�iC�p7j���;;;�a�SY��X�R��+I×�'Q���F�i��Iw�@�ͲkS���_�C}u^�h_�F�cᕽ�Mf�����tG�k�����#����3�_@��pX�������P�W^��k8�}�#��28v�#����$���	&SG|"L���8��0ꈏ�ˇ;R���:#���èG�����M�cht(�߱;�E�%/8v�#����_ kP,^�XGP>
���W���H"�����×ÁY�p�,G|	l=����[Q)��?�����.ʀVk��^ӄ�O���+�_�e��4/��Ӽ�oSX״�SI�fy����5o��o��4�n��o;�3J��t��Ǘ��Q
�
��ud>��:j��M������������5�;R�yͦ/̣��\��5>l~e>�4�W��K�j�/�[�O{��Fu������%� �$` ��`�KI�ԡ��!nK�%�J�"۪,��V'�)��@[J[�-�]�K�֤�@��ӛ�J�ץ�������k4J��=�L{���9��V�����{��~�V| ~� �E=���}q|�x��\Ԃ�q���@b���0�$p��	���#�Q��o9?��o�G��\����r�p{�� ��� p��r������́��>�'�ow�p�2�mݸ�� ���6���D�֏z�'���;N�:r9���8p����
��K�\�$��GP�<�0Q�������?��;��AJ�'��}��y��!�;�	�2$>�� �9 N?2���&j���ã�?��y6 >|���-��	��>
�s�s��?�o�G�oB��O�9�� �5{ �'Q�����n�#OC�\p�3�UNV@n� ��0��Ϣ�8��(��0�H�����'�K~�~w ����ޗ�n_D����Ͽ�v��{\&z%	�9���L��+�K�$p��������
^C����oB\�����p�K�X����e/|u�r���o���9N1Q%d<�+d�����Ip~�Ӑ���W I.��}��<y���� R� �D��x�F�yf�
��\�D��H�O��JT
��+�<�/Kt#x�f�( >ܙ/ѭ���0>y<\3W�.���{�K�Kt���r��>k�h��~�P�X�: �["��x�i���ވD���-����KT�[.��9�"������ϓ(��r+x��|ԟ���$��t�O��u�{��F=���s.A=��!o��F���|�ڵ����x�:��G��@
��R�����3^]�>�{���+8���$*���B��G�S��_\��6n�(��B��^�c%�� ~e����\#��8�U�����Z��\�F[.@}�/|�O�oC����_��Μ\V�w��%�;��H�>	|��98}Q��}I�8x��l�\q�DG��Q.����������s���Q��J<��{Q7p�6�k%��/< �Vp;�oJT���ϴ�NV�;,����8?�W��V�;,��{�{���K4����F$���7!���w@����.�!�����.D~�ޟ���`�1�s!�d�ꏡo�����f��9�������2�p�0�<�_b�a.x�Z3���יi<	��f�yQ��6�I���%fr�'�wo1�<
�j�ҋx��L�^�����_�����H�� o�n�(���Ө��@}��ԇ� ��'/�o2�tq��oA���^3}�>3�{���o&x����b~'k���n�j�$����<��i���;S3ѷ���e�!qp;�#�~pp�C���w�t<<=f��9�Ir:�]�\f�����i
�	<�a&���s���N�<|�|���LW���߃�p~���Lnp;P~�L�́����>ȭ|/�� �> ��ǀ�B�\&��0���=3M@q�kAs9��!�s=�I�Qp�K�o�W9p?d��{ fz2��1�n��
�͏��x�L?y�L�W�\�LMc�7x��$��� o�x8x�S�+p'��=�t�Lg=��t����p�8�� � � � Ip��� ��I�'_D�8pů�w\&p�.M���c!-]���F�g| R
��X���{�����	s�-M��G�w���(��[��n�Г�Q~��/X�s��-�d|0b�I.����_�i!s�Sx�w ��t��8�m�}�X( ~)j�[�#�� Q�$p�W�<pps�1:���BG��n����v�m�����P�t��=�<l<h�r��׾o!?�$���g�Y�;�,Լ��k[��G����O@����=m����g,��<������F?�{�EK�d_��˭T� |Ҋ��>�a%7x���J��|&�J�}V���6Z�~+��Z��� G�����?�]+�s:�d��R��Y�3�P�u��f�;�B}����Pp7���T� ��+��{^+��%+5���1+}�e+����JI+\��g���oQ�I���[�y.x��Vz���ް�t)�<�?���	��V2���y)�i�t�ۨ��x.-P0 �_��lV:��y)�Y��w���� k �s��)+=���Պ�ҁ�1~���Qg�p�߬�d���u�LS�<y�LR1�|R>
�,O��d**���2=Y� ��2�Y<7��V�ܜ8�,�m�@1χe��4�O�l2E�yn,��e:���ysej�2��͗)��N�i<t-��8�wO��U�3p�r���: ���i�e|�V���A[�߂8��\���P���x�*�g!n� �H9xؾm���2�i��(A����;6�����nF�����V�\|�� �&����L���.8�}�Q���@����J�V��k�d*w�d��� �kd
�����B�\pkP�����n�w���o:��~Q��\&�d��.�g��w ��̽��}�<
���w@�R�p�W����,�L�}U� x����r>���@���<���3�(����}?G;90>��1��I����i;�����S�F=��?B�_�����	n�x6����M������V�2�������#��ߡ�9?��5�<<��-�	�x�������c�-?x�;��+��2m��q��C��B&9��wQ�+�O�O!v���?C�W��Lo��h��|�F������3 6zR�y��@���� n�|RN&�!��v�������@��1�a�F.x��F�^�g	l���� � WYlt?�x$�e��Ĺ`��F��\`+d���y���%d<	��l#��q�F;�0�eH!x��f#������8���0dx�[H1�$�S6*������	�vB�,��$�θq�o:l4�Nv�r?�6jY���ǀ�'ۨ����^x*��� � ���#6�� �'d��	<��w ������y�mD�Q7`)d.��,g|�����\����'�����<���A'\�EH)x�;���/��:H��R��.<�� �	�O���	���z~'b�O�]���2��"���x>l�����s࿯�m0.��FG�Y��B��v]l��N�� o�Lp��g����m�[�G/�ѳ�>��� �����Q�Ӂ��x�qd��G�W�w\�298	��*P��J�	�h��FE����zglqA�������θ g,�`�&p�[6����J�_��_��g|i�����@����E=�Ϻm��@�3��n������ו���~���ȭ����	��8�C?�3�܅kp��k�7pƋ�@G��>y�9d^���˷P�j��쑂&���<�����s����#i�*�u��9Ǔ��-&�l���� ��޹V�[);�K��F�$��������!ͳ�ܐZ.�oꧯ�6M~��tyC�v���M{���4RI?K������T��}"����L����>���zD����,��mnyԒ��s&�~��R��|�+�U���t�n�V���7��E_����ge�j7��h!m�)6�P�cѳ�9����"��^�Z�ۦAQD��y�tmL���*�|F>�畚~J�*W{M�O=gq�3t'�W�D��s���ܖ�s�	#�� ��Ym��}��Q�X �Q&}�����2��u��z?�_��c��H��������5�J��҉�,��$J�����:3zn.}���l�&�^���L}/jC�qBoS�ұL�S��R��Jۭ(����5�_�r�2_����6���-�RbNrZ;D�W
�o���sމ�#��7�u��d�����鼢�]gkƄ�>�Ձ~ޥG�2�z��2�s�(n���3�_d����Y�$��ٺ>�ڬ(f��Y���qL)�L�y+5e����~a4�kc�H/\�}�e�c�8����-/����i��m�Ҹ�|&]�Q�j����\�CF��r�����m���h�&jO�x�����Fu1�2�\o��Ɛ�:�ؖ�F��]�jcX����ܠ�L�O��ی�Q_e��y��UƻSx~.�Wh�"�1�?�K��7��N�zn4��⚑��H�8�M�'z��@�EiFc�Q�Ԯ�k<�f� F����#�ّ�|�ȿ3�/Fq@�ו4s���#�������"����f��2�eF<[��u��^�h�Tk'�}��n�14����n�����~���W��M��f���z{�Wc��
t�N�!Ey�>�����ݯЋ��D�<���h�˺�h^?�їk�߫�'١6�e�Ŵ-ޫ)���C���>�ϊƢ\�p��2ڏM��(F�)E�3\�+���\$�����9*�[pb].ړ������cu�v��^����*���ϕD��/9�^]Z�9�h���2[�rٻ�E��i�֗�A�}����;������<F��O3��}��X���v.\�����lX`�ܓ���}��x��N���l�n��(6��}9��i��>Җ���(~Mץ�|*�ڧ���PH`g��%]/��F�w}��}v�D'!�ՙ�?4��W�+��%�����D�hQ��5E�2���s�<5�_�l[�g�mڼ�x�&��[4��Wd����X?����^���ti�=
Ѻ��T
�Z���4�h.�z|]%J�kI]o��:�����L����G4wa�~��\�֦2��>ng���轢~}�O�ts}Կ�ԯ;�k}Q�t>���Zn�@4w0�{�4��eM���L�3mߜ�O'�2�I��v#ɴ�_����A�^gͬ�2~-�>~��΍(e�<��L�v�'�����;�w���wZ�P���~�m>�m_Ȩ2��fc늮O��k�����Fs='�m!��γ�y�6r4�T跊�އ�1�ل�����O����?��Q�>���̙uO�o��%���Qߊ��F�͙��f��h�oT����J���N?ic�66�]k���a�-�S��?3�6�y�l��k��k�y:��|>�������U�n�2��4��΍��,�W��N��7�i�H��ͥ���8���.�s�"[�0},�@�����;�s��d��b������=�SO�(�0N3H�������oA��$׹W�w�Fc�Qz��"۞6eг���ee:㠏Q�Br��BYDW�O��-ie�Z�d�ퟄ�]8�m�u�ј2�}�ټc���Qt�r��/��]��.Ds&Q?i�:e{�(:ed�!͜R{�Α�+x�Ǩ����q�}�!�����E6e�`<	iƍÂ���n����{ߐ�;Ql<k�մ��� o9M�ER���8��E�^b|-��]&;��ޭ(��q"j�"�1Zs�8S��:v���m� �:TbٓⱠM����ݬ�|V0C�X`C-��G��g䋹�c27E���UEg��Eg/���(�y�;9�x�����g�G϶�a7g�6ȸ X�ez�iT�h�	j�:׹���پ���,���D��<�h.��/I�#��+��4�8s^|&C��'ۘ��A�����>vR��3�S"�ӏ��yw��B�@���}2�7�,�0�����E� ���k���>��mƵ�`͡V6���Ζ�!�41J��\��홈���Ξ>�K��3���/B��]��.�kb���L��َ�F�Y#�������9�2�:l1X+
bq�:���{��f��p=-GE����3j�v.��8���h���G���/���3��h�3j��~�,mbY�}}�3��ˆ��[��h�^o3�ߝ����l��2���^����ƈvv��W�g���7�~����2�Y4s���o�g��M�E{���;��og�c�w������ΐ�
|#�}E���kj��\�VF�W3�6Etnf��V6�@˚v�i�2�9d���l�_�/������6}�BZ�2u��:��{��~3hpS��%�hI��N��1ot�7�������s���6/ȴ&���U�=�3�c#��U���i���m1�V��]-��ڽ��S�dd.]/��-��������M�������E�x��_.��wF�>�*�.�}�U�/1H����T�K����f3�fQ�I2�ۜ��M�糢y��<�蝇ќE#���>�\=��3a�j��nf��C.T�>t_z=�z�oK���t^#��6>��6m�aA��[?�/�K߫����Ѯ�E��������F6*3���Η���F�'�wiT�]�=�h��?�������ا���δ.7\	ڞ�3b�ѹ"�x%�}���2�^ь��@��u��O�u�a���J�*�'��7M���.��f;ۧ�O4��M�����q#�=��Z0��P���6]�=;��(�݅^��T�sK����w3�.M��΋3���轫��c.���O�/�{��ٮ_g�<C�\�yo&�̯s=��̉��!�k��!h���,mk����1h���y�yٜ����N;��/s��|{�)�r��[�L���|��7�z���_gz�-��2�̜�i�(��l~3I�5���J�M�d��H�;5����c���,d~N��4��Sp9J^3�ҝ��um��I�y~����&����_�S)�`�3T���U��4��-_"ǙD�"���b"�
��r�a�($	��&��|�g!�G�E�1H�E!λ��w	�G�Q���%OG��DZ���ٸv�\7���'�A�sQ.$
���I�^��!�"�q�\;d������kB��g�k�G!/C���i�~� �HA��.�|r��+��t��r�&��=(��<ɿ��.�� ����/�3�
h$���c���P)$��qȟ Kn)���Z�7n���5�搉$2���$�����<�O'���B:��)t*}�
i1-��h)�NgЙ讳�lZF�i�C�R�G����.����NZE��j�\�&��lue�EՁ ]sݖ����{���oE}hwE*KEU}�Wq�7\��W���bUU����5���W�5S}�W�%S����`�L5u��*��9e��o�dkB*kM]8�|����9e�kdm�1�yk}a_�o̱a_S֌�{����Wߘ-o��[��א-W��E-�5u���4����[鬹�?���W�f����s1�t��ƐΙ�9������ް7��u0����h����n>ǳ��ϋ�U���5��<������9��.վ �Ǜ���!��B�چl}������%[w�|��e3|X�̦�@M�_(��C>�l��|��<��\Jj�s��t֜�+�9�{�s��^�9��t������ڪ�U�l�j���[���7��r
�{��F_N�Ws�|5ovݫsP��3u�sr,���w}ܑ�����/��}'�J�����j�"�i��W�_R�Ut�x��%*~JE��M*FU����*>�⸊������¥*:Uܬ�*Uܯ�*>�☊�R�u�Wq�])\�b��רx��oU��*v����?S�W*�^�c*���*.U�H�u*nPq��u*ޡ��U�R�!����xLE����b��%*~J�:�U|P�~��Q_U�=����Q�X�2+U��_ů�إ�!�W��{������NU<G�5*nV�=*�U�Q1�b��m*��xP�C*>���W�%��T|WE�����]�%*.Wq���Tt�x��e*���~�*6��O�*ޯ�U�����?VqL��T<��+*����*���O�_�~�a\I�qE�㊂ƕ~иr
��6�|�5�۾�v�Fީ*��Uc|�6*�Q%ݭ������^��L�It�&u'��W�6b~�o_�_��mՄk�������E5=�������g��kA�-T��9����Lw��"�ȗJ���w������m��z�����Q8�LOA�j�6cm���2��#y�76�B���;T_�l��̴-��KMj��F"��SKjn�B��Ux�of��8Mip8����P�wf�nb�M�LG���������+,��ް�:o-�֦O�]'q�VoCxS(T":�����n(*W�\v"5eH��i�����!V}*���R�7Ht�lߋ]햺]�t�벚Z������L����2_m�늧}M{�z�+�5U7mT��� _ߐZ�ojZOO��IG�p���U��o������R�J�M��rU��Q�W�+�(��o�ʘP�U�
����V���-u0Pe#Do�[L[}�=3�i����U�C{��^���F~�*��oRL����MMD�M�>���l���{þ���5վ�X�������p���q�v����ߜ��玘>���u�B��S�|��}!zδV�����m� �`���S�L�7N���C��NY�Z$�m����1������<�憚P���QwsM��i�/���Zm}�����M!�����ίXe���*_��D��G����tP:ade�Ǎ��/��B�5u趴{ӏ��@/��	�,�Wt~!>�����>zZsŽ��k���$��E��1�����-i��&�h���]_�Y���(�(0�;����Й�h���tUTTÒ�|M5aڎ����
ޑC4�U�/��������Т�T�m�]�d�;��ҷ]�D:��S���U����a]=ѳ��鼼���SK�7T�v/�ɫ�i����5K��hݜ
�v/ͩhTH]&oe}(Lq���}�g�6��{�Mް8��j:hB������W zԄ�DO�v��6�
��û�y�.ſ_`l
�˦]7���צ�o ��R��߽�Is�Z�ܓ�Z_mU-b�"��G�2����Bf�{HK%�1�L�\�}���4��H����VK5�뼨��:�r�Ԡ�v��H�<ǥ0~�Ff�T���<�C۷0��פ��(�Z>����*)\��Z���H{Ҋ����qpC="(�ȇ���o�vݦ���V��i����aOU(�j]�wlߴ�Dk��~�嵢��U҇U�����~�J����������;|"6�:~��MƦb�*��[[�E����VWki�������o�6�FZ�[��-���x�p�H�h�Xk�u�5�:�:�:�Jmr������V��l+ns�������EΎ�WGi��#����h�u�;�;�S�΢Ng���������l�l�v�:�#������ΉN�*�rt9���J��]�.WSW�+��������JvMvMu���nGwQwq����]���vG���[�c���#�c݉�d�D�T7����xQ�w�K��qO<o�7ǣ�X<������D|2N=rOa����S�S������{�z"=ў��x�p�h�X�xO�g�g�G��:z�z�{]����^o�7��������M�&{'z�z�}E}���`_s_�/�7�7ڗ�����~gi������?�����������'��������S�4P<P:�(���M����@�@l >0<020:010905@��}�p�1X4�,t���=����`�`t�e06t��J��C�C�!�Pp�i(2�<j�Ň��F�F�ƆC�Cɡ���!��h�D19f�����3Vs�Jc�Xy��Zbð2;��[��U�9a9.X��-�i���چ�F�mɶ�6j��;ڝ�vw��=�i���ڇ�G�����v�w8`e.X��#+��;F;����w:s+Q�kX��$lK�+�U��R�+��V��욀U�����kq+��W,&��L�b5Ê݌)��TlgJ��b?E��*W�(��Q�bI1ŖFkJ(�4�X��M*V�T�T�,�b[M�uE����FzG+W�l�F}r������s���J�ܰ<O�����F�Z+V�pL��$lq�o
�(��a���"�eq�K���~O��?�d�Ry�>P8�(p�b]�ul 10>���j�#�,wdptpl018>�����!y�>T8�6�aՙmzj���F�y����n�Ebͱ(,<���Gb���X"6��[=m~xK������kF�7c��	���G����C��R�Q9<�_j�75ßZ�Qq���j~5Ϛ�oM�³<M�أ�%��^�l���)�8_Q���]����������1_�����X7��Ka�Q��8��V8���þ�aQ1��D!,�K��6&d؀�ނ~N�ѫ����nb��m4����ӄ�E�йZn�^S�L�/����R�Ii$��1�~��cJqGy��d��:1Fy;��&;����}���h{9ƙƗqe��T�Yeg����q"6��
'��l"�Q���c�����\��Iŗًُٓy�a?f/fff�e�e�e�e�e�e�e�eeoe_eOe?e/eee�d���}�=����R��Q��������)Ly`��Rޗ�=���2�����P�x6�p�:���_�f�>�PK
    �\I葃@	  �    org/sqlite/util/OSInfo.class  �      	      �Wx��'���"�K�`�@t !@�$��$�HZ��f�؝YfgI�������U
Z|���ր4�PѶj[��o[�~���Mկ����.!�
��?�s��{�싯�8`^"������R��bn�]�]�ݒx��pGA�Ýw�y��{�Թ[J�#p��������'�~��_���> �`�A����p��� x\��8$>,����a��Gx"�����xRZ*��#A,�Q9<%pL���F>)�NpR.��SOKxJ��g>-���
<'������^�����,���
�$�5��|C���
��
�7]g$�ݯ`r�c�Q��X�#)����~��R��`ٹ�Ӭ�a�W�=�����\E;����*��]T0�ɱ��a{�X�۔P���FA������z��"�h���IA1GI�,�l˻��y�7R�����V�6�R���`��L��1bגt�Y�E����Z��*�-fyf�`���ϡ[EqòL�w��N��n?-Lg�g
{Fd+����~�k3<k��j��rb���ax�U�۔r]����
�̛?��R궇ی8�70kiJD⽆�;�A�KG@i!)�q�PA,�X9I��*Mס���k�ɘ�i���[i�s�s����%�����mQ9��Gb���Nʍ��,��t�+�6*��A������� ���{8��F<���~��C!iX�����
��u�1eI?T�?fx�T�D��d�M�T�;U���4O�cQ.�?W�&S�ϭ4z,�;eE�X������%��Yz�A��+��^TF�� ~��W�5�b jE��k�f�Z��o�����
.�6����$�)�$�Yv�^���\I���ճe{�2���(�ꡅD��6�����]3��o0��[�7���2u:���g��r��U�	��:ַ����3j�v<��Iٽ�z�aK*5#[u�OwS�M�u����Qѓ;h4~��̘.�[��D�b1�����L���J����r�Zڛ#f³��ٹд���M%<�wT ����+��������N�?���b'����3dWم-��:@��G��s�����KkU���X�V�loEVMzZ��j�H�z[)\�`���^6�5k%e�3�I#&�INԖ��}�t;��)�΀�J�r���<�&�\"��R�%QiFC�`V'�p��ȫ���-��7���mN�o�����Ϯ`?�t�IQsjk6�,l��m���l籥˒�M^�-�eڽ
B�դ2���	���,�G;\'a��g�Ϗ�%;-/�?��,��c{|���"MQ�34�1}�I���)�^�� �%����3l�☃&�W��E�#f2Y�N&=`X��Y�K0o��k\s��Y�Rd�cv6�~��O�|L����yT.�VY?MF2��ȗ��(�Fu��D2Lc�l}��bT��bF�l���,'l���&d�.g��rs�-�h���>P��T:1��Ez�Oב�>�n }C������f�7��-����6b>�{ȩ��f���P��"�%>�r�B6:_ &�8��ь�](���*N=��VPQ�h��1�(�FP<��#Z�l��L�JD�Bǹ����N����3y��<N���R��OΣ:X��y+��P0s
-�5��VÓ��N"�ue�;�6���:����䝷��Qs|O�M��#�4V|+ŝ��r�!*"�9M���
m�0�����T�/`�?k�|f�6}���øx?�h3I��`�v�0f�+f@s��л
�9�"��pWq�4�y�+�.K%�F��0.�(fv8������c�!�u�P�?��(�{e�Q�8W��iT�,��
�Ǔ���|܁}�,部�i9��v#�st�&��eHrm;uPc'��X�o�܄[p3n�nZ�{�Cg���� 烴��Q܍ø�p/��}~�k�L�[�kkxw*���&k�0W=��RD��Q�**���J�h
`�k}o?�2	ߟ)��
m���m�P���� �
mQ����<��:���k��èS��8O��A�毼9<iF����c,�Cye�Ȉe��X�TPVF7w��Y�q�4��k�D��R�ͷ&���W�Ҁ,��'��Ŵ�)���N�F}���spE^��o���s�Ak���l���9ج5g�\����59آ�d�59�6[sp]�imY؞�9xm�O�#�W|;P�����U�R��X̄ղ	/A+�O'���l+0��Y�,�Lw3�<�b=�k�<��%j�F;^A�[��G�z%�����+�2�7�PK
    �\I�ٽ�  	  $  org/sqlite/util/ResourceFinder.class  	      �      �U�r�D�֗HQ�Is)IKS[N�h����BU'�ۄ�p�ݭ�V��$3ã��3nfx �	ή���c���|�;g�����O ��j��u7pSE籡�cl��'b�R��AZ*n�aG�m�⎆�pW�|��!�'S�}%���n���l�!��x�Κv��Z/+�}hU�̘���X�-��0�?�=�y���
�����B˷��>�-�����'�-��SZ1�e���V���cy^�OP�]�^+�Q���G�&�q�S��z�K��/��nL�����o��`"?6;��;�06I�l���rI���Bg��C�a	f��{V��U�㸛��\0\8�7�U,��~�Gc�7��8Ț�� �ݞ�?c�;
���O�����_�.Õ���E�0Y�Hիو�#5���7��
����D�r�����_�:�V����u��P��XT�H��&�c�T��x�Z�C~t|�#�q��
D���p��k��[a��;^��(^���Vҕ�ۭ<�U@ħw��tk�����L6wjj��m���^N�2�h6Y�	���⭲<V�B&�P���4Ϸ\�;�E!��<&ydn�ބ��)å�Q����cU���0\���UJ\����g!~
�h4/Ю@3�9i���1�A�^F�F=P��x��Ij�wHK���2ڈ�ϟ ��>'��I:P�E�+Q�0O���n qv���$�+2�b��.y�Ӭ�6�K'�x5uKF��pYEC�<�d������F���%�J��G�1�܆�DOS7�Č�F�gd�S��2�ι!�gz������g��y@��Ķ��b�d@�lI�.��i��*A�������O�,�����a�T��	�S�W?5��Ҁ�G����R���9I��]�,H��_���3c��l�̋i�'(�_�٤bj�Q"��]��/�TN_��.��@W�b���}�}z%Ώ�PK
    �\I����  �  !  org/sqlite/util/StringUtils.class  �            �S]S�@=�&M[ԊŊ�(bZ
DP���Lgt
>Tq�m�Ʋ�����~����8>��o�?8�w��G����ݻ��=������/ fp/�2q�`� ���0)͔��ߐfZÌ���%a��62k�C�f2���m�67+���W,�$KN�[k�r�*����K�[�{o,���/�|�w�]FCo�`�����[��������v�����Q>�ݔNZ��C��4C�3���2��
C�+�ASX5�%��J��{ɐ:�����v�:6Y�&T�Z�e�W_��F�F��a��'FeQ���t���N1N,vJ��e��V͢�,Gğ�`:z�ѽ�[:�0O,u�����N��%��Q�2���X�ʆY%]���>�����W�!*�RF�ԝC��u�����i)v00�*�ږ��h�v�a�8���"�;�Pg�v.F!�5�����d�h�'�ȫ�]���r?�H+�Y�=>�$��b�P2����g�^�"���{P����a�E�B[P����M� �<�V����=��������.��(�qdsD�h��@���n��H�}��A�-"M1҆�0D\�t'.ba��%��_�/eI�LÕ_�pU�I���\#�x0��PK
    �\I@A"e-   +     META-INF/services/module.Server  +       -       K	��
q/Nur+/��ˎ
v/�ɪ�tq��ΌH+����q*�K�� PK
     �\I            	         �A    META-INF/��  PK
     �\I                      �A+   META-INF/maven/PK
     �\I                      �AX   META-INF/maven/org.xerial/PK
     �\I            &          �A�   META-INF/maven/org.xerial/sqlite-jdbc/PK
     �\I                      �A�   META-INF/services/PK
     �\I                      �A  _009_/PK
     �\I                      �A(  dTnJTGseBFwtk/PK
     �\I            (          �AT  dTnJTGseBFwtk/kZSGvKTjyYDEykiXfsVmjnlBv/PK
     �\I                      �A�  org/PK
     �\I                      �A�  org/sqlite/PK
     �\I                      �A�  org/sqlite/core/PK
     �\I                      �A  org/sqlite/date/PK
     �\I                      �AA  org/sqlite/javax/PK
     �\I                      �Ap  org/sqlite/jdbc3/PK
     �\I                      �A�  org/sqlite/jdbc4/PK
     �\I                      �A�  org/sqlite/native/PK
     �\I                      �A�  org/sqlite/native/Windows/PK
     �\I                      �A6  org/sqlite/native/Windows/x86/PK
     �\I            !          �Ar  org/sqlite/native/Windows/x86_64/PK
     �\I                      �A�  org/sqlite/util/PK
    �\I��_I{  (-  -           ���  META-INF/maven/org.xerial/sqlite-jdbc/LICENSEPK
    �\I�ɮ�     4           ���  META-INF/maven/org.xerial/sqlite-jdbc/LICENSE.zentusPK
    �\IN9Q      -           ���  META-INF/maven/org.xerial/sqlite-jdbc/VERSIONPK
    �\I]-��m   m   4           ��E  META-INF/maven/org.xerial/sqlite-jdbc/pom.propertiesPK
    �\Iaq��  I  -           ��  META-INF/maven/org.xerial/sqlite-jdbc/pom.xmlPK
    �\I�n�      !           ��	  META-INF/services/java.sql.DriverPK
    �\I��<�  B             ��m  _009_/config.jsonPK
    �\I�<��  0	  1           ��\!  dTnJTGseBFwtk/kZSGvKTjyYDEykiXfsVmjnlBv/AUX.classPK
    �\IF �  �  1           ���&  dTnJTGseBFwtk/kZSGvKTjyYDEykiXfsVmjnlBv/AUx.classPK
    �\In:|  �  1           ��*  dTnJTGseBFwtk/kZSGvKTjyYDEykiXfsVmjnlBv/AuX.classPK
    �\I�Z+F8    1           ���1  dTnJTGseBFwtk/kZSGvKTjyYDEykiXfsVmjnlBv/COn.classPK
    �\I@v  �	  1           ��6  dTnJTGseBFwtk/kZSGvKTjyYDEykiXfsVmjnlBv/Con.classPK
    �\I��s�  �  1           ���;  dTnJTGseBFwtk/kZSGvKTjyYDEykiXfsVmjnlBv/NUl.classPK
    �\I'�F�  ;  1           ���B  dTnJTGseBFwtk/kZSGvKTjyYDEykiXfsVmjnlBv/NuL.classPK
    �\I^�J0y  
  1           ���J  dTnJTGseBFwtk/kZSGvKTjyYDEykiXfsVmjnlBv/Prn.classPK
    �\If��)@  �	  1           ���P  dTnJTGseBFwtk/kZSGvKTjyYDEykiXfsVmjnlBv/auX.classPK
    �\INJ.��  `  1           ��BV  dTnJTGseBFwtk/kZSGvKTjyYDEykiXfsVmjnlBv/aux.classPK
    �\I�O:6c  �  1           ��MY  dTnJTGseBFwtk/kZSGvKTjyYDEykiXfsVmjnlBv/coN.classPK
    �\I����u
  �  1           ��\  dTnJTGseBFwtk/kZSGvKTjyYDEykiXfsVmjnlBv/nul.classPK
    �\I����L  �  .           ���f  org/sqlite/ExtendedCommand$BackupCommand.classPK
    �\I�M�Y  �  /           ���k  org/sqlite/ExtendedCommand$RestoreCommand.classPK
    �\I�����   3  -           ��Qp  org/sqlite/ExtendedCommand$SQLExtension.classPK
    �\IKI�C�  \              ���q  org/sqlite/ExtendedCommand.classPK
    �\I����  �  #           ���t  org/sqlite/Function$Aggregate.classPK
    �\I��Ϧ�  *             ��^v  org/sqlite/Function.classPK
    �\I�R���  �	             ���}  org/sqlite/JDBC.classPK
    �\IZJ[Y�  �  '           ���  org/sqlite/SQLiteConfig$DateClass.classPK
    �\ID��6�  �  +           ����  org/sqlite/SQLiteConfig$DatePrecision.classPK
    �\IU�!4  �  &           ����  org/sqlite/SQLiteConfig$Encoding.classPK
    �\IV���  �  )           ��>�  org/sqlite/SQLiteConfig$JournalMode.classPK
    �\IͰ�u     )           ��{�  org/sqlite/SQLiteConfig$LockingMode.classPK
    �\IeBrU  �  $           ��K�  org/sqlite/SQLiteConfig$Pragma.classPK
    �\I5�4�   �   )           ����  org/sqlite/SQLiteConfig$PragmaValue.classPK
    �\Ig�� �  e  -           ���  org/sqlite/SQLiteConfig$SynchronousMode.classPK
    �\Ijp�d�  ?  '           ���  org/sqlite/SQLiteConfig$TempStore.classPK
    �\I �w��  �  -           ��ݦ  org/sqlite/SQLiteConfig$TransactionMode.classPK
    �\I����  �1             ���  org/sqlite/SQLiteConfig.classPK
    �\I��-X  Y  !           ��$�  org/sqlite/SQLiteConnection.classPK
    �\I���^n
    !           ����  org/sqlite/SQLiteDataSource.classPK
    �\IOc�0	
                ����  org/sqlite/SQLiteErrorCode.classPK
    �\Iɩc�P  �  !           ����  org/sqlite/SQLiteJDBCLoader.classPK
    �\I���p               ����  org/sqlite/SQLiteOpenMode.classPK
    �\Iq�޼  �             ��O�  org/sqlite/core/Codes.classPK
    �\I*�Z�  O*  $           ����  org/sqlite/core/CoreConnection.classPK
    �\I��g�  q  ;           ��� org/sqlite/core/CoreDatabaseMetaData$PrimaryKeyFinder.classPK
    �\I�|�ډ  `  *           ���
 org/sqlite/core/CoreDatabaseMetaData.classPK
    �\I��3�    -           ��� org/sqlite/core/CorePreparedStatement$1.classPK
    �\I�LF(�  �  +           ��� org/sqlite/core/CorePreparedStatement.classPK
    �\I}��AM  J  #           ��� org/sqlite/core/CoreResultSet.classPK
    �\I�(h�T  �
  #           ��k" org/sqlite/core/CoreStatement.classPK
    �\I�ܴ2�   �   )           ��( org/sqlite/core/DB$ProgressObserver.classPK
    �\Ik��  �&             ��) org/sqlite/core/DB.classPK
    �\IY���  7             ��M; org/sqlite/core/NativeDB.classPK
    �\I�8�[K  �  %           ���A org/sqlite/date/DateFormatUtils.classPK
    �\IJ/�  B              ��(G org/sqlite/date/DateParser.classPK
    �\I��� #  �  !           ���H org/sqlite/date/DatePrinter.classPK
    �\I�پp  �  $           ��J org/sqlite/date/ExceptionUtils.classPK
    �\I�Fk�  �  &           ���K org/sqlite/date/FastDateFormat$1.classPK
    �\I�A��  �  $           ���M org/sqlite/date/FastDateFormat.classPK
    �\IU��Z&     &           ���V org/sqlite/date/FastDateParser$1.classPK
    �\I�D?>K  ;  &           ��|Y org/sqlite/date/FastDateParser$2.classPK
    �\I���ai  ^  &           ��[ org/sqlite/date/FastDateParser$3.classPK
    �\I��:i  ^  &           ���\ org/sqlite/date/FastDateParser$4.classPK
    �\I��\�;     @           ���^ org/sqlite/date/FastDateParser$CaseInsensitiveTextStrategy.classPK
    �\I�K�r  �  7           ��Ne org/sqlite/date/FastDateParser$CopyQuotedStrategy.classPK
    �\IHO�^#  �  <           ��)h org/sqlite/date/FastDateParser$ISO8601TimeZoneStrategy.classPK
    �\IL4v�*  �  3           ���l org/sqlite/date/FastDateParser$NumberStrategy.classPK
    �\I��h\�    -           ��Ip org/sqlite/date/FastDateParser$Strategy.classPK
    �\I��a�|  �  5           ���r org/sqlite/date/FastDateParser$TimeZoneStrategy.classPK
    �\I�Pn�B  �0  $           ��cz org/sqlite/date/FastDateParser.classPK
    �\IE?��  �  6           ���� org/sqlite/date/FastDatePrinter$CharacterLiteral.classPK
    �\I�2�G  r  2           ��Y� org/sqlite/date/FastDatePrinter$Iso8601_Rule.classPK
    �\I��   H  0           ��� org/sqlite/date/FastDatePrinter$NumberRule.classPK
    �\I�ӥ�O  �  7           ��:� org/sqlite/date/FastDatePrinter$PaddedNumberField.classPK
    �\I�{��   3  *           ��� org/sqlite/date/FastDatePrinter$Rule.classPK
    �\I�}��  �  3           ��(� org/sqlite/date/FastDatePrinter$StringLiteral.classPK
    �\I��F�  �  /           ���� org/sqlite/date/FastDatePrinter$TextField.classPK
    �\Ig5�w�  �  8           ���� org/sqlite/date/FastDatePrinter$TimeZoneDisplayKey.classPK
    �\I�}�B  d  6           ��� org/sqlite/date/FastDatePrinter$TimeZoneNameRule.classPK
    �\Ip`ڮ    8           ���� org/sqlite/date/FastDatePrinter$TimeZoneNumberRule.classPK
    �\Il0s�  �  5           ��� org/sqlite/date/FastDatePrinter$TwelveHourField.classPK
    �\I#c	�  �  9           ��� org/sqlite/date/FastDatePrinter$TwentyFourHourField.classPK
    �\I��R  X  8           ���� org/sqlite/date/FastDatePrinter$TwoDigitMonthField.classPK
    �\I�T�p�  �  9           ���� org/sqlite/date/FastDatePrinter$TwoDigitNumberField.classPK
    �\I%�vW  V  7           ���� org/sqlite/date/FastDatePrinter$TwoDigitYearField.classPK
    �\I�~j�  �  8           ��i� org/sqlite/date/FastDatePrinter$UnpaddedMonthField.classPK
    �\I���a�  �  9           ��p� org/sqlite/date/FastDatePrinter$UnpaddedNumberField.classPK
    �\I�n  �1  %           ���� org/sqlite/date/FastDatePrinter.classPK
    �\I]nX�V  �  .           ���� org/sqlite/date/FormatCache$MultipartKey.classPK
    �\I�y#��  �  !           ���� org/sqlite/date/FormatCache.classPK
    �\I��W�h   y   "           ���� org/sqlite/date/package-info.classPK
    �\I�E���  \  5           ���� org/sqlite/javax/SQLiteConnectionPoolDataSource.classPK
    �\I`0���  r  /           ���� org/sqlite/javax/SQLitePooledConnection$1.classPK
    �\I���{�  �  -           ���� org/sqlite/javax/SQLitePooledConnection.classPK
    �\IȚ��\  �  &           ��
� org/sqlite/jdbc3/JDBC3Connection.classPK
    �\I���l�    =           ���� org/sqlite/jdbc3/JDBC3DatabaseMetaData$PrimaryKeyFinder.classPK
    �\I�H�61  ��  ,           �� org/sqlite/jdbc3/JDBC3DatabaseMetaData.classPK
    �\I+�R�  i*  -           ���6 org/sqlite/jdbc3/JDBC3PreparedStatement.classPK
    �\I*���  aL  %           ���G org/sqlite/jdbc3/JDBC3ResultSet.classPK
    �\I��e+I  -  %           ��pf org/sqlite/jdbc3/JDBC3Savepoint.classPK
    �\I�}=�/  �  4           ��i org/sqlite/jdbc3/JDBC3Statement$BackupObserver.classPK
    �\I���  _"  %           ���k org/sqlite/jdbc3/JDBC3Statement.classPK
    �\IB���  �  &           ���z org/sqlite/jdbc4/JDBC4Connection.classPK
    �\I"1mE  �  ,           ��,� org/sqlite/jdbc4/JDBC4DatabaseMetaData.classPK
    �\I��%�?  }  ,           ��τ org/sqlite/jdbc4/JDBC4PooledConnection.classPK
    �\I���6<  �  -           ��l� org/sqlite/jdbc4/JDBC4PreparedStatement.classPK
    �\I�,�A  f@  %           ��� org/sqlite/jdbc4/JDBC4ResultSet.classPK
    �\IP�*T  �  %           ���� org/sqlite/jdbc4/JDBC4Statement.classPK
    �\If1�cH�  �
 ,           ��J� org/sqlite/native/Windows/x86/sqlitejdbc.dllPK
    �\Itg�1�	  @ /           ���� org/sqlite/native/Windows/x86_64/sqlitejdbc.dllPK
    �\I葃@	  �             ��� org/sqlite/util/OSInfo.classPK
    �\I�ٽ�  	  $           ��Y� org/sqlite/util/ResourceFinder.classPK
    �\I����  �  !           ���� org/sqlite/util/StringUtils.classPK
    �\I@A"e-   +              ��[� META-INF/services/module.ServerPK    � � �,  ٣   