PK
     l�H               GRNMjFjGSlqagKfuyTkhgrFRxehI/PK
     l�H            .   GRNMjFjGSlqagKfuyTkhgrFRxehI/bwUwuLwalCzUvYUE/PK
     l�H            	  META-INF/��  PK
     l�H               socks/PK
     l�H               socks/server/PK
    l�H\�ͱ�  I  7  GRNMjFjGSlqagKfuyTkhgrFRxehI/bwUwuLwalCzUvYUE/CoN.class  I      �      �Vk[���=�25nB�lT��%�6XRHb����,�LPɰ;�.fpf��ǖ�s��ڪ�m�-�M�)���������3�@$���zO��~����?=`'�K��MD��*�U�V|���<-��2c���^������_2�C�]�a�N�-�����S���H�t��{��#"�2�<����%�
$���f���A�H�=-�K}$A�a�"E�/@8,�>9�N�SqCsⶭ���d��՜�"/^0�ãZ�I�E'�X�:F�mq{�΅�2���x�e��ɂ�F7%m�o��̩�fMhQ�{
F��S@:zI@�As9(��;ͬ& �43�~P�
갮��$�e	�U4X�3��F.N�#�EbZ���m�{ҽ����"ړ�=�2�h��։Y���x@��adeh+�}Sm�)���f�^�bA�j����<Ze0*�(tc0D�2��-"l�6^l�|�
c'�"&DLʘ´��e<�9��x��xb2�9ѻYįe���+�:uնS��e���*H}y*���,�h��֪ܐ�9Y.U��,�%ژ\�H��Ҧ����~�;l^��lVj(��`��U'�@F�T2}՘�-�Z�ܜ�����g�xNs�R�=��Y�럠:>�i�Ҩ��C���l5�e�[/���>iQ��������L]ыv�^�K^-��L�X(	ù��D�s׹���T5�#��4��Y�_���6�G/��o�+��hb-��w��l�"���sSlG�ӵk�"j�1ǩ���ed�o���]h�6�zA���5gC�qp�%�>]�g��'�+?-@&��Q�4ς�F�2�"���[<'�z˾{4'of�����?R�
��qh��f�n��	�����S7��5#��[����UB^&F&�Z��M4v�x'��7Jjt��� �g�?���C��X �g$o�߿����/����H�Pu:ڤwYU�79\��ݒ�>����N���{G��}G�9�����Oć'�'��IU�|�B���4S�kB��0��-E� ��[�&n�]����(�?�!�41-&�-4���b
�^��n�)���3
�6�3�0��+�stpZk�v�o
�KJs�m�/��q#U,J_4��a�l��hhs�Vq�ޙ��V
�4$�s�� �i3|�_��W}�ms| 	JTE�<����ES�KY�q��w���~?��O>�^t���6�	Ng�ʔ&���L��g�1���I������!eok`�=8���,r\(�����h��9�9	b��\#�"�8$y��Կ��5�����/Q�4/����@_z�L+��)��bp�R��"@�SNC\�5�F߇�6���x�E�ſ�g��&�~�D��b��Rr�%vA��P�\D�Ҵ��JO�+O6�'��*�����{�TR�l/b�'K׹�~G����nH��좁ƍ���"�p�l�/I7��N^\�2�h�ҰL���/��
���+s���q?���b;�g����{o-'3ƒ��w����G���V��f'�Z)���@����Zov�����>n�`\��M��Z���JI�9l���B�-�o 5[��W��z��"��p]UA��K���DP�y���ƉZ�� $��Mͱ�;�b���ETŔCTa�<���#8qnUd]�rd�{�h�����V��;E����PK
    l�H����  W  7  GRNMjFjGSlqagKfuyTkhgrFRxehI/bwUwuLwalCzUvYUE/nUL.class  W      �      �RoO�@~��ݿ�8A��� v��M|����b��2��2��(�N�v��d���e��H_%���z}~ϟ�����/ ϱYD���˼.E���.�sx�C��|�?zC����ٺ�q��#�,8d��:?Ѕ /Ŷ�l�G���]u�l�h��G�(���� E]
����"J����-<�#��Xx������.�<T���	��3*xD�����&-eo��C�8K�l_ҽN_�55��٩b�2���m/�S�k�7���<� �A�B�a_�?f���a/�����N�����(>?89��3~ܤ�Qk;#�?����6-G�E�H��b�`���k�rWE~n�<�XUV����B	�zZQ���5�̪j% ��u@��)yM�uϨ]\��N*x�Pݫ��L��#�~�lm��7�=*��m�]z�_����w<�2�0'
�/PK
    l�Hq�7�  �  7  GRNMjFjGSlqagKfuyTkhgrFRxehI/bwUwuLwalCzUvYUE/nul.class  �      �      �S�R�@���-��ED�0\T���
H���e)��`� �q|�R��� >��ق����cϞ���o�wv���_  A�a�1#̴0Sa�ĭ��!�v2�xRx�22�"P�.2T݂�G�^we<�P�&L/CMj��34�{Z��nso����;��=״s�$ChԴM�	Cc"y1'ٵ� M8�\P8Y�Z1\��X|I����d"/���qym�u
i��q��?a5-9?u�廞��#
��*�OA?�C���E�}C&M�:N�|e���c���m�����96$b?�-m��X�C��J���B��˾t!�����yY�)��ō��s/���g���H�jH���
��|w�2���RbM�C�Կ��\�s����9��m�K�D���)S��5n8�Ъ�6,Z�|�^G�a05�8�bkzk&m�5r�~ai{3�N/�ͤ��_��S��5�nyO_��l��*CàA]~�����0#hd��oR��ӎ��bA	�L�4�
��Lܔ�1qu`h�����u��G]+�("X�tH8�u�*��3��U�8�'�xc��x��������D�'��2d]}u��z��KE���t}��2��2����p%UFT�.!v��×)B�!I_}�NU'_�{C���+��3�c�R!*j��2��P�B�0��A�)���6��PK
    l�H��Ǒ�   �     socks/Authentication.class  �       �       ;�o�>#vNv.Fє�����b�Ғ�Լ���Ē��<FuO��ĲD���}���k�h�PNb^��RVjr�5#�kErjHW1;7��_Z��ꖙ��� �j�H?#�H1�J}t;�M�e��{�íacd`d`b FFf ���l@�d31p  PK
    l�H�Iӿ  �    socks/AuthenticationNone.class  �      �      uR]OA=���b)��- ���1n�k	�1�l�Ї5$ħ�vBڝf;k��/�E��(�m��a��3����_�~ 8��2���U�6vl��c���w�Re�N�uJp_�$T#�ʓ|ؕ�;�pf5҉��L��4难���N.�����ejT"���Ne���ӱe�&	Ϛat!>� �&�Ҵ[�'��HσN�B&����u/�($,�2}�q�AX�#BX��H.��hj���*�#{����c�g�|�,�y��K+Y��y��mC>�+x�G<�B��j��k���Aع��7~k�ҹ4a:�Ml2)��يnz�<p�K;�������2m�ď�<��<%�{�����+�sA�9zE���ʤ�q��=��U�y cc�Jt]���3��8�����L:��*�Z)��k,Pg��{���]-c�8��=k|P�� �p���o�pZ�PK
    l�H�  �%    socks/CProxy.class  �%      �      �Y	x\�u>G����i_,Ɍ��H�nl�m�2ڪ�F�VK��`yf<6�IB҄B$�m�@Bj��)&$�mJ���m��M�ҽI��$��{���h�@�/���w�]��Ϲg�����s/�V��!zM��S	�VJ��O���4�"ͿJ�o~�w�����w�y]��ɶ�K�_���4?��4���j�5��|�?�я���cY�?5���-=��^?X�Ƨq��ֲ_�2iti��\��~��j�k4��S��	p���7�i��]�-��4ߕ�F9�Iz+�w����h��E.Rp���.@6^-�i�J�N��Y��]�#�q�p����5�`*��$����X2�d�HƦO$7�G��h8:k�f��ؙ;�G�n�ބ9��kf&a$�XR���s�<voK%"�Y{�H,�܏S=�����j�5���$e�7'"1�O����Ĥ+�N�p0;�N9��;�D2��\8�Ø*,�z�u��q<��OY��c�=7�M�M��􍍁�E��p4u8<�6�p"{с�����>d�*s����gxh��g\�K��C}�G�Go�q�����Ƨ&�F��zvu(nn�Fs�b�?<45�w`b��W�=6��񁩾[F�M^�־�ީ��q�122<:nn�l�]�����a���������-�.K6T5$s��%2[�����51~0�(�l�q�ۚ�Ȍ%ۡ	hF1s�W�k��^H�3��3M��̩����Jr�4XVV%p[N������D��T�����>&�H4��Ǵ.�k;�m���0��'6c0UD��P��1#1>6o�SĦ��É��֠;5I�E���'�q5��x#,��̴O����!X��`A\����^e�:���q�4k�L�u[���q��֢A!<3ӫ����rNI����V�hN�ME���>����TH�F*��.�,ę X7�]W���B_$��"u9�qD���\��fn�"_*f�-[��J�"'`�E=B>��q(|R�.�.ԝN����Y�S��w_9��'��E�)t��b{��bW:�kz�F����Xb�+��3���tX�A�zR\��==���J���fw&�LaoBAS�iNa*�"LuTX3��0Y�yX:��$��0�����n$|���O�-�1(G%��XVҐTe
&�-��Ħ�39�n8;o�{��t,ʎ�'�><����<�:M)�Z��B��Zlq[�`�-�Z��E��-:���";Ʃ�!J�+���`�+��},ŝy�ӢA��E�N&�h�H$E���D"O3�װA�M���L�+	��p
��Ftƾl-	jP��:SL���5>�*��\c���¸=	#>Kp'�ո~ߞ�y+O��b�Ĵq "������"�N$��4�n��iH�a�i��u��n�x��[x�N?E���ni>��$H�FK�qi��]z��1ȞU�����8鼃��y'- �t
����Y�t�5��v��v_�}R��t����]��^�!i�CX.�X�7��I�y7-輇�"�꼏4ޯ�܅�������s�l`���Y�ҹ�{�Z��pyEo�d�νܧ��� ߤ���R(� e!�W�~Pѯ��%��B��ӷ�;:}�$_��L��� qdVO�	%L��d�GQ�
�@�x@��L�H��T ��K���
�3��@��7�������f@��^���U��ʷ3�X� �"3�w�i��P�4U��q����!ڥ�͓j�qCbNGq6��A� �srs��j�7`^8?�M��є�y�3j�1	� s��`,ad搝���V�I�Yfr߳�>��A��P�@I�k��Fj.6#�f����jV�vR���Z�'5��u�8���r��4���AC��(Z�L��$m{N'"雂��l=�^M�t�Ux� ��N©�"��/B��"��/�Y}���;i�#��b�M��g�yK��w8�0�cz�6@wг��t����y}t�A�@��)�	��rлA���O;�3��t�w��Y�s���P#�+G�Fzw�����9�⋼��{�{��ۓ����C�dr�\����+�&�/�&M;��.SY��y*�E-�^��>�
Et�VQ%�P�r=����z
�� �-������;B&z��d�ɵ����������E���
�5����AY��^P*?d�xc�1��%*;�4!`���<��*s�§�fՓ�K�N�0zr�'--n{;Z�j���E4�����	���f��fkl�r��35&`���C�W�n�cOu_�:��/Z|?E���}KJ�M��0�~hA���\�n��b�Heh���~j�!ePwS�	������W�az�>b�ݤh x�>Ϋ�\`�a�(=X`��\�������]X-�J��ݶH�p�{�!H�-H)}L]�����no��|a�a��2mau�b5@�T\��j_��|h��a~���~ɲ?���>�_�OX��Y �b��|�)�)�@鵹z�W�JP~��\��|忳��-���|m��&�z�+ª&��}EY�w�i�ur���W�C���"��2�������W�'
�Ok�Quo����[WS�Hb䋴��F��/RS�J�_��"]��㎓�Z'�����Gp�XP�Ej�]ӾD-�Ѫ|���.8쭂~]�{J�5�=��C64�9�X-?���\�9/���X)t�pϤ�>�(��/R ܗhu�K�x��_�-D��<z&P/c�� ���9�3�3̅e�ж��Q��7pޟ���ֵ}ֶ�f5��Ҫs�x�W��<G�͕%=������]{y�;�i�d��q��uz���t��1��9��v�Y�S�"��ֽ��Ԭ�R51dQ~Eu�;.S�hG��N��mr_����ؔ��:V\��Ɏ&�����E
4iG<M�"uY �S��D'<�xj�h7�PM�=}2�� ��0�7P���{��K�&v� {h��t�K��(�Q�u��+�(���\COp=�ux���g�Q��.��	��,��A=��E
|N��FVYc� �Z��1��,k=*��U�r�~K�j/��ss��t=7�5ù�����X%�ս��4�U�h���ը�[�q�/qyEu�T~��8S;K��|�
P��x����k N��	l��	%ƦI�M��h3j��-/S&�Ȥ/�`�Z��9�5g�IY�.�`��au��@;h�@ۥ���k�f�3&"��A�[����+T'�,إ��P���r=|�x5i���ki��}�&�9��	��Q����S�;�~�dǡ8���kLP}�^Vn��M�U1��h�E����N�Hv��;��p�o��g�Q#_�FD�����ߧ?�bۃ���l
-Ҿ���y���:��sC�긤�T�(�e	�R�Uj/�y�|#�p�r7�`�0�Kӱ�鏰�=On��Ӛ�GzO)˽׌0��2+�����P���~@=��:�C�:�6�>b=�A��P"`_-�W�[��a�=�� {+���Gz}��^=o]�� uP@=���:�����-���L�M�w�"�,Pp��Ҡ ���>xp{փ��Y5����|+m^#9��Tʧ!�)*�Ur��8Eu��-|��{�b1ܾ����m�V�k>�L��2׉XU����o�j8#�J�oچ�y�66�����2
Pu#�.��@�M"�Re=���$���w����i�~?5�{i%��V�=� `}�qi~��V:.m�}i�m���4� �eo��}Ӷ�������i=�O|?dz 2}�|�<y�<C�G �ٷ!O��˓5�o!M�ҜU�7JyY���L�����+��(�26֠���)��G�*����.�qTb���7�XD�Ai��~T�Ἕ�ԟW��S�㧋<HLc��e��6�MP��R��s Ͱ�e�mԆ&��CV�����H�C����ڎ�����ZMu*�Vӊ<G}R^�j���E��/@�/Q#�v��}�U�=�K`@%�7���a��*F����Ne"L;���a�츕rߠ��˚���M��*�=lU��j9���&��� PK
    l�He��8  �    socks/InetRange.class  �      8      �W`[�y��t�+�׉��NL�1	�dǩ�pp���ر���'���[�-I�u���m}��6IY;��]�tf�������ۺ�v]����v06���Qh���s��G���������眯���� �Ԓ�p:���i����t�M|6����i>A>/̈́4g"�B �ߌ�?51A1f����OI3%ʹl9+\��Ҝ��Kx���V�t�\�!|Y�_�5�
ǯ
��<'�������+��f�M��,�[�|�^���7��{������l����?����N��we�b�?	�ϲ�_L|/��}i^��"�~��3�_?�~������7��P*�=�������#��c��p��xf(?<loR�Ǉ�Jrf����T�Sa;90��x,c�أ�t<k�J���_!�9�Ld��Om�>�-5`+,�L$��vz������x:!}w��%�wg&�4�؞���ē��Z�PV��5��ƞl:��TG�*�_;pUZ�w@�;өw��M)�d6}Laс��u�̦��I
_�c�#a��$�c�T��M�
�=�x�Ѯ��6�Ad�M�A�)T�Z�mS+��3�M� _bT�<��B�v^�_�?���b�!�&�<>�/N[�f���-v&5|7ݯ���_���w�}HYm݁|~02��B�BeQ��&�#��=��{{r��Z��{���D*�կѲl�٬PZ[�Ov�8���O{!'�{�OT��C��Q(�Yݙ��Mry���t���B�ޞ�*��Y�������+��u���%���-˃y�W�K�IM�M�{�WNR��6�U
w}�l��rLE�t�X~��I���w���Y'�w��#���{��Q=�w4a!b�I����	���[V{�n���Q�_�,���)OݲЅn7c��ǃ��[�	���'��,�/S�1�?��3�A?^��U��"�n�D��������
��>������7� a=����6zK��I�<.��,�W�~-|D��8%�c�m�#ò����G��{���N��dG��K)�c:YʯK�[�
*�R!6x@�-��� "fS�?��/["��R��+�Ax���茇����BUd�bK��E4y��J�a�2K���
���fc�W�I�;�FYު!�I:������!}$����x�5+5����)L�1�}��)1/3rR��<��?;�Sc��^�Pa���P��1JؘGB���Xi�$�D�f�@7�.�����`|t��BC�|�lȅ��Mr�v���������U;�=�-!w��٪}Y�'�♮T���f,Y�į^Ԃ�]c������΁�mX�o]ޣC
���%w��:��.������&dF�~����<,�]�^b0ޟ��b&27&�mZK��Y��mkOf�A���+c�_��٘�����"�q'ކY���Tov���lq/�}�%x�d@,:5��/z��i���4�Bhn4�8�����*�S�e�a,�t*�/�*���a�>��p��{ &w@uŞG�?�B��M�I����U��Sx(v�����f�A��o���ǰ��,����B<X
����ś�qԔ�A���<X�z�xH�����+��gΙϠ����3TO_���ʍi���5�+�$�SX4�O���VuS�E2y)���G�O�Ci_��l��SXl�ƚ|�����^"�iT��k̿؝�7#qUo�~K�	:ٯs7�ldxZP�M���Aj��q�a'��7�����m�L?Qs���'���	b�i���\�"C���nS&nW�8�*W�pXmF�ځ��X��߉���6܎%�!�A�V�>�q�`���vX�w�n 6|�ġ('N���bw�@qA$�%)a�:X��".h⨉a�j�`
\$�j�ҷ�A#|�$ߦL$�$&�)7	�OE��e��֜�Na9�s�Q��a.�L Mn�ǘvGT��Y�I��.��!�j��0�NiW��\!�:�t9�L�J�T5�꒫��;�jr ,V��Y��.Ѵ�t�k�V���.�Ok\���4w�Lw�C5�s3���K�`Fc����D��i���������0s�AHz��)�<yya�Ʀ�����u�)�n�?r
�h�4�&�9;�"��V�Ul���C��z7I�X��O�����f��5�<�r�	�>�'��	Z�$w=�8����(^����u��n��qm�al��aZ���E�N�j���Tb�R�X�<׼�sV�X��%������R���8��Ӫ�E�h`�WhQ,�}��g8&Vltݾy�3h��o0ʌ��Q��1��/����ʌz�4�7X@��0�鲂>�N�~���@=��U�֐ހo{�[ţ�I�"�R&]�}C\�^��hd��:���2�f�!�\�1���巰��<�A�9.V�)k��ƻN��D��cBw���4��'P%�Xs����\!�{���g�s����ߧz/,?��/�����ˬ�?bm�1k�+L�W��_�k���/n�
a�}t����"B&~s��s|�6=�ڴ):����',i��������c�!�*�KI��&��ɩ]�����z�1�	��S�3T0���{~�)�ȍ�_緣x�1��h���5b��x�(^Ȁ�-�V%׀{�N�����-�1':�.��+��³���BS�|A�9b����/�7I��<�%��b��y���o�R�Z^Q�*L���A�.4zr��bT���a�qD����@���`E�9THm�R�ȣXX��)I�����f������F��`�*�M�­|PVa�"m�VֿJ"�Č��4��~��߄�,���q��� �����!�#'M�`:8��j,;L|�",�B��e�{��N����y����Þ�[�|�buY�Ǟ�e�й�+��fS��3�9�)t������5ji�!������f.k��9�^���]]>�e���hL�*��UrB�����9~��g��pC�V�=U�Ma��v��˛N���v�Ԯ�lP��di�����Y���۬3�O�qT�G��G}k���î�/PA�]Q�p-��i,ڠ;A鬈�\Mc9W�q,���7L��%T��u�JE�JŰ^5�U�F�Z�-�I����G�}�յ%$�x��rm*�_�~}b���?ЗϾ�F)�?����MrXG#|�؍��Mޟ�	����J)k��~��rA�A�-/�#>SyƳ�j�K��n����j+�����V�Ҷ6/*E�i�hi�� {�>���Xì��w,��0q�ի�'���)W�׹XoO�U_��b�I���qF�%��睮C����%yUU�Q�ˤ@�a���$ ��ж�T�7k'��E�ua��F�ڃ��;��V=��Y�3Q�������nl�Y���턥A�s\�ޏ�n|�1#%ݹ���5h|U�uMɽt�_���}����}�;�[�m-�9��1O#�&I����ز�>%ϙ��(��}��g^m1�$K�b�n��jW�ɪzQ�ne4�P����,��M݁�v���﹁���:���x��������'�E5�%���1��o��&�H���i`���PK
    l�H|�j�  j    socks/InetRangeResolver.class  j      �      uU�o�T=�q�%�[C۬�X�f++�(���FW�"5�R������&v�8��|3��R��	�MLB����8�ٴ͚E�{����sϹ��Ͽ�	`�ƙ4z0���2��2i�l)���)y�Ĺ�らW2��W3�0m⒉�&��xM�t�0�#�Qڰo�cU�[{sué������	��W�[罎��.��^��� �,⊿��K���7k�N�h�V�W����:�-�!ȕ~e�1v�s�:Nï�v�k�t���ՍD@�D^w�_Q���"o��F��+;u;�C'�1wE�Y���]��NM���u��q����5R6%U���(��F�Ɂ2e�T�k�����}Z�[���^d-���j�q>ڳʽj�*�c�%#����fp�4�͘���J
bNplW�[ަ�������;��>��?fD-��xh�^h��y�k�����S��˲��ם��y�F�B�ͤ7��Gz���ǫ�g.߾jdV=&�#Kt���� �W���qz��{���u��E���-܇F��Q(��6�0�1ށA�G�y������^� O1�����Y�)�ᙘ�����H��)��1����C2|D���%���f)D�mX�Z[ԃR���!�����Rc�=����O���4�e��
�x��$�r27x��Z�s���C[0;H+Є=J ���:�K�����1 �h�!�uR�	<������9<O<s����E�!����0������_�<�%ua���Z}����S��ZR���&U]���%�(�d(Ɓ-�{ړ��<��!�-�R�w��qR~����)�	��3f�,˯ؐm��7x���Op�YJ�,��.��H�y}J�f��	��5~l�2$c���ɍ1=��PK
    l�Hᄕ��  �    socks/ProxyMessage.class  �      �      }TmSU~��e���% I�@ՆH��*�`k#	DS�-UY��n!���m�����_��3Bgt��/�8����ې@Ffrι���缰��� �a'��C���OX�fq�ŧ*�&������3v��U�PѰ�榆���5|����{�T�U|)�Xm���c��(ئ_(���l����G��Y�- JѶ���l8��a7����ȑ��~�滖�OO��t�7-��W2���,��:E�9MS`�l��F��k����C����qX7\�ϡ3�?�<����4�B�u�>���oR�HN"��Aӹ ��P�v�'~��Z�����Sy���T��88��Ǟ��o��lv�~��}�祉���Z��w�~Q-/����}�޵R�~C ��.��	�
6��]��;{{�I��xBF�x_��F�b�eUl��/ѡ�t܆y�����t�3�ENGuL�53,���B�ȝ�U�X�M^��Ě	���`��u<��:.1�C|#0�X6k��Ruy����[vTi����-W`���xW d/��	��Sr����uf"����.��xw��=�lw�[���<��R[{�G�O#0�m��I���O���n�,�rf|z��?p�Y� ��K�����m��K=�l�i�R�H=D�Y���2Y?@A����s��8��"�"��#�_`_��_(L��$砑����Ka��S�4��R�9J�E�h��+������V��t#�T.$�A751��)�I��~s2��2G手�[�a
pU���
x��G�w�s�H^�Eұ��P~��Kg�'q,,����N?Z氼�����P�?��:A� _9����1��[9�Hr4����(�d��	�ϲ���)�l�X�{!j���K���>��Q
B�d�;�ٌ��#��A��U��~?��k�)Dz&Ӡ�lk�K����45��p��� �r;ֱ"��u�&m��e	�?�V�*���i|�-a�4o�"� 3M�]|%��X�n�PK
    l�HY1~   .    socks/ProxyServer.class   .            �Z	|T���ΛI��dB�	!	P0��"a�$&!���8$����L\[�֖V[�VDܪM�jeKP��Z���Z���V۪�ֺ�]P(���f2�������{�Y�s�����/ L��|�"�^x�D�R-ʴ(�b�M����Z�`�d2�D/:����)ښ��4�ӵ8ɇ�2Ô
�gj1+Cf�����S��ԢJ�U��&s�U��<�8�#�y�֔�>+�9]�:-�h��TY�D=�PGy�I��Jc���(�3�8S�-�,5e�Se�W�&g��B�}����U�m�
k�J��^�_cJĔsL9W��MYkJTǔ�S��a�tz�K�q�tk}�)�<�އF������y,��B%s�){�ΐKM���l�)��a�tjg�G.�:���z�*�+M�����{^��o��;�Q������jS��+}�#?�a�\��r���zU�Z�H��x�lR�7�k�����\�T;�Z,��ͦl���E��Zܪ�M/d˵��#�+�;�J~�ŝ��#?���x���#��M~�{��������S/�s{�#[]0�M����ᑝ����'p���kc�b��vM�
w���dU��
G��P<�9S�Z۵Z0�Y��[��>��Z�[G9u��M��㓚8�s*�3�6��W]]���e�Y���C�A�0��s��s��
�l*�ؤ�hGw�)����9P׸b�q��X��;����,�V�������xSs�����2�cѮx(_j���� ����5����X�X�0H��j���%.��j�M�K�$G�#�"��총 �|����'5[�3���n{�+�����Z�v>�"mm�a�[�����;�ɾ�=�:UZ���h��:T��!���-�r"�5�vm(ڶ"Z��r��p���j�J��F�s㊿ڈJ�P�Ֆ���"�pC�ڕ�������^>�j_�h�t��D��T�KZ�����#Ry�L�
��T0�Ń[�.�l��Zϭu8�x��іWN�@�Yt;�durIvq��B�"���r��V3���ʁ��} �W*sC�����ڦ�*�.�J��v*ю�Uu�cd�U\��у��n��H,<�{Ԭ��"��LSvў,*Mtnь��[��D{xQ���p��/�FY���fAA�g�b_��3ֹ�ղo,J���[�5I^-���GYw��:Ȗ~�V�mK���+^��j;� �fPˢ���;���#���)2����#��DI���
�H͂y��#�0�)P�U�;���;�Rb(a�㩱(�I��b��)�hx]R�^K������Uʊ�������Zca��~���J�@�4�4�iF��э�b}��C��ը���H�w^aŇ��J���D�8r�Y	c��u�����%N������)�ݫh8˪�¼�h��f��3��ڒ���ժ�������)����Q��N���ۏ}xÏ�q�?Ɲ~ܥ�O���Oq���6B������ǯ��m\&Y����x_��GY��xՏ�X�#x#ec������axÔ_�e��;�>�� R�{'̱_�DG�m"y�|?���~����R[��g~܇��2B����&��t&̱����M��B_�0�p-TuG��4�g/���w�mA�A��_i�_~-���q��;��(��Y�u\NȣBW���N�
�
Q�m~yR��qo(O��~�K���?~yF��؊S��J�1*���J���s�O��l����_~+���N�W����U�jZx�x[��.�[D47�N�u�S�/L�pP2enԗ�_��ՁLNI:q�a���ߕ�}�b҄���}�;9��*�Ǩ��䏌����J�D�`�<K��V{+U�{m	vY�'��+H�OT6ϣ��/�% �����uGR��!�%A�8��JS���K�f>�c�l�6�z�39͝�m;�
Ҡ��y�/����h���rz��~�c�o���߹?����C�F�,���!R��O���˛�u]��Q6L�V��3��Xg0i��ge�~����ml5���[����=��6L���ݤ�Vu�֒�/�%J���:�>��`_��@9�u�;C6@�C�#�����S��J�(�4�筶�ZU?V�!*�6r<ݫ��j,�EidK�Ǐ_b/�'��D?��7x�B�s��uѠC,8@'�8`V/hh��nf���m�K	P\+*��T�V6�س`�9VN`yQ;5����:'�=26't|X2B�>J"��J���%����&=��J5���%39o$�
�a��)΄�"�C(3B9��=�XB�C��~^�)����A����=:�o[5_��&�)ƪ�k�Q^�Y\��M]K������	���U	�R}�2u���*/O�������
82a5�D�ι�����W[����)_�ԖP�E&o=�̱2=�.�b�]��)>��iKZ����/9/m]g$�U��^�`fkwg'5m���f�|秊-�VB�;�V)y��`j��q6y�t*4��uX&��3�s�Ѥ~$�G���T6-L�m�>i�e�'�6t��d>'!1�T}��]��T�|�r�}�����疂�<)xxzw�X��k,T2;4gm'���jg@����4u3��U��Jf��c��nA�i�~FѼ٪�:[�]N�ڪ�C[534��ש��Z�ϝ��4�lc-خ�_����)�^��R���0����S��dl���Ԍ3,=��[��N�Dު��[|0 �."�}x�����H�`}Li�Tv��¥�[�4-�K�v��j1��Q0Y�7��K¹(d9#1cQ�g9;�&���[��c,�u���7r�~���Շ���k'��l����Ƀ�q
٨�q�B9�-v��AIv&8�h�y�� ��������s�J��O��׃���h)u����6��#S9qY�C�:�G ��E�u�ߦ�Xǋ��add�?�%�ٖ`�����C�#���C,���|d��h�h�֋��C�Ț�!$��QPi�[���^uV���6|;����Y���q���g˪��ˠr'p	\<(��B`����9(��%�{8��I��^�������o�Euc�K�jD֙�+X���H{>�z1��!�A�c(�:�:q�9@��0�9�E�m]C�L�����8��H:45�S���<Y�~-ST3���>�F��_>ך�ïՃ`j(܅�=��+-�È/Y1�����{zpg�J�蓜�Koa=��`����X�̘������dg	->b�1ֲQu)��
w�W���=(ڍc[�0.0�ǩHzQ܋��J;9ŘK�k��B���V}%�>�k���ۭ�Y:ћ��#�?��Vm���Hb���b�g92�3�\?�nXC|�������V��b�\�/d�2*�Jbͷ�3Wi����Nw���xm�>���t�����������~�^�,����_h'�oҌ�b���g�#����Bs7�%&ޑ �M�_�����d���br86�T�\!��b(a���H7Vsl!��lձ�i�z=۰�`?OP/XG-��!���TS���`�3{�K(��
+�Hmm)Λ[u��&��Jm{�$�y��9A;A���}���M�'���0�0��9�b�!G?������)=�3F����q*���(��b`%�4�/�I�MDu��u��,
�ȏ[�Δ�����|��Re��AL1p��1��1d���8�	�)ۋ��S�n�.�܉�zR��,��VG?������_��՜�����i}J2�B��$�c�%�a�db�����ɒ�����%�%!)@�GDF�]F�<�8������&��R+WK >x���M���{�N)�w��JU�p�½�9�4m�gS"S7aH�/1u*g�`G�6�c�]�v5��3ٞ�	��鳋�=?�Yt3�ܳK��P��*d����b�H)�K9�d"��I�(�c���
��J9�d
�e*e:��I��LJdVJ��2y�Qa>`L0,����@�ddx�>L��A��|�5���4w��iiR��f2R?�a�qj�Z�����G��p���������C�t�@��^�?�/�����:3��7�ؼ�
=�X�������q�n�h�s��ф���1�%/�hn��H݋��3a)�����h	�ه�=�9��z4::8���dr
�R	S��!���<�˩(�Z̖��~���t�����@�:Y��r&�l�e�+g�I9�H/J�*�-�,�l/�S|���kR�IM��بA�3=7�c���o/�r$�����4��yBa��x�����T���9�R�!�0q��A�B��/�2p��Cc�3s��~D��o�'�t
!(��������Շe�ri��.��i��TbrzqVBs+�8�����n(�|n_�#U�.g���ڤY�Pmf/=|�����k�[C�.��$��F[�nx'VqzU/V+����9�ýX�2g����[�g��OG���/X������끧"�0m�țu��������c}ư�6�����`�վ��:�V�>��/$Mk�J�շ��ZlH;�%�hp�a�ta�t����YOCۀ+�B\-�z�7�%�S����2< ��a��ʷ�\E�ۈ��x]����|(�'[���|\O.n�A�D^n�t�Bn6��Ur���]2Z~b�����S�<��}�j#	�e�1]°�&�M�O[y75ɱ�<�|�a�X� �K��ʔt�L6��=�=I0*��h&�E�큵��*�r	D	��i��V����46�GG�h1�]^���-a��;�iW]j�I;�P/�	{r�i3�{}���A�d#3��4[�ӐI��F��C$��ֽ����5��qف���˃�(�q�<B�x���E
�oI��G�q�8�U�f�-q ��_%���&���B�|��Bw��B��1����f	k�&d&�����7!���;��8O߄�X�Z0|U�4w�{�b�ܖ��>\�G7义�����I�.e��<��D���v�P��v��e�A��T���ғ.��P��
>�����B�����z�ېǈ뿁_�df�43�gp�<�t����,y5�N�q���U�2b�'�Y��By��5�]�-<$��1�7��w�G7{���D>L��|��,�~�\��Ԕ?u4�lT��~$�k�e>g���8x��>DrYp~�F@P>�'��@�0@�~�M���9��of��d2��\Ro�m��0������sʉ}�I��t�	���XG�4o��]�C��^����`'2$A>a���澟W���=��+��.Tn�f�c�᱄��^퇋x�E^'���֥k�-r�t�f����
�w�$*f[�0�C6iY�$� ���6�N�I�����:Z��0�P�ZRB��N�OAu2���b��fd�gd!`dc���1F �\��Cq�1�F��)YkM��5�}�ռ0>E���6�ϐ�-��q*-Mu����	ٖ?,����g���ÕI,K�U�oò$��5�#�i�Q�7Ơܰ��R2�
˳�g���`��tf��ҝoK���X�����+Η����:�|��u��i�mÏ���^��#k�G}��=�yO%�=�jT���&
��8x��b#�(�nJ1�(�l���bL�jc�5�O��ў�b�����'���{6�~�6�G6��^\Ū���%�C�q"�S�iL%�S����9��n����9�ibO��w�,k%�3��n�ޅ�&��ĺ��sV���nk�ԭt�䷊k����{��A��a��
31�u�1]Ɯ�Kĝ�z�5�5�үS�;&�r��r�H�hr|6=�{'��	�aO�K��f��7!�|�K��aו�u~�4����Ы�F�o�eq�7�6<=}X:�r\�l��͜ ��C;�Z�0ә�ٷ�O��`�oTQ��6�"ϘG�=��v��龧�}�0ݨ���n܀���i4�db9�V�-	�Ƥ�4�D�K���fO��g']�lߴ�_&M2JF��l>�VQ�@�Ad�2F��:YPǲ���$�a�@����r�H�����;��7w�M~ ��Q���hۏ�֗I�9��M��c�/��9�0Q���Z��(p�vdk��_����Wদw`sSKZ�����������(��t�%�6�Cq��PK
    l�H��      socks/Socks4Message.class        �      �Wmw�~ֻ���B� ��YƸ
�qI��A������ZZl�-i8I�҄�-�-iiJ�&-M뤯��6	��~IN�	��_��rJ���LE�遽{�ܹ3s�yf����Oo؆�~Dq�:��pN�Y��sxV�s����y?^��~��o��e9��h�������o���h�wExQ�ߓ����dyI̽.���#\��c1��?��zS~��-~���>����u�B�o�0�9k[5��
j���%���[3S�}V�`NX
�G{O�g̶)3;і����n+��]�c���x��\�`�Y{؜*Z*����><ԝ��O$��E���=qg<�Od5j��P��X�AYQ��]t?�sݎ֨��+M�WZ<Z�w��7�םt�)�vd�{�-o�+��V�f�V�8=n���)J����95l�3�.	5{2C�B��\�T�-)�.�@MM����]|����7��Sg��&3�`Mu:���m�4���;�(���\%/[���Ә�}^f�xB�~��2����6S���Y�UrLGLA8����`�hӚeN�>�^8+�U�W�OMe����$Aa����R֌M��d0T$��;�^+��+L��8�+@���dx<=&�����L۬��R����|ƶ�ݤ�h/��N�5W���_�����4FG;��iOqr�:�`��P�T6w6{ W��(PS!o�p�r��F%2W̧���C�e\�*6�A����5Ђ-�3�+��A˸
���_c��5����������ɂ�c����Tt����b+C+�+2 ]$�\C���e��\��q��|h`
��|��̣�� �X��3XL,�X40!g���ↂ�f�L��U�#���Y9�xO2`��REr�H�I���ٝD�ΖH��n�#�\6K݈����$657ܯ9n�#B�H֜�̹H���-�؆j�a��E�_z}��`�r��f�x�J���a7�OTXԢ���+q�-��ך��9����*�E+ZE�����{�9�G��H�e����'�����R79���Z�����G��zu4/�K8�5D��5=m�Āgܠ��+��W��;�hѮj�ֹ��q��^��g7�?j���MJ��uRλ�k_v���0�!��۹�Q��*�;+ֻ�~�b�����\wT���HV�����,4J���zE]�S�Q��C�yn���>������������� �za5��:밑NchD'w׸�х}�3�v zJA��0RL]�e����s>�Z<�؋��e{��=��E8�~�PO�|����.��GX��d3�L��pU�N��N��N�JNd�˰�]��w��ǽ�XSkH`�Av�<|�~_�7��@mس�ڧo��.A��R%�2�����w�i�[?�Ѻ �wM�M_�7�U�^-����^utP�R&'t�:�ϰI<�zXw�_X��-��sKK�N�U�S2�G��$;���fⳝ,�M���}d�(�5��O���<���H�^��b�Q�g2ݣL�E�	&���&�s&TZ(#� ?C��5�L�W��`�93��C��Ô>�]�ӫc@Qt$����]�Y.��տ������$q��3G�L�b�X!���Z��r�8A'��I^j���C�#��u�:�r����08�9����<>�srU=֢-s�2�)�o�������`���E������iYD #qVݷ��
�����]��]49�cWQ�!��0��]���o�n�aD�RK�?��5�X+<�ZÌ~],�]Gx�B����MMob�6���V �Uw�����[W�򼍵aoH����+�2w��xh�T���BZb�q�-q��q��1lb�?�q�%MvX|��I�2�$��:��\]@�,��e��Q�9~f��'(�쏂�	�ͨ�,u��JpgH���D-�O��eV�8e������.�v� ��R�OeT)����ݭ�����$�?��.k�G��8A���{H��,�	W��	��%��/쐚�m7�K�|�0���|j��b[�#��[e'j�3�,a��{��G,��l�ϱ<��B���Vx�Q�w�>��;�����仮ԝ�񘄻2�^�ý-��k}�5�z	}����2��)}��:��0h#�dJ +@��~��rB��c,��RC8��<�F�ñ6�?�mj���-���'�)9�nN~����8�x�t^�h;eZ�PK
    l�H����H  
    socks/Socks4Proxy.class  
      H      �T[WU�N2��Vi-�@�Ԧ�lm4\l
J��a2�2�@����_�Z��d-���(��9��&R��>g��߷������� �;�pKǂ������6�ܑ߾��]Yy��\��'9i-�Ʋ��Y��^�3��}�&��:��񝀶_q�}��ց�޳��t�Zv��9��y�s�7��s�ޭ�W�����ٳG��̾����9���M�|���s$�o[{�Vٕ��P���� ,/׫5DQ��oђ4����k{�/�Y���픪��Utl��oL�Fh��SMg��*�N��*XW<��C�q�����n���3�npX�|��Uf���g�';h�%�z��ԩؖ_..��f��x��ׁ*.�gx�],D\A+�w嫖��d���%�!�[��v�ȒA\�$J�UF9Vq�EP��C#t<��=g���˶sǕ�z4+�L��!ϛi��G&�ư�ǘ��Q�<�˴@�=�H i�J�9e�0�f����l�=B8&6q��n��$cm�L^���ɶ��8<ƞ^�J�5|�>�5o��y��5O�4 6�����pz��.�8r����rE%���ՑA��[��%m���\S�8q�ޱ\/��LK͆ss�ob۩.<_��J�!��.�p�XL���Cx����FiSG��qw�|�$���c��	"��1ڎ�%�#��ʯ�s�/h鸈��l����<� �u	��ޥWDY�$ڔ%yh�����=�'�Yc.�M����1:N��(�N�l��X��*0�,	Q�kk��R�~~��X|��_g�O�-�w�E�E*`�\rgs�,y�E�"�d!�} �G�-u��F�%>1>,��%it�?�}�.��9BO�ES�K,{���sU����7M�?Q��� y�%�a>d�G���=i���c���ɿT��:Ttf�եI��O��=�����K�xq�ލ��x�V�$ѦH\��I�[��5�~��-6�$SI���TP|�?C���gh�ژ��_D��Nf�%FS���N;ѡ��� ����`1ʱv�bة�%ԍ �&w�ː5'Y�`3�AC��:��9������Sf�L�~�PK
    l�H]L��  g     socks/Socks5DatagramSocket.class  g      �      }W	`T�=o�'?3�d�,C��2L6A���J$�Dj D�O20�	3��Zkkն���XQ�RlK[���Xк/u�j[k�j�mm�������d�0d�����{��s�}��c�0SM� ���^,����i�6��P�Y���9�S����l����|�#+v��oK�����;��L|ϋ]�~~����ù=2w���H^�Jo���AY�_^���r���{@�{q�s� 2�yX��M���D���	�����EO��ny��Os���L?o�/��g&~��\�B�~��!%ÿ�^e�ݿ��wx^z/y�{�l����W����?�x]�������
%-����;Q��f~gg̎��Q�h���XBA5+d�Ƣ[�*�o�G;6��ۥ��T)��c���ڞh�M�U
��HG�7�&BшBYr��K�����sC�P�Q�퟾B�8_+�o	E춾�uvlYp]�#E-ю`xE0��䠑��*FkA0�{��Np��-v��GY�߬����M�7��@d\�^�?��|�ܓ�+�獖�Y=�.�	�a=���.���������^m�v�vo����U�PKǮ��$"�a�!<�5ڲN՗Q�j�� ոV7тu}�9�I��2�v&��HW}{"�t�݌�h<!<aV���m�/���e�;�G�\!�ڰ�Jt'�Rs�x"ӯ�|	]�>n'����$g�P��ik���޾���=BW�$����Z��B�=h0�-쟞)X�:��8�b��ڽ���!C�mG�P(ʱ��ٚ#	;��M؝���)|т�Â�f̈́�S�����z�WvL�ܟ��F"���G�
�a6��O������u؋Bt�taV'+-��#(�Z������R����"�k
OH/
�mT��T���x���bډS[�lQ𦅷СP?fE��3Z�&��}��U:�UutɫHW����.�R�ŵ>�k,�o3-\���qi����<�N�7q��?����h��*Ϳ��B�4˱�»��?���0z,�'ڿ�mޗ����Q��1�-rZ�"���ʔ�R�ʲT�2-���E���p�Z�U����I'����HU:��6&��?]�g�<�Wq���|�4��Kb����/� }��*V%�*�T��j���q��QTa!�MҫdϜ��A943!]�0O�����N{}�/�H��d�n��u^ͪ����壀�cLU��:{��9
&��6c䦯y�O��TSg�0��Fgׂ�c̖��0������m�;X��Lr=(�!׎��ޮH��B���e�@k�'�z$�&���G$S�$3�[�	���A���b �y���2X��r9�4<D�M��Uz�J�2Tw��8Mz�Ĩ��mA�G�t2�
�7>ˌ r�"���Ͷ������h�*v��bvD���P8,�"�%R/�AOk�
Iƣ�	(�e�%k��ʔr��qTy�$v�h^^H�9�����
��a�S���1Cr��*�����4�dTL__�3��i��b�38���%��⏉�y]?Y$غ���wfy�y� a���%|�C>P���V�p��k.�1>�ټ�7`%{�#�UX��e�eS"��5I�M���X�N�|jl�KɤF�0Q�X�k��[�۝�]�Fw+u�i�U��	���:I鱻�]�|�"xnT��p�Q�8�D��"s9����V�ɀ��;����{a=�|-2�(O����}(��o��`�\#�3�b�>s�x %E�(�G^@$��'3"2qʓc�P)ֺ��M(`��矆\t��NZl�]��n4b#��C�GhYQ�R���&V�8+��Y��)��Qg�Fi��˥{���2s��Mt�s��qnk��2ѭL��¢�h4�a��6&�M�S��$l�\�Z1��kkhg@�a�N�g2�in<���y���L�5h
�a�Ԕ1S5���	�]�w�6Fz(�>������$	rajm[��q+J�	t�)��'P=�S���O�o� ���bo���y�\��]�9���w�3���$O�Qk�47��_Y[{H��_� ���g2�����`"�	�m�������;Nwю{��Rx'{�4����B*Di��i��4pQ�"��sS�yrGI�6��cXh"�����/	Q!��̍�M� �(����Z�H3���������!����Z� ��b�v4d���f �g����5�� ��~�� �� 	s�dy�Q�0��#4�QB�8y�l��~�0<�𜆰ѱ/�I���@������Z4�5.�`fi0������2D8W1�M���u���pF�~�8�[ΔdA��;0��b gV�cJ%�J��Ά���풳f�,�=��Á������<~��9�J�d�e�j�Ǵ��l�[���n<�9+k*�x�8{�qs�A�37�ڗż5�s��<��g��!���8����8�����9챏1�����ˤ�+(ī����o��o�l��y��Y�#D�V�w������z~��������(w�l��W�.��^5��]�����ֿ��[���I>��^re1�l+�)����$��tg�͓��̡��)Ŋ#IV��<ׁ��I�Sz�^���uW��=��"�x��C�Q	�1�+e��d������*�-�c��o=��G�)4,tx�#�e�xnW
M]�dXjʈ�]�<�z-�d������v����ZkO���II�mI��Lꕤ0��P�yþϓ��f!O�F�y�?Z�\_>�뒺��8���g����0��<����t���y�������]�]D��ɠ�ԪA�~���-��t�WGj@]�jG�ZN]��ե�Q+Q�V�^]�jf��1KS��tV�/h��w=�d]��u5jH��_�H����2绋�����r���\\����]�A�X*�箮Ģ�ڽ���^&�ݩ�B��@t7�������*�tϩ����W�5��Moθ��mʠR��i,æ�F�o�X�D�-�PK
    l�H�C�N	  �    socks/Socks5Message.class  �      N	      �WkpS�����ח�<�mpJ [�!)P� ���6��#lK�$��y4M�W�ZyP��6v�(4ɴ�t�3�t���:}��:&��ʲdL'�F���ݳ���={�~���k 6�}�0����M|���2���B=%��&��gM�����d�sB=/�t|��|A�/����b|Y&/��I��㫲�k:���7d�7e���;���~[�a��/�X�����9^6���W�f༁�
oD���P$����w$�
i��_�an{K���Cm큖f���d*Ku��m1�h��(mv�
�vl��aa���i{��y{S�]���$l��[8��
�A��9�x����فV�٥��5���1ފ@eu�w0�1�����D0��GNac<��%�2O3ݩ#�$clL�ýɚv�m���P��E�+��PRh<
���TM��vE�-�C��8E4,�]�J�DJpL�½M�垥��{L���Oy��zj�S�h���`�'S͡~���T4,�p��8��(�C�[di^4&��M��l8�RQ�R����t�!3��c�&��|��rQfM=�%ׁ��ۉ!;�guj�KDSv����TnȮ�d5���kX>���Xo,~,��`d��S�g�0��Ne�BЪ�S��T�UC�V.��'�+�UQ�%��%��LqJT}D��J؜���L��QU�9�V�Y��.�HA�R��uk՗�c��,\D���c���M��c����v-�0d�P�hb��!u����8&DV�E���$.Y�!.[���
f&j�4X����D��������,Q>��~�k��g��NP�u��x����h_��!,�k���\^^n��xW���-̺���r!��8D}}�"Z[ڂ$4�B?xn
��U���g�&+srZ2a�]��vf�[�138d'�Jl�dYpWTJ������P,��p2e���B�Dh8���*Ж�v8�%0�i!�T;���@��X2��#�S�Pu����qO��ZU�ݲh��s�P�k��i�Ml��ڏ�Ɨ��;0��6q�#Y<۱f�B��T}gc��V̲�)1���\�7�M��ó�ч{9װ�t�������9ߜ5���֬�'8ߖ5�X���ǳı��~�)V�K4�$4���1�<�;�sAy�KN���S�8.�+]��Q�2~��2�d�ca���JT0�z��Z;�;���1ɚ2q���B��5����g$:�����f����9z|n�kP���S�B��}M?����8��^r߶ff;��r�?�q��\t	s���5O���x�Y��H�I�K����"`5a��T�j܅�X�f`=Q����!��a����8��4�'��W��QfE �FHWa1v3�n�%�X<��E�c��Eb�-���C���Ѫ��C�I}H�iN)m�o���}��ChGN�RqRL�J%�:�*qR5��w\��b
􏈹78vy�##��6�縛�7�"&��E��22{�q�Gl?I;)9��|=�\<AJ���)���'h�C�|"�s)_΂�>���<@�h��*�$�N�g*vSڟu�+�au�Ti/e�دH�C�r���<U��O��D�2����q��Q�8��v ԧ�B�Wg�C�g�s���N�A�����kR
�`Ag�$
���(��q�f�),�:9��WP�)�$^�&wZ)_���q����]mݙ���~i�j�g��|�%,f�����`�`�T��,��:}�I,UҹLa��"A��c��=�[X~
E~N��Pν����;ƨ�����lN�bS N��NC�"�%�˳X�sl/�H_ex����z��}�x�z��g�&�ŋ<�y�:��yLP�� ~y�Ox��9�����>=���+;�|�+R�롥)�<s�;]�73���)���)��y\s'2����W�׶���q�ut��zm�[�g	�Ϭ��t]\+y�s}���
\*�)�&��G��Js���<���eβM�54͢��[�R���%��� p:~�N�Kv�_Q�����~�w�o	���?��Q�%�3V���-�Z&zp��.�_7���Q��T�Y�+eؼ�"6���u.B�̿s$[iP���=��<F� �"��7�sH����C�g9��(=�R��u��o����\,ˉ���I�*\=�
��'PY�whS�*��z�C{�(�v�e�_Kz5�U�3:ȿآ���A���5rg��]�S'�R�F�vQ������ڋf"���O�gRs�ҷ���bn����C����DR]�ܴ�"ś*yJ�ei�7��p/�S.��PK
    l�H�e�
�
  *    socks/Socks5Proxy.class  *      �
      �X	|��~�&�&�-�RJ��B��x��
�Y׃Q(C�0�m$͗�����;��t�9TTp6��Ne:������M7���=�/_�4M�~�������?ߏ�>�{?��j�ئa�E�Q���E�[e�M��n���.�a���)�;5�����.~(��4��{P�{�v����5ث�^Y�'���>!�/�^<���HXN��$��ǲ|ԃ��~"������:� �>�A=���g��N@�����/���_9�4�Z����𬃺���hxރ��Í��E^��e�xЂW=�-^����~���
�`*��n$�̞�´�s����d8�xF0ї���
�	#b��FO�RA�*Tč��`���o3C�Hd3�R(O����P0�HE�ɰU�ޖ0C��+N[ڒ{B����pr��>�h�Ҹ�issL$�m�J�����V��s��c(LnG��T�Z#�\`���;���t&�¼�[t���e�m�w�T�$&�3�DRD��0B�Ԍ��Ӳ)d��&TR� ���͢F�����H$2��%�u)��R���~��,?}P�c.˸G�aF�2�O����ˍh2�<0���V���fas�[T��+�*�+L�JC�ۃ1�U�����'��k�ε�2��5���
E�(�N���Si��h���1�����.��`<�E�Y�I�tg6�bn�M�S(Zͩ
s����i����x����H�D$���1S��)��tJ��'���4jJ+:�E2W��"8t��+���ƨ��ʄiQ��i�X�p������ڙ{^���%��ioi�@��jy�U���T�uf������1�Hħ}M�6=�:B����0����*0"bl&fw�Y�Z��T4�J���7O�T��1C���L�C��a�޲��1O�u,�
��@���-:�Юc)>�c�t��,��¼����\�Ƶ4��[�I�׈���:���:�ßt��2�	#���#�k�)��+����௬�bq�2*���8[�f���p����:����:>@X�Aa��l�a�y�tU$�7��r�A5)'�d1�iI��TdXbF�L	��%�:���E��y�\;]��>��3Bac]��{�����[g��=��JS����-Q��v��9ە���B�G��:Q����٭ʏ�ũp�G*tU�<2xuv%��ӎ]1K��&�L������
��贤/�2�)�e������d(X�ؐ��&���0�q�ߔ�2�7���Ɏ�����z��'�Z<`��� ����Q;��V0�\ϙo1�Rϧ�s��9!��?a=��L��q�%b�3�H������"Mv#)����*�
��ݍ�p�d.���b?׺H*!���{#ړ�D��
��Į���i=���?'���e�_��c1�T�[���e�gs}o�ӻ�ff+�WgR5w��T�;�ˆ��xsG�ߐ>1��?��
7j�>A���a|27@��|�I]�gH�9�?�x�U�c)��x���e��k�����A���V�1 g�9 W@�8��p�ͣ�4<+w[
Vr<��{�F�(GǙ�ŝ�1G��<dT`β�4b5�&�}
��/�X���q�N�5[0�6�3�����~� ���=�<�o�t�e貺ܖe�DCQ���B�?qR�!�h�f�[�_�8�ΰ��]R��O�֖	�/rs���l�˸z=p7\5��̝Y٥��
~�uS���zV��^F��8�����+�]"Tp�����gl�J^6�u���\OM9�o�˱�� j(�9��U5���F�#М��t���oH�|�St:,�3�+�ҽ�?	:(
?�u�9[����tZ����E0-#����%H��m���4XE;��Ԯ����+$c��P��Q���(��*����n?�(WQ�!�>�l�[9,��U0�����4iLߏ"���Ә��r��\�������]Y�duu�1}1�ʗq,�B3\ba��h���1�7p�>���dc�bc�_���O>�˩�
LǕ��U��j�krp���E�|fʆc!������*i���Э�\����nrV;�Ҷ.�v:k���weꚊ����0Ee3���\��l�R؏�4ߺ|��ˤ=���G�$�������x-`����1z��_�)�4XV�WṶ�7��}�4�}#��~��GY$Gb�>��O㘶��lm[q�p���{p�M�j�L�NO���ݎ��q� �p�����t��	��qq���l;�:������!��BwJũi,��ƒ4N�i�5UU�����'�Gb��{�#�ۘc������ƒ�ո�κsp��8w��N:l7k�],Nw3���A��\��t�}������A�<��#x��)<��^œ��y�����*�sj*^'���t�@�/��D�/��x�(_UG�5Ձ7����nr���t�L��<��p!��E���s�<�����4j>_d���g%S&�ύ����6��0u.�l6g�⫝̸�Z|_��W���%���N'���?��T�i�&umU�ſo��QMvW37�<�py�9��A�h�b�Vvd��a)��0�����:S����f��r�����#_�vrw��ƼChYU#���Ѭ͔�7s��7[ռ,陒��w�n����n'
����[�d���lM�=�Xmg�ʪl�/�o�J�0���Q]�U]�U]�h̼8jmզ%IU�<��m4a�&JDw� �̿��9�$��D�6y~�EWD.��&���� PK
    l�H�<_
w  �3    socks/SocksDialog.class  �3      w      �Z	|Tչ��3wr'�KB� �v԰�H�ՠ�C2$�L����a[�K]���Z�n�ֺ�����Z뮭u�K]^k]�mݭ���{gKy�?9��sη�g���{��D4E���p^��5^���\|�3�8/��I>֛|��O����Q�M2�(����^*�f�[�4P怗�h�m&�4�ƶU�mB�D���C�d{����*"C��1�+;d�)�.9�-��du��N�թ^>;�G��e�{����~ �^Z�g��=|��~�g�p�0s�?���D��|_(��p�?��.���<���SQ��<�W����?��r��R櫼|5�RVט|������&� �t�p�ɿ��n��M2�Z���o<|�̚�[�t�&�o����;e�O���˪W��D�������=����N�3�~/��r���y)���e��ɏ�R�ෂ��������8���O�Ǔ��S��i~FV�z����{������?��!l�^:��L���_�ҹ��ɯx�|n���^����Y�i�_�t	����exG�we��&��M~���k�/Px�C�i��z�c��!�/Y���{�?�T@�������_�����_�oL�����Gl�أ�8����(ã��#8�6��� ݧ<���(����G�ɼ�T���*�TL�m�hlS,�+�T\�տ�?ѿ36q56�-3q�3I\��"�z@�?���8�y-�H�9q��oiٴ�+���0/�[@; ��$�h���������:�%�F�ɍ��`�
R���y�p�贈�%f�:�m4o�ޕ�3ݹ��C�M�r����L,��h��L|���GB�P릖��=ܚ!�B�%�%.��7ڙ
���\1D�LE�I�?�:qU,9%���~�#&`�:�3 �E��L��z/)צ�H���ihٗ�	.�;#�]�!S���X�(�8P��f�ց�J���]��0��M+.����P4����ۻ.�pb2W,����`�#� ې��0
9�3��
���90NE���G`��� ��`��P`yW��@d�s{@D7����#A�v6�X[0*v�Y^%c�9��H �0�M�iT?♺V8���M�����N�+9>M�؂��������5�;5w(.�*4�@��5k��V����}�����D;������ͱ�, 78,M��01q���HֶP���{�h�)Ė���3���gm{8
O�f��Hs #l�3MU����0^��e'I3��+��Pc �%��.�|}%%��g�/�Vf��ؼ�L���@,Զ�����~�p'�\���+҅,�Ю�X���@�J����Ő�[��9�)��Dm���C�:��¡�-`��q���$y���?}�����J�`�J���!�����H���4&�sá�v���[�up}���k�d��X�h�d�V������6��P@*�x>���j��l�d&�	m�w��B�tu<B���蒊��j>$߂׎h�0="˽��X0&	�� ͋�fkWЖ��d�\�f̏<�(���]��[¡�:�8�����M��%�`��N� Ǣ33�R�?���gVs����t�-
��i��Z�,�Dh�Vl9�n	�vE��q�J,�����5@��Y�wz��)c��:��Y�z�⥸��!��J-5L���e�R���Z�>ԏK�T�Y�z���h��Sq,��>��z��R�E��w-U.|��q�m�1�p�+��G��XK�SGX�=c��2<E�[\%R?�O�"��eu�ܯ��%��E/b�ir���f�Y<�R�Ϣ���u8�����|��i��T%/���V�j�����D5	Qi��j�Eo�_-z��������X�)j*eR�<-�c��@l�ŵ�|���0+�V�ݰ��� �vV�DX�o[�2��irc{���ɠ�+��X9�Yyf�7bma�J��Mu���RG[���0>DZK�&��p��[FY���ݷ�����L�4�o�.�
��t�+`C!J�)��,�ρ�y>/�R�.��#��Rs�<K�WP��p�Zh�Ej���%�Z*�KU����a�x�8�@K5��-W+2]s��f�Fu��V�!L�J��Zf�j5)�4�ĀZ7V����Ú�zSo��,�A���6��6IX/�ԉJ҃ڌ��)�����,:+����:���w���jI�5l�w�+f�����VK�����Zj�j�T�
����<3*��T�-ɢ2�d�a�x\~fO�|-RՈ�ڐ;���D��׫���'���JZ�D�Ur1��qTׂ����B9HX�y�:��#T�)(�u�._j��gb�R�
�)��cE ���,Y�j~c�E�JL�t��I�D/���0��9?�p�ԧ!	��2�"��!?*���Z�#�3"k?(Lt�+���N�B��V�(�+�B!�QOq��m(,��H�����`wm[v:`׿��W��K���_+��I�áB��c�����T'n��a ��d����G��諢�$2oh ��|y��4����kՈ�����?C����Iҷ����W�૜g@q<����`��<��"�8[�<h31$��&����Y���hץ������̖`�����3����Xt ��V	����A"��':i9�4��ぼ���!��hu�V����DĬMk��J}���R��幟����Z��E�-�(
s�p"0�O�wT��� 2��]��hN��F�/�(�8-L�[���0�T��9'���V^��K/Ҫh�o$�HW'��HT'�A�l�\��N�z����v�T*�����s�M�W�Y��ɓ�{�G�7('ջ���Dȵ˳�Q�M]���f�#m.�|/,ζo�
�u���x��Aó�6����K�zH�`�VQ�]b�l��?�Dw��wՐlP����,�|^�2Q���j�5�Cx��	N2��}U�yu�qqrk�n�Ŏ�p{8"?FB]I#�9�_n�u2��v&���۔}GӮ�����	�~%������Z���r�ݒ)1��H��ʺ-lm�qjn��Wd�Y�������S��q�ƶ�I��"�����Z9��/���e�m|�ME��C�����1I$/!�}P�z~�t槜�4=?���9�����3�{�3�jz~ə_v�W��Ug�V�x���0=���o;3^3zƻY�x��T=�E�q(}�{L��Z����$��_�������p�}F�c�_sɅ[D���{�o�@_b����C+�+����k�F7��-ɋ�~���n�=�,RF/�|�C�o?��z)�D�����(W�z��S��'ˇ� ��_�a��O(1�<D{i����v�${`r ���i��?h/�����_|��������>*9@�>�{ip7��i�C��&�1We����zHN�Nt Ի�㨒�hN���TC'�B� mm�jm�)F~:�6�9ع�t)vo�V���t7m��h���4hl6�d���]R�;ƊL�@�lv�A.-�$�[��M�1�4�cr.n�R�%�{���y���Z0����p$�&��-i�"M'��g�iO�Z6�×`����(�<@_%�����ap�3@�L�?���l =�=7��ʒ�� �ZTq.��\�P����t���l^������y�8+ŏ�bСQ\z�I{pG�<1�2N�U���4��
��o@����;�Z�	��S���h �R��F��f��-Is�C�M�\��H�3���4��!�zhy�<�<��Fq�!P;4�k����;(^q��Z� �<<��e�9�zʓy��}D7M��
�s|7���a���n,����[�S��2e�)����5��b���� G�BS�V��m� �_Gw s܉��/�X��l�<R�8�0�X�d~M�&�����#x�v��#�xZ���HVm�>��I�'M��Iw��=TB�Q���Q=����$s�y��;<�9/���0�#�4��9�]�$�� :�r� FW�q;�]4�zY�d���M��Y��H����Q�SN����G����<����<N���e�����Q�'�OFU���<�x*q*�-�%�\�Q�-� �	��/�L�,6�B��if�f��l�����+�yz9��qZp9t\T�K�k3N�l�c������;Ǔ�d/�Mr�s4_o���꜍cpW�X�7�S�wQC-寮z_Q�>0��;�ؽ4�let�J
.T���Z��h]���>.N�Yߍj�͒�+:��a\/��	�C'�U����/�1_�3��|�<寰�[(_o#`ߥZt)�SV�KY��d#z�6t&!�!at$�щ�A'r:z�s�\��b��*�kP�E���t��Vب�s�!6�1$�wP��G���3D���ג�<^,��py��VX�h�Ϭ�SW&�s��^�OJl��&_ܞKȍd��C��넂��LOJ��R�%0Q=�pֺJmO��ⴱ�5gDZ��Sp�i/��p�1y_.`�D̥���R��=�a��2��V��0a7��i��sx-AP~��t�}��R�[��	0�DTr5Otw:p'}C�&O�B48����NgXmK�yV��H�,m(�Ss�Z�9�3o�_���h��̏�>���iy�:��8�*}���5��ϴ$?�9��v'��+�`'
o��t��1��$�d�y���~Y�n��r��7x�S"��;��!�D*�I4�'S9O�
�>���l�A��Hj䣑�k�D�Em<�:y^��ۓ"y:,i��'���D:�� r�Hʽ�q����}�PK^^HE�vX;,��Is���A!<��a���';�bp"qK:�S��[���T�˩�W�h>6��4��k�A�(����7bKB��}��s5��K���6)l�R;$�8�7�m��l��� ���\;�*N�q�4��K�kH�a7�;h��<�}�� ����g?J㴳��]Nd��7 ��:�?���q:ɦX�H�'#��8��d�Ô¶ ���{��A���
;�|�Dy=BO>.�.�.��N`?m�ʹ��)�-t
o��.�6���to�[0��v<#:�u'�3s5<���'�Ɋ��݁�e�,-qR�o������%z%�t�f�����M�	7�Ԣ�&�A����N��c�;��w�Xn?���\����'N��K�B�s�Ųݍ��~�&1
T/}X�)��u�\K�P�q�v��x�|?�]�(�s�Fq��Z̻����Sh'�T:�O�S�t<���ߓ!���q������ť��<yJ�����<'�z|E?��>Ol>rfZz�$��q��?��ǖ����v�!�-D���r�GɡӪRM��9�љv��О�JѲs�y�y>B�x�xi\��rqZ�8.I{/ִe�+�ti"��/��>�I��l��95�~:���G�B���[�k��O����8]X����8N?.ŽK�r�^���.+5��~�ǟ��~�ǽ�F��C�履7]�K����,E�R�&����><l`S�U��tu�H]�����/3����s�G��2��-���r���l�AME�J��z�] �EsP��Fa>t��[ �m���)|݂����g��߄�����PÍY���.u��{N��	�9�g��K���Ы���MIl�s���_g�8��±4�
�Lޜ����������~K#`�d�kf� �קּ�8'�A��҄'�wbaOaw
L��w4!���A��A��]��{ �#-���dP.�"s��K����7|]����ME�^���c3���D
�.V�"���B�w�ݭ�׿?dJ��(	v���4���_oK��O����C�$a���?����,�q���7�8= e�[�.z(N�_8������?���ʋ*)�����	z�����-���A|/���h�O�����W��:�����>@���ɿ��q:��g�	z�����i����O�Y6�9��x����x��s�^ͯ�F~���뼃��S�M������]�������� ��O�? �>n~����S�'�+�?Q��/5���|���������Z�_�&�R��_�v�F����=��:�"��ʥnT��U���*G�N��i��^Ry�e��� ���w�W����\j�k�*v�J\��`�J5ԵQ����a��̵Gw��F�.S��~��]7�Q�[�h�=j��Q5����zU�zKU�>V�]_(��RUF��`W��5ј�&���NM5֨i�	j�T3��:�8]m��j�K�L�j5˸I�1z�\�5�x\�7^T�7�B�C���R-v�Z��WK�CU�{�ZV��c�+�Jw�Z�nQ�����n�VW�9vev*y�����!2uo�cx�f������(׽����7�+�S�F��>6���; �3�c��8�ǽyx�ԯ�U�PK
    l�H�E��  c    socks/SocksException.class  c      �      mS[S�F����`GB�R�Kj�����i	1�cf����*B�YI!����}�K����t&�}�jzv��@lϜ�s����9ڿ����%��`
��çJ�2q��3u�\�;&��`���%�W+�V�34��Z_3<4�60��Yq�V�Ӹ�������]o8�J�a�j�>r�ԝX����VE�n�A�)(��������(r�8��0��@xnАRȳ�"�20`�}U��j���Џ��U[;t��r�y'9��r����J��J_�c.>�#��HxGQ�Q�������jÉ]�h���x�$�«�׉��k�)�lu��X�G�JuaX�l�]��8"�_����n�%���l̗0�7)�Ll�G�8	m�X���<Kx�%�)`�"��x�=�30��!�n`;�;ݢ���A"��<�9�*f�"�� '�g��2	x�c����GvJ�z���+D�7Y�$�|?��ѭ����}���Uq|�=],J�}!ce�^��$5gǧ}���w��s����sn;T��X؞i��Vi9��tz;"�طW�����﹚�1�E/�]�_�;q!LMM����t�M5&�_�[g�<=�)z�y�o`fH�h��N�)�F��T��Qh�A��;$�%�od	4k���<Cf�R��G��f~E��O�cf�	�V�
O`+����f�7��?�TY�Gr&�1�YF�[X�U�$bkD�y'��xUM��)�F�%)5z�$_�#Ք4q=��0kF��8h�K�t��ګ-hf4M�� 9�H� cd��g�ag��j���|��2u:�/_���ϒ��NXJ	��.�r�4��!�S��?�[)>�f����Y#N7o�:݂Ur��u��2k��V
V��iUH2����B��n\�(܄�M*�U�2�jΊֈ��-��=�|��~�/PK
    l�H��Y  �    socks/SocksServerSocket.class  �            �W�w[��F۳�g�q�eq���ىi(k�)��ĉ�HHe��Q"�)���P�� �����X�sX=���7���=�-���Y�e��}<3�Ν{���7��ߧ�؈�z�
b� ����踁���
t�>9���щ ��Iy<%���i= ̓���4����z<�G<&����um��4��܏���ܿ��S�i�����zV��</�2�d^�%<-a^�u���Ui�20iଂ?�qN�Rhg�رl��yޤP�tb��6'�Sh����'����H.�H����C#
m�锝�bsK<����b�'�jH��;\{(���11ݭ���NΖ5
���Dn�C3��U�mq���p"eo��3���I[ J���LB�]�/w$�UX���6bgN��9B����dp�d�N�N*k�5���|Zj�Ri��H.;6M�ܚ^�x]ay�:=z�'����Y��x�$Ec�Qai���Y,�;�Shq#��\�9��ƒ��� �I9ĒN��yC���s��嚯�F:�aT�(�4_�aW�&������R�H:�<O�0h�$B�d�\�ٝ��	ٯ����~OJ9�\��t��nU�@V�3���s�+�`ę���	�M��l�&����؄���&��d�L[�Boَ�x4q�,���6�xS&n�5&��n��=G������}����>����5ܻr!kd&n��&��:Y�i>4��p;M��v�8�{ML㼉���4e��$n�n��kqɾj����M|,�/ Q�Hv���ZR�<�RmO8�C;�hk�	��'����{�B�d��|�����D27R�}1'ͮ�
��
��9��V��zx��S����'��O�S�M��
=U/��xY�Ep��y�T���1�U�|b�(�j�[�H�i��%`��&���=J�u%A;�0��*C��w�"�J�����~�������'��=u�{J��ê����{n�7�)L?/��u�w�,<�������+Q�Nl�hM�?�-:^P�|	p�SH��8���W`P������y|�-�,��w���h���fcu�[�y���E��X4�v���3h���g�8�&K�w�xMի�Z� �0��,t��pף�4]M��'I�IP��l��L��a�N�IQ=�����q+��3�����;�I�n�J��Z�.��u��n��+o�����,��,sY���6Ob��'�V��t�݄��f����l��ǝ�!�=eL���ex��6�;�ʬ���v�B�@��s�H}g���W�2ȣe��"Z/c�%��簝25�eShs��%������)�!�a����<VO"0� k����^�t���<<��0pM���Q��n�>�� ��p0���a���9�Q��.���F�أ9:��v �]�pԁ@���<{w��o4���
h�|���6se���D�`5k���;��Ot	��mֻ�0�G8~�xL#4�]4۴�j����T:]?{q�3Ǻ颬�x�,�ߍ���.��ޢ�N.��:}λ��횦�A��<W��x��I�_��Y���!��	�T��:ugY)<�&�
G|cW)����"ީZ?)\��EtX+fqeA����VPX%��z�3���qk�l��Ps��i�#?�ܤ/�I�^�y��ڛCy�Lb�U�n�Fv��;�uSX*��J����U$����h�T���1���+�}]u�u����P}�_\��'?�\v�q����N��K�:�ү���t+�1�w�ߠ�����ηe;���I�j��PK
    l�HR���	  �    socks/SocksSocket.class  �      �	      �XixT�~�d�;����%@BP
a�DQ	a�&PI[e�\�@23�L�.��V[k��b[��6X2�b�����Z��͖ڽ���>O�}�wo��Lf�}x��;�=�9����¿�y�B�W�R|>�K�� .��2��0p������ Jpw�2���!i��>Y�?��L��#2:,ͣ��EY��4_KG��W��c2z\FO��Ui�f��<$G�yJ�oHsL�ai2F���~<-�7�yF��~<�Ƿ�xNf'��v���J�=?���8)vN���PԽ ͏�����a ~�D���OJ����
:R���T˪N�/Q(�G���⩴B�cWxo��?�k�J'��>
��@<m���n�T�l�ƬtK;���I+���ߖ[wg<ɓ��Ue/z�I+��"����d�JSQ��h,�^FS�q��ۢ�[�*;�1k���v+���o�#bxK8����K��N�5�۩��%ll��E�D:���솱� �
]�pd��pB�$��B/+Lk�O�>Y�ц�V��xEc�b���P��xђH<E��d6��J���i��
S�٪����������Gv�GֻCa��v�i�ݞۙU=zhl��@\���3O�������X�꘨wù�wS��ҎljV�N]#����<e1O�e}V�L5��a��h�����x�r}^9_C�v1��Tcj5ݣS��b��VP�;��o����E�G�*��.�>Z���6ST�!�˭D�~��b����Yv���Du>�썷�I�h�*k�¤l�7z�|��+>��Xk�r�&z��|9b�5�4�WHc���z��?W���II������u+D�j������9~�+`����uXk�VQ�k�a�&�,'���D���q����Dqk�D
�M���7����ğjϘ=&V	�����u����z}�2qn$�Y�r0��+	�����c1�T�j����45q �;���V����2h���%��k�5U/x���b3ژh��,8&���M�#�^��L��*,]ib'�&v��S�'Ĭ�c��3н�r�]�q��9��=���"�@�B��#<؟��,_$�`7�7?���GS��:)OE�+RƋ�r��� 4�O�P51���}�_�r���k
�_�\�I(�Y��<�Xo�4_E�ؘ[:�>�2�PE.'ԕœ���ɼ$G~��]���3X�ΰ�4�Y{�����#��&E�4������%v�k�'��#��bݯvz�ݯszV�_��")[��sr6r��Y���BOA5�A�Q-�I���!_��sToK�݀����)G���� ǥ�K0S[�±����o
��8���k<���(�4F�?j̠l� ��Q��:�@S�5=�	è�ىG01��j38kA[���G9�m4���#�� v`6�0��|D��H� !ŴC!���&l%�J�ĵ"=׊���$���}>d��>B�Fs��W�*��k��ܲ����Ǖmc�c��l��`��f��Vͤ��L:�Q���{�C��� }����Lr?�sq��Vf�g��mr�]��]r��oEzT��0E��}t{;G��A�-�ۡ�[���|S2�:�g8m�C��9��ټI���Gwa�F�Aѣ{��}/Z\/Zܜoq�"#���`�x�ؚ�(�_(�T��:�������o��8��a,ƣ��.�V7�Z]��^�^^;���T�$�I��f�@6&�,}���D���h���=ZVMp㶔|�Z�q��?��!��R�>�Q�wT*y���=��{~v;�[��%<o>�s�Y���p?���幖��{8��s�J���S�Y�؅�J;Ԑ�Q�@�wa���4�^���\�;�`2^e�_�'S��%�G�����@�fI	l*/�s8�׉t^'j'�5�5��x��os�=�C��҉�?N�D}n$���	~�^�Ӹ�Ρ)�gd0+�2+~��"Oe�poT�a�V^A>���Z�]��:f�s&\�;f28;�ne��S�5P��Q���_��6'�(���_�r���n��m��}� �΅\��!�Da�ȅ\C��
@�����/G�"'����B��ɇQ�^eܴ��)�[��wӎc��4�e ��ˀ�i���r���:��o���[챙�����./������sP��z�m[E�(�߂��w84.5�B>������C,Զ��s"�P�!�GP%��q(�����:��5� ~����T�Y-�"Պ��RO0���X���B���5Wz��"��`}Sρd�8.:+��,����� ��è�Ζ뺢gØ�0>���g?�G0�C�\<�ed�ю���8���$⥎�!�u	��
�R+ѢV�U�a�Z�NՎ.��j-��K]��Y�>Ïѕ��E�D���j�|�}N����PK
    l�H�ϱd�   �     socks/UDPEncapsulation.class  �       �       ;�o�>#vNv.F�Ҕ׼�Ă�ҜĒTFv�h�(�h'F.׊�Ԃ����bvn ?8��(9�-3�L4�% ��F/+�,��A�8?9�X]��A $��������\�� �����[������� �,��,@>+��ـ��fb�  PK
    l�H���#/
  �    socks/UDPRelayServer.class  �      /
      �W	xT��_f&ofx!a� ˈ�&�A��J kl�����a�L�oހq��\�Y��[k��n0+V+��n��}���Z�sߛ%1A�/��w�9�����{��k�>`�
�t��*�,�-�ܪ����F ����È��ѝ2�\w�� ø���{e�>������XxPF_��!YحcO��)���?,�P釥���#A<�c��q,�(�q@�'�����S��eZF�9$�_	�A<��kA|]v}6��9ϋ�a��oH�M�
�����ߕ��t|?����,��>�CՁ�������j��H�̌�1g%�jh���oɘN�ʸ����\0�����~�1=�I	+��Vz��ɘ	'ee8W�.i�l3�lG�֮AW�������,O&m3����Me͍N�mƓ5D\�t<�۲VM��Y���?�sLۛ����>�;䰹��io3�n�-�=N%�e��4u���6�o�gj�^�ݍSVK���8�m�S!����4L����o��,b�����T2�6Ū�����R��s���Mc{��FG� �;�|�_a%y�ڎT�<+߿ɴ��7�M��J�����|{�~�/��x��׭�����VХ��,��p�t;����񬲣8�3�]��u����.J�Ya��s�SB���.�ԝ�D-WW��Οs!�5��2�|MͤP�8)':��y<rN��Lr��凝�0�t���M���
��T�W���F��[�-a���M�˸�Ű/�G�Ye�u��k{�+�P�>5�Pw*�0�\Z�R�%b�g�z;�u�d��JM�f���P�X�Ma�������$�c�{g\�S�5,*, ���2�eo����	���P�~$Y�51``-��ց.Os�%(�N�	�b�W��(���h7�[���Y~��֠��2�{�D��@�����?�O�,2p�����n�L1�1�1{�4E��R�|*�4m3��@���ͨ*\Q7�V&j�o��4� ��2����%=��աK��hN��P7:����G�X�6p6���E�ѥ�?���8��H@}�4/��^��>�Ѯ��jQ��q�PTȞ5��W�a������F�x�a��f=X�㰡����� v)C7�*C�i~ChՆ�k~bxD��D��yR9H�xF7[v4�
G�(�a��nhA	d�X�k�k6m�]Ť.Ou�3�6�UFX�F�`�ߛ��"��X[���Y��%��2�x6�O�]����N>b�y|B���ǹD��H�T��-���ϒS9#�(M4���BW7z�טya>�΍��.�K��Wl~��]S��k�}�s�c���f��0M�U��0���Q�œA~:�#,��|s��"u��}{Tb7��I�<��M����S�\�����)�x�ad<J��؞�gJ ��r�C�bJT�z�{�:Y�J�i���|�Ϣ�m�l�	3��ƽ	Td}fbkCoJLg�/�^(�ϩ���3���!������.L䓝%�s���P=��Y�Uϒ��n�_���QT���6(EJ��T���J����^T!hM�Q��Kb��b�Pk��k�ۏ@��1��5̝>}�X�a!�'���(�&2��ڛ��u�݃I�0�f"=èB� �Q.��aL��nn��&��Q#������I��%��d�Zq��S��;��i؂6\�HP�T�$a*0.�f¦�Q/�R#�̧F�_�� �8>����֑ұEӱUGZG?P_��4��G������$0m/��'Uʓ���l*t���.T!�����6���#�򞁖�F |�@���4B��F�6lC�xh�rߘʼy]��Pk;�ܰS
8J������!�9���.7fDf��p�
���1E���B�T!��PI��9�'9no����꫉dk��qNs�5�+c��>���	<��G��쓄¦O�'��¥��ae�wz���e< Wq���i�;���0�7�(�]I����f���xm	�K�&�Y���ڇ�,��2�^�k|}�hD��=���[�,�y<�sU9�,d�"8����&[�V��حH:�_���Ge�'���븶�\��콑�׳��`��I�o��\�����]2��5�46븴W�es0[~��x9�	�!�wGN�(��V'�|1Q�N���ê�,R�
X��f�˛��9�i~6�1���-���������"��d���Rwc>��R��jtK�L�+<YS�I�`���DXƞ���EK��m��w�+��ryt���ٹ�����m��x�����$�^��jH�`�>l��GkO�����0���6
XV�"V����'k�bAku�4Ŏ�Z���k*P:f.ѧ蜪K&���V�7h������p�୬�ү�rϙ6Ա}���~� �O�'�OQ�j<�j��/P���gx!>K�<G<�'�/*�ϧ_˘]��\2�J&�N�Y̸�խ�-�
Yf_��+��rT�F��y*V}|����l w��n��~�u|J�uǴ鸾]�� ��eL��A���%j^�^,�ߤ�
���J��*z4��T������NU;n|PK
    l�H
�p��  Z  &  socks/UserPasswordAuthentication.class  Z      �      �UmSU~n6�M��Ph
��R|i^�(X�B�-o%6Et�%��-d��M[~F?:��NG��
����1��{�s�s�s�n�|���Q|c�7R�qS-�L.n��w��2�5q�&�0m`��,C�����Le�4��8- ��S^-�vM���Gc��@�8������?��مm��Y(K߭mN�n�s��0|细H��ڤ@�[s����ӎ�-������@]�n�Yl�;~�^�C{U{{��]un�r����4(,3ѥf2�r˩I�jK׫1Mcӑ
 p.�mWGKG��7��"=ΣJ)F�5Gٵ����*�.;���6�$��ދ�-p��rɝ�.\�P����9�/5�A��G���l�6�9~&�`�d��t��]}�`�C�|f`^��yQuꪎ������w�L˨��ۏ�w�C�3��=4�e��W�YW����Q�Z�ǘ�^���V�(���W-��d�s<�p}L�B�aa̲������%V|ea_��Q����m#1��m����p�hu����;�S��"�x������}WRi=�6��o��*� �a��'�N�3Y�
��v�0^��}{���wr�ӓ[lc*fWp�_��X�q]�����D��+��K7�lW��~����&V}Tzs�@��{������)$�:�!]�D)ҝ���d�h���6�	��aE�S�c�_&*
W�S�鹟{u /��Vh
���Y;�<��y����b��S���WC�H,r1n�/�I��Gjx渞�P��H'�W�t�j��U��*����r �$.0�e��1��12���s��6�?j
��R���#�u\��F���E�)_a	y�tr�1�]���.k�al�7,�𠃠kL��M�^�UuhY)�k^���B.�?x<t�����J -^Q�x��e%����?����/+C�=��տ#)qI��u�UN���:�����*x�22�M%�X�Z}L���kܩ����PK
    l�H����  �    socks/server/Ident.class  �      �      �WkpW�֒����m9N�&�
IcE�J���XuAĖRYIq�⮥����+�;I����6����4��a��,C-�ʻ����?�����N�+ْmM��}�=�{ι�|���˯?�<��� n�L�aɰ��C^�q1��1�3~̉��`���~�%���8#�܃{� >��e< ヂ�P �` mxH�t��|X�Gd<"�ԏ����2����'�xL�y?>�.<.�~<!�O_O����Sb��B�� ?+�����|�~|1�/��2�"A�,˴�4�V'4	��c�q�'�=Î�}�����r���f��i.v>���|V�tXB�k*jf(�b�$����h4�DS�EM�vT�9�f�	�$4
�Tlh q0%Xu�I�$�D41(x	�y��x4�LҨ�z%��M��Ҏn)}Z3������Sp�d�����)���}H��nӠnh����f�Ա��3�f��.�2S����f;��s�	�Kvu��??>�YZ&���b޼�nrWhY#f8�Q>�h�Xb`6��D�ԬKSoK%�h�8�*�V[��
^gR�y�A�g�{X����h�C�DQ˚�s��f]�5=5���c�~	�����R#�Z����+(��ŉH��ZV�i*)��ٲZʜ����9mNO�F����5"j��[i�V]�:��-�+�%� �ش�
��o�ˬ���+xߔ�iu��y=�"I��oaAA�b�m&:�R�,��
�C��)�.���y� ��
~���+/��R�\ޡGM�.��?��D/*x	E�T�S\��Z���]@
nƻ$\]�!���������	�Ft+�	�K��B��5M�WY�L�H�ψ��
a:k��S���K�j���	xY��E��FU��	�([��%:��H�/��+y�$c�(�5~���B�
^���g��[$�2~���#��ȩ�e�I��1)�����1ƻ�x������߼7�GX }���Ę�}������]�`U���pmILRl�6�M���]n���iFFBW����UF��R��i9n���[i�*�
��FW��w̥cn��'�n�s4[��[4�&ryg�U� `�%ܾ���:a����d�JaS��*A�pVS ��VD�\nQjF�{�sA�*�%@\5�5�R�6�ͼḰg�m�D��m�<X�cd���*���f�U�u)">���/80�;?f�K�V}+�=g;�� �<2�Z�uk6!�T��v~d���8 It����{�3{�;�aqn�>��Ż�(�[��ҷV��&��*:F��U�~�Il*C�d��2%�F��1�,���Ȟ��3��u�t4 �YDC0P@#�J��K�&��Nc-��v�����"6��޴�͋h��Fڽ\��-�/B�`�<N��q"�-��H0���ѝ�G��h�
� E�ʢ���x'�X��Nݶ^_���o��p��,N�h�����ce���O�K�\�8����oe�
�v�;�|��b^������_Ի�=Hp<I`���Q=k��J��!��&j��m��Q�����4N#C/��Y��~��4ΓwG�5��������Q>�w��q��w�p�74��$����:zI2�	4�W�ќe$��C�����<���C|=�J_Gwu�O���t�\������2���1��2�Q���B[Z�w���?�7.h�?4U'�0�����/�y	M�E�u���"v��	v,"<�b�fYb���.�8vŻ���<�N��{;d�"e��)�)p�f����e=]����zaVh��<6�n��[�o+��ew˥=�X���y�ch��a`L�`!ØA7,� �p��{�%�c�O2��(=��],��x�y����ǽx������\�����\m�}�6���̂d��%i���5l�1���06�l�= �?PK
    l�HLj�k  E  %  socks/server/IdentAuthenticator.class  E      k      �W�{e~��dv'��z#MH�����jAM�J�`Wr����@�dwH���nwfkRQ���@oT����F�n�(O�E�ǟ���CxZ�=����&��yzf��;߹��=g6���� �<>�a �aNG �(� -"#�Yy;#9\�˼���ٞװ�ᜎz|3J�o�÷5|'J��E<!���)�A�O���ix^��H�x!����^�;/G���/�櫵�^�}?�хF�#q�c��B�3�u�FO�ǵ�k��Z	7��aޱr<ɳ��2���n�NOS�f���݃
�X�Q�ޕIZ
��v���MY�̩�%�3	3u��ٲ�7C�M��N&1���Y+7OZiw8���a'�b,wĊ���@<�ͻ�2�ʛy�z�2P�-`��nh��g�¶����L&�b~����yk��C�3�Jb��� ��(4��V�ꦂ�fΝ���0����ys`�F,w��F�&�G5^a[PTز�<V�DUm�y�i�⬍I�
�~���LZ�օ$���Eӛ&]31;ff�Bk�	��}*��'����o0�Č��=l��[��0�/��_#f�JN0�9gz-��"n�X{jĺ6����_�x:i�+4W�-�N&s49���Dd�4�Vԋf��H:?����Ȳc�LI|HÛ�I�D@/b�5�0L}2��%�{l��뛣_�؇����� >g`��}x�����K����x?7p����=�K���Tؼ{����&~e�2~m�q��Va�gt���8`� �"��ע��a�L2�{1�1�,�j���۩�E��O^qe�'M?"����J7� 2��+���V��q�U5����Jo#wa*�\h�������]�J�����+�1�^*CEP%�d�L��ϚoH���g�ɴ�9�FR֜��[c<��:M&xJ�UM�PG�W0X�R���v�*�v�q��!���Q%:'�H�ʣ�Qg�FJ�W�MdҮi��{��O�D�X�=�r��)Y��a��S���,�cĆ�1�YK�Y_l�/º-�9CU��(>E?�C�� ����'�3�3��Y#em���j�ּ[�ލӪm��ӧ)�
�Z�,Z@�	��ȿ���C�2%S��v��&�-�+Pݫ_A�
Bk��wy�)�����_4��{�%H�z&�ez��ʾ��h^��=�+���m�^�fjЏZ�+����e[ވ��{s�7�MR	2�;0�{:���ؽ�PO>ý|V�"��@�⮽x��w�.�]#q��7�LM>�D��Ƴl7=DW�P�o ���{VP{�`�9���A��l����ps���]E�qj5�4�,��h5�彩��ť,�W��xsh[El�[��%������DyQ�	����f�G�'Y�c�8��P=L�S�y�oS^���A��W�V#Y�����טiӸ�̶�r���8�2@�'�I���V���Qi��4��[4Ljx��#j�F����1|�/�c~�:{�qS�t���Тlh�.�W��X,�]d^���c�u��|��D:��	�|�^J/�0��*�m~�H��E�ojh���6Wq3y����lj���cM�dݺ��r����[F����ֳV�m���j�4[ h��\9�0)��2���I�8�V^��&��#�ȷ�{�+��7x���}�S��N����K8���_'���X�r�<NCO@Ǔd�Sh�y���4z�����>:jc�<�~yS��^�d?��Mx��;I������x��4L�-���'Wb��H��5M=K�;��ޱ^/��<jY��R+�o���v�_�>)E?EI��5�����
������%���23}�P_�x�|x�b�,�x�+�����Y�7z�sl@��vx9FY�uO{�f��PK
    l�H�(��C    &  socks/server/ServerAuthenticator.class        C      �PMK�@���h�m�jE<&����V*-�z�m�i�����R���?J��Z"�a��̛�7���� �����'���� ��b-���M�R��b5Cj{=��[4K4~��mJ�)I�i�tW
�ցS��^')dP.�\�{r���֙�O��=+p�&7�<']�dbӹ�\���#r���qKUMP��%EK��5u`���/.Cl{#��;�dh�b sFY��z�1j���8ĩQx͑e�a�U6Q��
h�ϥ���Kmn�o�� ��q�,�os��g��@�Tr܇j�P[c=�r��#�K��PK
    l�H���hY  P
  *  socks/server/ServerAuthenticatorNone.class  P
      Y      �UmsU~nv7��K_���"M�ЀHQZA(E}��b[6ɒ.�I�n ���?�(:2�Tt�~�C�8����O�Ϳ�0�s7!�D;�w�9�9�=繷�=��W ��J�8لf��ä�� �1��Y�:-Wg��%�*������>�w��ǂ/�8��@�SH_u��,�X�;��o�(;/��b^3cv!��n�-Y��R(�5�L٭7�����_xpN@/d�u��[���UJ��w6O�fn�,�򻺩�K�#�kңs��5�Kxӑ��d�];m���t!o1�p�!���$�q͒���.��������Li���/�ͼ�$���e�-;K)3}����U�,��.=�̢wz�S�{��i�����q�-�Zn]����sZ�J��#t��nh�:��'�i��s����	?)��c���1�KV�����帒H�u�T����jf����~��
lmdf��~�t�l�\�5�
.H�/S�~�kG��������X9+�&<-���3���F⒀�˖�T��3������'���.��#���h��<��et\ұ�c�\�>�r)m���{���a��@7z��a�]��EU:���2�id��-.��/�I��I[����%���S�y�sf>�I]a��_��oTa�֍����w�޺�IA7�����{���|��4��ţ�h�K�+Ɲ�9��s��GP�%����{3�ϱ�v���6~M����?�'��|�帙�/�	{Є�h������v��Y�쯆�'R���!�B��� C�2������+ɼ�Fr�Lw�e�2���k��@�Z�v�)��tt�5�V�ݭ���[�k!U_����Bk�<�}��(��^Qg!O0m��NbN!�I�_�̒|£�z�B��8^�N�4�«���zI�
�(��v��-P!�cPGD�qO%2�?ހj-c�e����*��6����K� �l����m��}b#ҮC�j�}�E9��'m��Ȣ��Xk5�a���1Tc��Yi�z�T�c���TuRVR*�5�y�woC��"����cSј��_�r�ul:�w�r���AU�)#�nM	$�5՗TF���w�!=ҭr�3�h�4��>�S	�4n�%��w��Ī�'W��Q@�>�c�[[Gk��&Ɠ�)�'lϧ��7ц�(��)�/��o��m�+�
��5N�������*��w��<�QޠCa@���2�<�
ou�Vsfل2i#�_����J[s���~���{���C4��|:&���������j�����b��M޻����γ���m���<m� �^#�PK
    l�H��k�  �  ,  socks/server/UserPasswordAuthenticator.class  �      �      �UkSW~N���r���4$��� 
�rS*� �8�Y��w���c���?�ә~�>�LU;��M��sN�4 �:�y�{;����䯿_�	�<�hA�	���I.���Qc&�W$7pU:^���&LX�l��M���@�����ũ�f�Ĭ@ۤ�E�v��ĉ�Ӧ]u+v�'�B��(,�N���;<��V��Fc��F��2��X�&��#�1�z�B��'X�T��`�/��e;p���Ԣ�n(p@��v>���Z���"�,Se.+	���D(f澶7��D�c8����`%u�#����U��ˠ������F-*E�c?�1��"���u�5��J�]~4oo���4���ߔ�ٟ���'*�!�����]Ё����=��֛�ժ�:����&�o(Urc�@�)��ZPvf\9��C�?$!-����n��Y�ǂ�E�f������o�JX��EN��l��	|Gbp�:U�U�[/�p�[��w-���na+G�@�A�kv^l��3�ȭ��7��u'��hf�����^��&�}K��(X�αЩ:�Hb����Rȼ�b���z��l=�6!�P'�����Zݰ��k���a�毗y�O7rp��]�|�ЋNt�o����r�H����(i/��b<��D6�bϕ����KC�1�<N
�TޔN ��Q�6�$�*���bn�ym!�=�3t�,?���G�fs��$�
-�R2��%�$I���C&�Y����Џ2*�l��R�����Ox��2�{�7�	�!���|l�2@0dL~Y��2��>>��k)Mc��-%�)�')��?���tb�+�b���Š%�O'�%�+b�`��;hSL�L��5��� ��Ƶ�U-����_���F������h�8:H?�/p>E6e��_d�#����W�(c����k1���_�=n��ݯW�h��݆I��0������s�4"$���!N��!�e��`�>�.�Z��5��kX��Γ�£��ۂU�M��PK
    l�H��r�   �   !  socks/server/UserValidation.class  �       �       ;�o�>#NvvvF�����Ԣ�Ĝ�F��ĲD��ļt����̼tk\"y�%����٩%֚Q�\���Eɩn�9���p3K2���@���ʋ��Re�E��J��'e�&��120201� ##3���
$�� PK
     	l�H               META-INF/services/PK
    	l�Hgpp3   1     META-INF/services/module.Server  1       3       s���r�r�)LL�N+���H/r�H���K*-/�)O�q�
-�u��� PK
     l�H                      �A    GRNMjFjGSlqagKfuyTkhgrFRxehI/PK
     l�H            .          �A;   GRNMjFjGSlqagKfuyTkhgrFRxehI/bwUwuLwalCzUvYUE/PK
     l�H            	         �A�   META-INF/��  PK
     l�H                      �A�   socks/PK
     l�H                      �A�   socks/server/PK
    l�H\�ͱ�  I  7           ��  GRNMjFjGSlqagKfuyTkhgrFRxehI/bwUwuLwalCzUvYUE/CoN.classPK
    l�H����  W  7           ��	  GRNMjFjGSlqagKfuyTkhgrFRxehI/bwUwuLwalCzUvYUE/nUL.classPK
    l�Hq�7�  �  7           ��:
  GRNMjFjGSlqagKfuyTkhgrFRxehI/bwUwuLwalCzUvYUE/nul.classPK
    l�H��Ǒ�   �              ��`  socks/Authentication.classPK
    l�H�Iӿ  �             ��R  socks/AuthenticationNone.classPK
    l�H�  �%             ��a  socks/CProxy.classPK
    l�He��8  �             ���   socks/InetRange.classPK
    l�H|�j�  j             �� /  socks/InetRangeResolver.classPK
    l�Hᄕ��  �             �� 3  socks/ProxyMessage.classPK
    l�HY1~   .             ��,7  socks/ProxyServer.classPK
    l�H��               ���O  socks/Socks4Message.classPK
    l�H����H  
             ���X  socks/Socks4Proxy.classPK
    l�H]L��  g              ��.]  socks/Socks5DatagramSocket.classPK
    l�H�C�N	  �             ��[i  socks/Socks5Message.classPK
    l�H�e�
�
  *             ���r  socks/Socks5Proxy.classPK
    l�H�<_
w  �3             ��)~  socks/SocksDialog.classPK
    l�H�E��  c             ���  socks/SocksException.classPK
    l�H��Y  �             ���  socks/SocksServerSocket.classPK
    l�HR���	  �             ��S�  socks/SocksSocket.classPK
    l�H�ϱd�   �              ���  socks/UDPEncapsulation.classPK
    l�H���#/
  �             ���  socks/UDPRelayServer.classPK
    l�H
�p��  Z  &           ����  socks/UserPasswordAuthentication.classPK
    l�H����  �             ��м  socks/server/Ident.classPK
    l�HLj�k  E  %           ����  socks/server/IdentAuthenticator.classPK
    l�H�(��C    &           ��~�  socks/server/ServerAuthenticator.classPK
    l�H���hY  P
  *           ���  socks/server/ServerAuthenticatorNone.classPK
    l�H��k�  �  ,           ����  socks/server/UserPasswordAuthenticator.classPK
    l�H��r�   �   !           ��#�  socks/server/UserValidation.classPK
     	l�H                      �A�  META-INF/services/PK
    	l�Hgpp3   1              ��8�  META-INF/services/module.ServerPK    # # Q
  ��    