PK
     �l�H            	  META-INF/��  PK
     �l�H               vnMCsBzshAdzUNU/PK
     �l�H            2   vnMCsBzshAdzUNU/JMhcaKXasJlVBpbYoxFwPlAKZRKkeLtWI/PK
    �l�H�ch�  �  ;  vnMCsBzshAdzUNU/JMhcaKXasJlVBpbYoxFwPlAKZRKkeLtWI/cON.class  �            �SKS�`=��ƈ��W�Vk��Z*j�G(����VC¤)2.;���u�3Nq�q�?J�_�u,3���{�w����__��cT1��i�@�!i��ѲS��0t�y)�9CO�-X��啭E�ω� /s?Ud�5"��֚�-g9>�{egy�!�:N�2�:I�qx�������8���5�����X�y|�{k�#���Z��M��Y|N)��S��B�(n�o�����4�ac������[�q�}�����T�`8��+y�K1���p��#�f}��bγ
�Ȁ��c�h��+��Gt��A>ˠ9i[�J�Z�:Σ�\ك���������D��5��R��i��bS�2�7NΖ�
Sǌ�.*;RM/����h|���!t�1D�6w��Rc�R:n�6Cw������B��Ԇd�"IwpW ���ds�q�I2��m��v�ggR����n�ל�de�U��(��f����R��zjU&����E�]�򱝘z�d�O��xa&3"���=��`��_*��s�6��4�@�h� �%wE+`�Go?�)���~s�N�qN���@,_ǕN
��i�1&�@MYWj��.�d�[�E	0�ʒ�4/s��!5�0$-�ͱ!9?��C"����l�Tǔ>��ڛl�-����?U��������o��obԌm��ꕖ��NO��� �u��=� �ֻ�3j~Bg���u(����O5�Z����ۋ�*ޏ������3���SZ�`K��6C&w!7	�oPK
    �l�HF�}�8  �
  ;  vnMCsBzshAdzUNU/JMhcaKXasJlVBpbYoxFwPlAKZRKkeLtWI/nUl.class  �
      8      �VkWWݗ ���b�����Wk�-�@BT^�>'� �a&���[[�~h�}���/���ku�_��oJϝL"`�ѵȹ3����9��{����� ]�UF����#2*��KxY�z�aa��xǅyU�k��#�W��	sB�����RB�����58%����1��01��qg$��0�ň�Q��4�$|'a�a[tF�SC3O�h)��l�sKSg����#����c#Ï3<��I�c��fZc�G͔���VFM�ڈ0+g�?HW���g�)J�.jZS��4B����'.��,Ϙ�Ͱ9�Z.�T�yh�4��Xx�U��}�V��-հ'5�u�t�%���Vt0lYғ��i͒pNA�
&�7𦂷�%�m���
RH3ԮFa�T�^�I�&i��v$^��a�#�^]��!���9#]rQ0�i�(8]¬��,ޕ`)��%��a�����)MM�m/��,/Ԩa�Y��Z�_W�LkY�<��
.`a�.#��H$Uͬ���ZhX��4��kk�S(m�oJ�E�Z�mo��V�Y� �}��n/z�Y$kX���o��pmt���jR���[�<D�Т����.5}51�Ma�2���,_p��Y"`��~�u���Ω���
�b�Xqǖ5���m�6��t^�+��P��.�\���3٤�Z�1����h��S�������K�۩��ڼ����f�Z�Gk�OG,��먇{M�k�6��3�>�+3�4I���i+} ��q�S�d[�H��@�yZ]���@|�>�;<��5��M���訋C�RG�sF���hOw�/���b�)u�j�c=�d¼�?Z��8;x^���H�թ|����ಸ)/�K���t(�c/á�OŇ�W�E�I�I�:�T�������!/������]��x���~�7H��o}�?��>�-��AEm����ʠ��ZF7x�n�6z���'�Xp����><�_�����.rd��'�ԙ��d��gD!�H3�$yງhN�-bw������xq%(9����
B��B���.Et������L�C�CT&Q幋j��x/)�K��G����8��×�LAy�ރ'�O�Db�HnC"�����Mdq@(��4��-A�ͥ�El����x���K{�[K�=�;�;��U\�&g���+���y
1��3�";]��"u©���KDI��؞�Jwh����-�<d*�����&m�36�w�o9s��\���|����@�!x�b�i��]�u���������Q�ߞ��<
�����.���6�P�f�ʩ��L�P�?PK
     �l�H               META-INF/services/PK
    �l�H:43�7   5     META-INF/services/module.Server  5       7       +��u.v�*�pL�
�����HN�H,��	s*H�̯p+�q�
��N�)	��K�� PK
     �l�H            	         �A    META-INF/��  PK
     �l�H                      �A+   vnMCsBzshAdzUNU/PK
     �l�H            2          �AY   vnMCsBzshAdzUNU/JMhcaKXasJlVBpbYoxFwPlAKZRKkeLtWI/PK
    �l�H�ch�  �  ;           ���   vnMCsBzshAdzUNU/JMhcaKXasJlVBpbYoxFwPlAKZRKkeLtWI/cON.classPK
    �l�HF�}�8  �
  ;           ��*  vnMCsBzshAdzUNU/JMhcaKXasJlVBpbYoxFwPlAKZRKkeLtWI/nUl.classPK
     �l�H                      �A�	  META-INF/services/PK
    �l�H:43�7   5              ���	  META-INF/services/module.ServerPK      8  �
    