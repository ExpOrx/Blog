PK
     �[�H            	  META-INF/��  PK
     �[�H               _024_/PK
     �[�H               _024_/resource/PK
     �[�H               qZMgjTcHLmV/PK
     �[�H            #   qZMgjTcHLmV/eZMeHmHwZscExclOFqAlhz/PK
    �[�H���}�  �   _024_/resource/RDPWInst.exe   �     }�     �}	\TG��02��C��# &�d����
&H\x��x�>f�3	����fw����fw�jL6�a��&�I�8�%������� �����~���3ݯ���������߸8��i9��9#�(��cfn��4��ą��N�w��,���ڬⵕ��+��(X��V)D>RYa+���UD.[[;cXP������?K
�-�r�/}��urOWk���{x��2R؜�!o����/����u�|�Q��OG�M��&����s}aXϏ��!��v��V��t�\�-���<ע��jӅ�M���+������万��e���" �A����@(��&��(�g�8��G*+1�\
_��75�xkA*�]*��[�J)=*��<��*=*+���9?�g�^QTZ��c2�sC��#����k蓑��c���� Z�Y:#������MfN�X^^ZTP�A��_jAie�Ua+��|�R(Z��s&�h�s�*�&TP\� M���@Y �p:�ќPx1�5����
a~��U)���[����+(-�2������e .z��EK��^��EC�o��e��Cۗ`)_�*8�]�O�M*�(\[VP�����G��9��{�LUJذ���YX�=�S�Q.����k�--¶��Y��I(X��4�P��r�#�E�y��$�**���<γ��/��-S� r@���Z��Á�|���"�/���\�G��k�B��� ׆���0�J��%
����l�6`AA���@��SP�� ��v<��J*-��l����0ϴ����EY��s�C���e�O��F,�N���&�h���ĳ��ɟ=�23�gO3����@3�h��Sa-XS�R&T<�����a{Ƭ�e��\����??Y˝�ƨ����*��r���BH���Vke��@h]�A�׭/�W$ u�K��PU�)/5Ç�B�����{��W
A�Ϥr
�˩6 �k�*�l�?CzY�����B��O��K�O*/,b���d��X�0�<�6|6�={��0s^�i���e��c�O|r�>Q�f��-�X�v��&s��Ӑ&B��I�v�Ϸ�di�Hߢ��i���b�}j�35}SM�Q�i�ޣj���~�����5� ]���|@����*c�`ڧ�hzE�M�*�hzM1�Ŵ_Y
�B�>�P��b�
YK))Z#L�V�$��*�
�"�:a5�*b>��Ԋ#�=X|jE�O�<Ƚ8��ek��V
ek q��w�Wq�k8�k��uAmc�{��?��dn��:U���bn��V�3�B⒂u�h
�Kf�j8���q[�N����J]y~TK�j��p�ފ�������*B&ey��_f-�Q��q*����$��v3��[���³(nqQ�Z�2��|�OpN��p�s)X7�3d��aLA�VUVz���r�+�C��m�o��,�T�P5�U<>�[N� ��:`Zu�fs]@Ő����G��7�>�+���j���,03��>镵�6khMf�#��Ӂ�1���4s���Pk���n5M���r1\�͵���q��o9Ab��PA�:��*C,5��)?����MC{H�4�NM�8�J+�,F�7�g,5���r�b��7���Ԯ�fX���;Kٴ�h����LǕ��B�*o�ǌ�:��\���3y�r:�
�L*����a���е%4��Z^Q�\��+�хH���r}���؋wSU7`1LǂG�t{��^!�E�[)ȵ����⿯>�.|�K�6�l�oapp}4����f�n��О�?��h��$���,誃ǔ�p�A�}s�uC�s�$U���O{PL�����=�q,w̗;���Ǚ�X�$�3�D.m܀�p�Y��>�7ƛ)̭���3w� ���g8_ܗ���/�3XO4���M`jF���0�Q��"�6�-⏏g�v��U�$C�w3��o���տ��7U�BY��f
�'��<���������
��Q�G^�Uu��^�p��_j�
0�jk���Y�e�]��	qNXHH8�s+*
O��C�K��jH)-ZK�*w�Xh���7�j�]��7l�Pz4�W��t�:������Ƌ��mjl�D�}4|� ��6`���Aj� �ZZ�h� ނU�q�ת6�����<�VFCf���M�ycʻ��κx�#O��gn̒_�R��	�(�,��PT88��G;> =U>6s�g��5p�rY�*, ���� �Š����y�P-~�
�����*.-ŘP�.㴢��j�5��L)����L�nTU��]�XY�F�ꖺe a�����L"* �[-�j���e��P4Z?u��l�cģƸ>�3�����|t�T¹��0�7^JT�YMd�R�S� �C!عʁm;m@F�FoxV��Й�,�<����"�ۙ�F��~8�AΛw����MK���`��b��	X���S�MeCBq�vb��-wx�����ʃޏ��?^U�@�K�՗�	��EkY\^h+-zy���)(����h�&���K�6	l왍u|�����P8eŀr
��*6 ��P}�W.�"}�WY�o�p�Y �F?�hM񝪭*�LȰ��eÇ/���;�8�/Ӵֺֻ����.c���ڇ�N4��R�:�N2�+w���gjڢ�մIM���SM?Pӽj����R�7��5������&5}��e55���jZ��O��5�Q�*5ݢ���TP��jZ���jZ����^MW�i��f�)���o��OM-*|��v��j*�i�Z���f5����h�)���� �F>*�,9�'9j�F�3�YM\����.�/�]3պ�j:���x�k̇�����ő����F��E�#rҚɑ3��gFN�dV�&NEQdiQd��5�E��FZ*ʭ�rAidf�U�Atdrц�����r�\<�)ڴ�����uE��+�ETF��Y�KD��H��Y@tr%.F�����IkTF��Â(^%��P�:�"�F
���EbWJ*-b$Xm�N�#hY^].����`[֔{7*����Ŭ��5��2�
E9�D�xb�Kx)Q? �`=I3�IZ`�M?Q�$PL$-��#��Rb�vL�(�w�:�#HZ�� �csD�fS�f}���;�#I�$i����C�j��tO"i�҂��7c���vG��Y҂Y�oQ�Ǵ��xI3K��o]��M��@��ǇwL�t�j�[B�sB�:Ӧo4'�$k�Rr������u�M?^#�Z��)�U
�
ZWm�{I2'�s댻��{��Q��� �u�g� ~f ����|t0�՝�W�W���|ǁ�z�9�#%����������\^йjon-���@�}�:Yb�H8�{md{���]bZ������-�:)�_���U_Ef���%����NK?W��Fx�D�%d%����$m�SPP��rTܥ�J8��k�bw
�ɈIء�FM��ピ�"-���J��5����	�S>�(�)GI��ت�	���yi�rW��u,�u.w�V%,~�($x&W%|^�ݍ�v���{�w&soib�r#x5NatI�\:�����1�,�ȎwM��,���l����� �;�"i����T���F���r�54��4��<^�h��V8�e"���W-���6��'I�x�$'AM�@LRx�Ί���S���)ƀ��ˑ�^���c�C�a�3��"�ů�b��q��(���р��g�;(��qC�q�����˞�v�6�@�K£$���Je�4���(����Nr��T�	G�ĳ]�'<��Q<�C�֝�����'�=Zr�ϛ��.]�r�������(�[��12���.�2�P�0��Q������)G��|A�Zx"�U�%m(y0���)��
��4uv��Z�����zҢ�7���|��l$˛�_����S�xn�V*��u�z������8���a�=�C����A�C��$m�{�%�/�	�7T:�6��FrH��x�ZI��������9��9���4��5���??	s�1��Mf�9$�'����`NĝF��͝��@���I:F���d��{j5u�I��IZ��B@b��Ky��^��a��S���xzvȓ(z̗k���	L�4��Wn�Y�j$� ��͜e^����5�Q�g���@�D�!���@���a�����D	�48f~�+#1�ш?hv���)��y��K�xiv�1ۨ}Ԥ��N1mƷ����Z�m����A��T�j��Ę�W��M~�Ó� �.���H�C��1�g�����J�'ߘL1$Z�ø'i��(��1�@�L�����W>���X�/-�qR�t���oL5Pc\ir�F�9�5R�^�;����l}?շ�2Z8T���,�{@��ۃB��N��h|r 8^>
�U�EKtE�4����eK7.8u�չ�{��:�y'[)�x����3�γ
扺2u�I�)�2~�B��&�����U-��1t!��F-33�`���~O��&j�����,�Y6h(Sy4���m�nZa(GJ�����>����(�Q�g�_�٫�I](��v�Q���tKO}�T��s<U@�Y�SM;c+K�:a��	��0k���B@�s�ƅ,��p���åLԨ\nj��'��j�I��q�e�l:)ɰC'���~֎���$��=?0���3`d������d��o(	�?�%��C�8tn��}�ܸj;�չ�S�g�L�g�jڥ�9R���ɱ�8-ɢ�~�}b�^�LOj��f���ˮ`q$��~iEl��%���z}c���
C"���|R}��F�܋���Z��o�!��R�|
ި����mSa�#����ШT}��'�a��iF�Vjk��:r�ߘԏ~A����4���j����5��Vg������dB�����Ѩ��dĵV<���q�T�XY:*��K�b;R:.�K.�_�C��uH�h�E��ˤc1�ɭb�rG�����P+�Z�˂N�ԧ�T�.%s�؈4�����������	��C��Yc܁l�F��aq�V��j��թ ���WB%�����׺�����_Q��8Z��'���9u��w��I��SxIQ��a-B8̾���؝��=Ҫ~���Hc�e��Q�RL,�Q�1U-��hmV��J��_}����t�Fa?����E�&����2���%]���2�n�$3�i^�cͷ8�;�S5q�Ov�^����C;;���iO|?X�RմZ����Wږ����F!��!X�Kϐ�T/��:Y�i�Q&��ǔ;�5Z���8�������b��^�c�s[m��5�߱Y'm��>Ve��9 ��T�?T,����Ҵ��g�o�B��ZU�F'Y�|��2���O|����ԁb��ì�3ӑ��g��{��5;�u��T_Cb�a���/~>\t�7�IA_:����J�H+��$�\�J�#N��Gl�X'��X�!�!#P9�[*L^�>�B*y�ir�!�."�~f���Hi1�'�lz����7lM��)�Ó����N�$j��I�qb$��$��A'E�f�����3u�mRk��_�s�w�?����Ħ�R�xE#v(u�8Zn��p��y��Ҳ�[���e�[���e�[�E�2�e��l���Fb�C�.�e�*��3�<�jU�ߓ��C��X,BN�,
�M�3�֛�Q�x\�z�<RyĽ��D���=��6�\ȄA���6����!�z�q�4ŷn4��z����;�Z9
�b��]%� '֟˰�%߂���7u��A�zS7��0����z�@�������	إY��=��m�,#WI[�"����0-�k;ߐ��<��2��9]=DI4E����m��h�4g8>;�i���"ٰu�]���E+A^о��\&��uJ)]ٱG�K.V����ĵ�|�x?��p�Γް󁋾x�䐂�.�xTLhø���1B2��ױHE0�@ub�����«g�xD4�>@7Si��y
P8ֳ?l|4l�GX�.>�	��3j�� bZ`?�ebb���j�6��"a�H%F)��'����5޼���J��X�Ke�P�R�	��ew�d��N=�	�;�\�ű�͑}�^0\�J��$�$Ğ=��h�e��2ʒўF��Uʼ
0�e���$}v�h��Q��M<|�c$���d)ݐ1�1k����!��F�eZ��ܻ��4���[�9��')��*�L|J��F 6���`}�B�k�P���6AJ��j�YNГ�jVd%�"�.͎��J��,��v��5Ք4�p���G�S�%u����}8g��S�i�XE��8۽��>����9%�9��@R�5<K�v�����9�`�ە�S��Q����6�/�A�0|8�a�,{�Fc?~�%��5��w�������6�Í'�<|�� �J^	�{T��KCp���s@��tE�R����'ѽ([No �٠d{��C�T�/$������.�"/�{ ��p�*M$k�#�A��J�S�r�3�mO��|��{QF{��Ѝ�h'L��mM�R�4�&с���w�]�W_���0��w��E+����4�{�tqȐy-���hd/�|�
Yr�k�w�j�h��f(r���B���� ��p 4�~�����#LN��ޮ\W�یON��r�_�6T��rb��\lq�d��ӧCT>�YMտ(Q[N�nXR�.(�P�q���G�t� ���)�0�����0�;<I%N�~�G���A7��leME�pG�0ۓ��'^~fъ��׊�i���>�ce�^+ŧU�2�ı2I����𼉵���z�T���%�7�)�=a#UM��'r"�z����1�7�Ȇ{�vU���+*o��
d��n�-���J���u��{*��*Ls���a@8l09`t$e�;��牴�_b;��z�[�m�>頕bS$ǽ&���Yf�5d�W>� gY�3�gN���	ԅ���m�{f�}�#�tͺ����;v���9�o��1U��o<`;�z���g���1���7�fM2s��sRR��a�'u5&]@7�I�Z��9���A�3u�+��b��D���ľ�~{��4��9�#��aV��`���o�����=����4�0̯�Crէ)��hF+��{���-� 	��H�c�@��ﭽ�Y�+�a6��pE���@G>�臦?�~��܇xʹ�nm�K�d��z���F?4�i�;���f �b˲ߧUH��=a��W#�er�9����l���4��ZI���p���z�xTi���vN+-��!�Q.�u���d�K<S.E��l���<ĄN\����0��x�����*�b:�^P��F��a�#�Q||�#1�>�S��(���9�e�.�;�v��6\�;~���ˮZVg-�a���u���,̰",R�2�a@��I� �׸�f���y�h@���"����7Pߧ��0�1{SL0���TѭG��LW��OcI�>��dы	�ԧ3�2���Q��V{���<j��|*r��U��.&�i� �VǇ�v�0�wX�e\�<ƪkc6w���_^,C�|!�$��ع��G��El�H�Wc7�U���\���t���G_0�%J|;�~_C��B�j�A�?�E��Dn�"����(ǫIfϺ&�W��B;����6<iSO�:�B���n��O6s�����x�L��}�1�'�c�#Y��X��1)���x��|�Qږ:f�w�vm�ײ�u�Gx�&`%���iO�MnU���X���r��R��J�;�Z��HԺ��Ӆ �y�Z	�} f�$%�\��y =�9�щN�q��
S��*^���8Ul��I;��':yOg,,���V���@���V�`����8�p�Gn����1��{@�$6��3�**l��2s�P:O)S���Z�Fv�������.�N1s�Jt��#�v(�#���$������Ӽ���t�O�3?/�P2���p������3�c�1o%=���}e w��7 ���v[��T%G񸠌��`��Zy� �m����x4"��\�A��[�qW�7�C�]�arՊ���d�[q(��Q��A���]�F�yP.�;�D�:7�1!����23{��tv�9-����0�5aױ
k���6�oE=�� ! ��
X�J�*>��ن�ODp��Ƥ���̠JfuK�Mp���ۺ�c���"�\�����PK��B� �L
��E~�Kz"�_�>�:�?�V�耩٦�Pi i�k?���3�K�aF @�3d0Z��4䫱{[��xRQҌ��4<[��]ǈN�a�+�cvzF�#5�8�T��j��T~�?��s�&D�	�����l���F���R͜�n���F8� :�15�0����*nK� �-W�b���%\�ő�f�ǜDi(�\�$k�6��cF������S�'��X��}FJ��g	��@�lVv�Җ� ]ڀ�E�@�O3���pm�k�|��,tf�w%�nrR�j���6<���4�O���ܘ���݋�I����[����R}��(���%�m���v�%!�u�ǄQ@0���h�ا����b�q�rAQYSa���E��g� �|Im�qOo�v-�|���V�	�(��cc�=���@���� ���xkD�����e��X�ɻ�u�X"�?x׈��=LG�y��^ԑ���w�u̚��1[ j�8�S�f�0�a��;��	���Z'��Ve��{J9�ҡ��Za"�1q�m)K�xI"���Y�SO]�3��b=�J�Z'ܿS?;��D�3M3{��v�A�3M;{��6�nu�f�u�f�s��<&x�κ�{�`�w|��!�&2 ���/�7}�}��2K������p�-MK�	,֛�t��&�ۏl��X�U�37zO8³���)gjk��8���O|F�'>a�1�'>��ʒ�����z��R���4ֈt*ƴt��A���&6h��H��]P�kӄ�=E���(A��MB|�
��m�Iȡp�F�n�&�YEO4@7N���x����85mjs;o|*۝[�=� ����m[�i��ɧ<y7>fh�_|�{��:�@��L�'�K}C�B!��e]A���u������Ԧ�mˋ�i�(�X�S���d�W_��5̸�o&�tp��a���]k��Z`�H�EAT'��{�$&N���M�}F�}ޠ���>�)\��@,�)C܁��ar�%]j���2�'���9!��Q��\T4i����Vj�W���+�m���lIO��g�����|+Z��\W��㟽����݃�Ը[GZ���J�G��vdj���\>�6�$�k��|԰��(M.����qE��C��9�?�P��p\���]�eRcL��O���f�er�yG�g�[w�R���V�|wޓ��d��l�qպѦ�Ŵ۝[k����с�X�������L�3w��N�G�Q00x�R����o&�S�'���ښz3�+Hd揉\A"���	�����~P���v��r����k�,���{UkVsM~��U��3�bPs�Q�Eu���V���H������,7鱋�;W�/DҜyOҾ;i�����4w�75�ރ���ȯߝ��Wc�w��h��5�}z&�>������ ��f?|j6�d���q烐{�͏=��6��Um�g�6�k�,���O���w�=4����׾=xhl��%�Wk���y5�?��}���6�6Fv���'�r�5���m�{�z������?��k��K�?m������	�)�-��E�߾�~���7k͟��2��M�Gͯ����}�����O�������s�2���S^�;,�����;�$F7�9�����ħO]��5϶��'=uoɊ���������K�ﭩ��|$�������M������~��jr�+����T����^���_8����_8���޸��gC���WG�}=u��V�ۆ�����˸�����m�W+>^O~�\���^�tf��
H>i�k�t��Ѿ�w����_V����ȝڌ���e��������~�	W��_�e���v��_]����~S3�ԣG_�|!�����_�q>���L��I�]���u�X���.L�z��>ܿ�F{)�~����C�� ��H�g!�1����k-�4?�������箛��]��G-A����������C���[0�&����DD��V��VШ�[�'�Ot���y�֫9���.9ʏ� o�+!S���q��%�M������{�[�W���,ArI��J�q�׹��/�5O<����E:C�	!�&�,o���'c=��}&�_N�EO*M�g��'¥��k�|��z���r?�y�lh�8)@N��Imॸ�69ڏ�N퓭�WЧ��鍊 �G�:�r�r��4�i��NN�a,��a���q�ĶK+��q	��4<�]9%p��;:F�$5o����x�q���N8��{���INDAV����A�!p��z�3/�H:�L|Vo���QΏE��@�����vXP�_�ZJ���Cu>�����-�LƩ����o.u{eF���&=�\dF|�-�T���y��T����mzRa�_o��N��Ɂ���:_��M6�r��K��9��hr�4BP:ϸ{��^t�/�Ҡ�@� q��y�1�1�|J� <�Eڻ4L�������n�oW�a�=�t�Q{��!(����+W��D�y����%�pr#��
Z��<��{����S���齔��0�U>~(/���j����ɱ���a���笄���W@S�����*��*��]h��s�Ԟ(Ɠ&`�q�)�q��:�\N�Ȭ�&�����oq$i|(��Җ�-Ρ�:}��Nh���{�.�6�[���� �0)�m|����%�����$Dsh��{&�c���c�p��˸��\���g���1�=�*���B1=^u���2��Iծ��	0�39����x��?�@���"ڂ�1�1�|�6���������|�e��q�}��qy���K�
����d_-H� ��
���SBL�R�%F�-��s�xd��7|���3��ǳj۱��������ܽ����~��gFzf͑-:��sı(�TH�H����ƹ��9?�5JA���]�3x�5����!D�V��f��F�ɏ�$bR2���i:;=�=�]<|���<��s�����3�]����?>$?��\M�sЮo׸,XW��u���,�`X���^�e��{mb�~�&>a���$�!JOw���S�%&�� 	��+!�x{�*͆P�a�w\�6D���FY,Y���Br��Y%�w���hQ*y�tNxa�L�~��s3ئ���8�`������s�ztb�����ϳ:�1�8���X��}-��l�xa����<D�-5�n�(���2�Q|������0(ճN�D��p��_ގ���ۏk������x_�dEȢ(�:����B�d<��J����0Y��H�g�%]��m�k��+u���4�'ڗeU5n�Va����� ����z1�ׂߟ�,����� �J8K��g�2��,�5I����'��*~�r=Y�7��_D��'[�f�Yw&�%y �-T���\�� t���p���}�n��zPJUJ�&%[��^0G���n�.�I���g����+I�L�C��	����K�FsY��L�͉���E� �[��bk�mN�[u�qH�
2ns:b��8y���1�:&�i����c�cr����;�X�>hp\rp��}㰜Īy?�I��Ⱥ^�'e��M��y���[�C�3��&Cvq�r4;��ҝ��mK�L�=�&���'?�L��o��ܼ�?<F�aP�H�����!"���0�Ov�W�v��D~�
u+�D�펤�"eo�@�8{۰��P/?+{YtC��*	(��0g���\����pe�IYoP����]�D[2d�׊"��炝ё��t��ԩ�G+wQK�c�h�=�������&Hb�K4���չ>�$��=݊"H/-�p
�)��I�]����nAH/oś��0jj���])?t��s�%2)��Jk��c�
���&<�q��S�	Ocf��l�NaŴ'Q�	i���~?S��DY[q���Hx1C��i�D��i��4!�3{�u|�W�������<��j�L���g®Þ��y̮c���y�v�yBv���:���u��ݥw;I�A�𜢬�繛l��ᴪ/F�G.�i��"�����pJ��LX5`�V���
�N�"��&����ˌ�E�9�4����01���lE#��8�8=\
�rk\�-�̧t� ����Q>�V�b}�4��co�c��0P���� �E�+�����~� S����kv�C�L2���7�r������mcJ�L����	��/��ۿ�F�p��
� ����y�]�����\���rȬ�v<�Z��k)�ڶq�[�lKb�j+���s���m����c[�����h�C�2s�~8
Q�{�u��$��ؑD���xtsώ߼�������lQ�q�l]/dr��Q5g9���@��=�9�^5Rc�{fGZ�cL��my�(o7��x�8/M��A䶩�J(�Ϯ����ů�{}��e9dN�C���AFjN�%x�0_�/ʷC'=�?�]���`Xj;�j5�'p��@E����1���x~���d�m��Ë�����RUm���@�@R�B�N�=���S\��h�]�=k>�������e���n$�#Hy��q��1�<��~���W�8���F{�F;��hTjӫ�C�e��Ik������ń�5�D��]`e��Ճ�����~����b��÷�H[<�3�I���;�U��6�6����&��ɫi)�}�=X|�޵���Qz�	<�<C��0��
���01!�`��E �g�'[��pH䙰���%����%x?�H��X��|���Dk8ʠ=�o�U�cU�;�&XƑF��� ��L�f���Bn{����Mo��k��M�dFa��Xg=^7��lcĄ���O̼��-r:�Ց.rM$7�ǩ�w�:��}cW�3~�k���b��?���k�}󷘺�}� �#�[~��8�%���cu>���G�O�+G��	� o�U�ܣ�ɰ&�eA����A��oܓ�Mߧ��s3HZ���0��w)�}O"G�7�p�K�ݒmI��~��y#�"��%^ɷ6&ko�G�4�K��Fs.��f�?k_:`�,��Fs��w��<���7��gܓ���oA]�a4�B��y
W	�s\,�є� �r�M*�O�C���>������T9!.ZY���$+�`�1Sv�5j$��|����|��?Z���{(��@�ǈI�`�����A�:z/�I����qZ!�i�H����>|u����-��9qk�=��w`�=9x�`�C&)}���,��3�)kz���L�����M�m��� �'q5e�U�� ݗԥ!���O��c���;2f	�f/���h���t��X�{���D�5r�;�w_�i�� !�F�7/���?��{Ή�Z���nu����;���T|��Ȃ~�;����W�H~��]�;�E+ߡ7?'?���l���;,1ͳ��{򞆼�!�N��l6�MnbxA�җ�浹���7)�q{�f���"�1�Y��j�p���*�� �':i�u&�$��15IC51w�� �_.�`_ܯ�{
n�}��t��؏l{�耣��	�/�N�M����s����KOƋ��4�H�~��(��)���xKY'��o ����eP�X�՞{���d�t^���wi&�*0�=H�{��v�P5�~J��}c�t F�Fca����Jp��4�*>ѣ�J`X��gq}H�p��N0ݖ��i��灶,��B�]��߃��2rŻ�ۋ�K>��y�V�cSpW��Y�IO�`�D;�yA� �Y^N/�������7�?��n��� �p�`�Ɲ2ra��bL�x	�Xs�;q��3�-�g����/�E�ťg������Z�T++�=�8�p'z�����ƚ��W-���u�,�@��-��GY|O5��C�~3z ��TM��q[�͡�B��!2uއ@9C}�}[��Z�H>�Ӂ)O�c���ʗ�Ъ$@������jŭx[�j�^�J��>ø��_bo6�Ƞ ��9�}։7�9_�!i���Qw�[��*���!�;�K��6�qς�'!2p���g�;Eacλ 4��b	j5� }}�U�g"ұ��֖tP�,����r�F��>��<^�!����] � Kx��L��b�~�2����|�x�k%!Vr�0��8=�)%�H�	�1��dջb���u��n��U�zī��|�O���[�䨽{<A��K� �=Y��ѵ��g������e��C�����No6�"�E��AB����]@��4�I=L��ct2�ρ���������^�>�R�8Z��ݭQ=�qԣ���>o���|ϱ��O<���OFzi�����o�ey�9�ko�<��������x���u���5�k�W��i}��T��ޛT�>� ����j�W��	�T��`tr@`W>�V�����ʐΰK.����^�j�t.W��̒�o�^��æ�m����v�Lw�TA!A=�x�폺�9�@�o}b�q�%��|vD]�O�D?H�w����X�!J�w��l����K0xH�N���1��.�^�]c�7o�ާ�e��㫮��$�5$�Nv�<���K|�v-q���gp�\W�	���� n�o�ŷ�"�v��R9�1���?Cԅ�r�P�ݏ��,l�cA�E��Z2� �u
��%'���N�O��@�\��%�Y?E�Y?݂�#��k#���9�����;�1����cnA� � ����t
>v�;kqmۍb��p�}�9�;$�Z�ǁ�@��.�(Օ�C�D��fFɻ��ۡ�̌�����IN��jo=�tږC[:���Ȓ~2���U`��#X�.�~r'���	kk��sD&�^��䤫�gTj��=���+%����8G��F�k��M��X�!�^���Ӯ��r�TX��J�,H�n�C����*��H�	t���+���������p��$��R���2��|F������&�<�v��4��o=��*� &:�z� �
�^��JWau��>�~�z�.�{3�s��u��)��WԿʰHGc�;#�^���>��RI~����z'�]x����RW��f����<��g1|�>1Q�n�~aݳW�OF��.�<�BB����F;�Wwئ�Q�ށ.��9E&���J[e�֯u,��e'�"����t���]@4��oZe��,ɾ ���9���݅��)�]�`��`Q��)KQ����2�J��5^���E�^�d��B�2��_�o��4����$�4��Bmb��2��z�#�q-��J8e�5��ãd| ��
��pHQ��Q�����CN�7-��}�}Z��w����{zS���힀��.01m�����CA�oʵ�^�ܠ7ȃ��(�p޺W��8��pr��=9,�/��	�Q(�2�<}V��Sx��mߠy�^4�_^�<s��h1�X$�1����͖���̰+ۦ/!-S��r��,�b"GxŔF���úfY�'��qC���/�7����İ@>}e "���!�o֓��ؓw�f�>��fA|�5��d�|;%Rc;���C����Fw��?3_��l�ƹ>�D�ȿ:�oQ��-ɂ���q���c4�`1޼�t��a�t��2���U�,�_�r��H+�S;�u�H\�C�O ����ϫW	��|>�k�ȗ�&���(E��Хޟ�߱��W�}�0^��%n��Ȑ�.��8��{��g��w��]�=t�}�w��S�O�nШC��_
^�/6n�Ʊ��h�;W5`ba3����?G������������"{����'-3�i�׸.a�&�;r�[���H��O��T�O�7}�'����ɶ�OJ�Ʒ�Q�i�����/%������<�'� 3�6�?�����6=��}�h��~|#���tj?�*):1͙;hpIv�AdK�?�[A�i#a�Ɠ����߰5�§9�7��ј#;�w�hb��	���Is�	�	����9�BȜ0!h�;q�y��7Ŗn��H��B^Z��D�i���<3���I�� �M�b��,��O��'AW�n�Wz¡��H��
Us���ݾ�Hmj�"&���n�23�]&9Xt�W`"�2��{
���Y}M��V@_��	1����1k^�4�^H��`�W4R�� 9�<��x�J: �������~�:1o��o��F(y3eR��~���=�o%�����رLb�)H��=�9I��ڤK�K ���R�K�Nm��5�UK���	^�E�2�.��T�s�\�c�>����8��>��ƚ` �N���AТ�Ҝ���������$̮�,�W]	������+ÄuUW@�5x�x��<̀x_��.-=��	�Gk��D��Ћ�n�����U�g+�/z�
�
�ڋ�'��1�0�!T�fR �y�s=���t���j��H�5N���<�R+�R��t� ��/6�{A�y � Gx��K~�I�����&�Q�;�>�,B��B��C�l�"y�+��xE��H�茓�r�L���~����8�\��`p���5�ق�B�S�Il0!�$�7N��d��*yy.�����d�j(����^�j�<�n�,�N��]l��3���s,�����p�A�������V��r�?f>ٮP�� ��?Qhꍊ���qsa�AS�0��˫�s�ltDVD��EQ��6}����va��)}a F��i�l=��E뱸�*�7�q�*�&�����7��@��^�9⹌�ŏi��{�Z�M8F�9 x�Ơ���׷#[�=�����6�ϰ���#��'��0iP�${R�R�A�j�lĭzζ�j��	zk# O㒪�ҟ��ȱ)G�[�6����������m!���V~�#��lo�~��, ��&����,�k |fŦ'�详$*lIω"-����#+�$7�k���(8A��H��#�Vu/S�O�m��TG��o���S��0>�oI�4�t��icJ7�n^��>i�[��<\����Uܲ�F��]C�w?��x�� Q3�3�'qs��Sl�yok~/ڋE���?� ��=Y�n�,�tC���Ut��� k���r5��Az�'	}���b����H��
[�d�c��m+������9��5�4��7�(��Nt�X���W �_1\t~M3a�5�=ߋ�=!4}��O�e������U��h�$T��HA��3u�=��Wx��E������:y5<+��륔.)�{^l�{T�����N�:�������`H�7X��{�A֌��|
 p1z+I��C�
��e������͔퓙�!u�y�܀��_݂����Џ���ԇ���@��szt�W��S�4KR���UE��)�%.�t�{0�="�|>��j������p��/�!�ӣ{�:b�w��(i���:��va����h�?ӷ��9�Iz��M.I)}de�h�]�>���]�<�����n�s4��bR.�ۅ`ܚ����xx��T���4�V�>G,���d���ػ�IR:իħ���!'��N�N�6�/ �����'�<�����xG�EO���}NWO_�r�����q�dw�[>W���R�tt�q���R��Uު���@��-#	J�jk#�K��ka��Cr3,���d1`.>G���zz�_�
�5��d��%��[Ǧd_��R���rA��zЄi��6]L�����ve˄y���;�)]^$ �/�-x3�k��k�߾p��G��*���V�egO]��>����y(Y�(��E��
8�S!�e���!P�#8�Qr�R��B,�%�O�s��\ɴ��3��OzV��J�&>a�lS�����$����_���oi��|�B�WAl�P$%�H���3��9�����#�_�A�z�/����_�X�GO�����i�����iY˦�wZA� )���rZJ�j���������d�ԲG���s£Ӓ�(�����
6O[T �M���q65��ue�/�
߈	)�Xk��TPV9-i.�0�%�8�g�+��/-_3��̗/�Z���,\%-Qy�Ty++���!/��NR&��V>2-9e*$S�+���2/o�eЉ%�'Vx6�c��>>�M-�P�H[x���mJۆ��y7�Y���dje��x�M4�dM&�e��)�޾��F��WF����zj�TV9-u>�U����ee��l(MZ��-N�c�8��l����W
����[E��!����K?����:����/�\q?|ɣ�7������PX�D��h�$Kf�J��%���닠���+��+�

-EV�?
��/*({�V�h����qE\Wߥ\,7���B�Na.�?��� ����+h���0����;���771)9%�ӽF����cΗ~��e��堽��4[��$r��t��K����hl�o�2�`+�G��IGن�����6��{�����������K7�������wH0��~c�`ML�]r��N�S���F����*�~��G\��p^�A������&A}����Yx�>�{�]����Ϣ=��lo�zu���K�Q�~7�`>͞e��.^K��Ne�Q����!�Yr��mH���7��6*�����W m���y�\Ef�'s~��.���[�+搕ݺ�V�5~旈X�G�-���}���$�����J��y+�s~P�r?4#���ׁb�w�䱿f��3�d;��#��<�S�r��(
�^� %���n 8������?��I��.B���9�/S��ާ-~�"<������3r�7�v�7�j���|��dtLV]"���ô����=.��?5��mÍ{"��cl�[.b�v��g���ͤ�헦��b��
3KpV[Jf)#�t��C��)���kW�9��_h�xλq㦌@#b�oV���L�nr|�#�<9`O�{���'���E��U���;�E�(kѳ�}amL����)�b�őr�R�+#Ѐ�4�W�������v�;�^�$��*���s�|�T|�4�7������w���_��;��l������O鳅���{2)�2޻ ٘��u[J��
P{�]�n��w1�d��M���^-`F�W/��G#o�$��C�M�J���l7�b�X��`��f�/�ɉ/S�Ի$�K��2��lv����/ccm�$�Sm����R�G��K�'{���s���o�?��$�c1��zg�R���/y�>q�,��`F�<�s�v�wk��s�ͣϔ�_D���Z�B�U���v���7�Ψǰ��&V�g�^�Y��ܓ�s��E�`̏{��_����0���v��)}�A@��Π?��og�����&�
�=��E'//�����5QH7U+��3#�?���<95ee��u�Q_��v�&�?@�� �^�CE�qJCk`�p:�9�6>C�Ł�%�Q��]�yŋh�^��G��^�(�Gf�<�"�|/V����Y+�WYkVb��^Lq�YT�����ȞAt���Y�Fzi��1
�kC���T/|��������f)��;[�yטsx��w��}�-���z��n��P��kd����вgb-�I�Z*O|W���٣j��� �.������:�>Q�<��`�~T���k��R����}u�d��6�J?��F��{��G��}ȼ|��-��F�h~�'i}[,�<�8�}��o�u��h�`��O� <�C��Y�ܽH�i׏� }�'�}<����m���]t�-r�/��: ͞���>�lD-^Zt_mF�]�2�r��	�F� �J��KH!���a+�E Y�R�T޲N"@*�� f[�-j�7u��<]�skoIA��2���.��+��giq?s~���߮N�K�]����0���S:��x�ޣs��R���|�E�W��P����~�!�ß>���b.ݔ��� �G�ۛ@�hd���}م}q�w�����
c��x���v��"�{��H�o�S�v3}��)��~��yC�5�n���鯢.$�<:ѥEs/���F���U��j�[��)��M��2��|�v��:�����{<g�40���;�dskfv�8���S�������q{��� ����?�}\�U��w�����B���Y"V*h ���>C#a|�h�%
}a���l�[m�[۶�n�&��#C�i�h�⃔m/ɨ��Ϲ��03���������s�=��s�=�yp�j ����ɒ��3�ĩ��9��yw��Z����?���g�o#��-؜�i��"%�W��W|]���[�~�}[��C�_ �\�8��_Qqa�d(Cqb��Z����Di �?���s{@bx1&����f��|���cנ��]C��ʨeKc����}�� ��3�R|#��́�IV� �������P�`�uӠL��E���(.}}ō�Ib;���G�fYd�$�ޣ5�܂�_O�Q�N�4�}�K�
�w�^��5���*\V��yT>:�cg�5��2�{yX��S�?l�Sñ�9�<[���s���'�g�S�[�����t�6����WC�y�b�����5[r4��,	��ɝ��Y�BKB4F�)��Yi��xӶx��t�Q�*�3]�>P�|� p��j6%�
h���E�����,�1��Y�c~1@�K�ĩ���(��^��#�����o�}�6�g���dv���!�j�q<l�dk���X���ګ.+�v^\�a��3��lY�;<y��Ɋ�@/p5�B��OHʟ]���r��Cfkr�� �P����<r������+?G#��ʙZ����t�[!�*�qBѼ�J��ε����:K�֠�4�5�(���\�
�:�H�9ln_��0�7U�P���˝����Lם�m�zUf�#z�:Զ)1�`�"Yr��npڰ��+�*g��۝�����tޮ��g�~����w�I��yM�� �� ����i�WV=6��3��{�ғӚ�7J�:qBL��N��6c1:���/����@��&\{���*�����t�3��k�S�F�O�)v�v�u%�Zw�k��o��д�~F�|��ګ�o#���3�׆�t���:�w8�֣�d�R�!ѝ|;u��w�7���(V�Ɓj�o:�<o���}/5B�w�y�O��%r�뭗Æ�++o�X���w_�1��_���џ�݄O���1�-�$)��4#y
��Rk�2ں��MW�WY�z��l�<�J�ʻ�Va$5��Շ�W�
K\�(�bx0�}���.*h���ώ�( bq�3��Z:��C����f�'ێ��U8���Z���wv.���R�ؼ���� ��q�}�����sR������0Y�{ ��8��߱LU m�/�:�?'�Or���r�����2N|�$���ޠ�u�7���J�i�@���TBI$Z0�����	�Ϫ�X�0j�ý�!�d�D�5����*�j2'���g�j���^7��;�6u��3dI��'UEҾ�A��-��B4Xp�%�隟��?x[ի�/�;�l�5PM�P��Hn�7��p�(�����ߠ��}�nw���.%K�EG��4K5K�����I7�^���[Ɍ߀�U��֘}��< �|��A
��w���P�O�� �fy��S��뵥VP������1�ή�.`��h�+]Ϊ�X~|�ɤW��9ب48M�trn�����07q������Lc
�{!p���IU�(���H���5�o;iD5��H@5�N@�eά����ig���*-$HO�ӕ`��@�*)�J��H��R��0g6�s����&{/Y�W�AtiM�NiI���`z8_��26�~���Pf���UT"9^�%�v�R�Âr�ΐ�L�����ULh�0b���+@��84�1��z,�ߕ`s�Boj_�)Q i�"�׀�1�\E]�<_cL'_"�|C�,�E&�t��iJ����I��pA�M'�L�=��#f��˘�p��鳨�l_���_Y�����Ė�g8MM���%��0M$�KzȦ�gQ��l�d��ln�l�-��q�X7��̙��sa�%�v�R?N��֗Y iP�Kk�q�\��׃�!�O�f�
	�s���M��Dl��&������ �x�(��p'��+�3ɜ:m��
)I�G�P��g�8��Usp��#58âz�9'�ۚ:s���`06F�̵����h����a�_=� ��
��l��N����/}%x#/�~���g�3���u��V�4�?�����5?:�ݑ�l���v��C�a�hf�!��cr�59��4�q��*.`�z�J�A�F�i�cv�Z�6�4��҃S����S��æ�r��8[*���ѳ�7��#*l�b�f�}84�*�0o����e�ƽ�!���㍱7���H��ct0 LI,	�74 	0�����}�DA1P+���2�?r���O^ᰝC�W9���u;8��a'�N9���^䰉�s����p���%��p�-��q�=��㰎�����KOr������4����,��8<ϡ�ÃVrh㰊�O8�氆�C��S�px���8���/8����~��Nwq�!��9,簂�=��p�q�1��9<���n�������÷8�;�os���p;��r�O���{�q�{_��n�p�D�V��/Ȑ��@���kS�[����^RS�3�f̘���jtcފc�~I˖�=��j�0�9`�1�	�K�%����.�����wL�l��������i�	JI=�q��Y�0#%#%!>uA�>!#e����I��#\t�=��������+sD�UR'$Y�?!?7[\�?){�S��sS�rr� .�u>T(d�[j�_�0�� u�§
�WJ��b���|KXa���Xd+���<��{�_eQ����\d������=�/̕3��i��ご9)y�Jak('=	��#%:dF�BS~AHބ��N[��$o�����`�&=wy���+�Bwn43rr�W�� �e���$���3R��^��p�@p������܌%�y\�֐���K-��|�B�
u�c�9��Fvm��Rw�~-��D�8��p,�c8���p�a���q؏�P�j8Ts(p����6��a���&9<�a=�'8���(��8�����GVP� �53������e8��x;8|�÷9|���9����n氌�Mn䰄�"�}��Gt�9K*jI��t�<9HBM��gҁ�e�\�qv�D�>z��4�$���q��6�Z�ь]��@�,s^�i9\��2s���>��l384p��a2���q��X�p8���0���9���j8Ts(p��u?��U-h�K�����t��ps�a�A���7Bً�~�R\��TN��6�mO҄�Mt�~B�|���o�����9|��?q�*�[9�3���5�8,��9%K8,��7��Í�9|�C��MZ8|���q��ç9�簀C�C��8\���r�@��~�
������*�֕[' ������[t�I-ӤH26�{�H����ڃ�4rp*����M�lVK_�T��`w�u��mN�[J$��C�x���Mmg��ƌ�^�o3JG"��}f���l�@����3\������+qxW�<=�s����d�]�8�8��� ~;
$�f� �s��s6:�yx���4i��wȷɟ�4fJ�%�͔|���5�毡����Ue�g���&�i�		B�/�2�w��*���S�3�xvϚ��6ᡟ��8Ol���:�\I�$�����Hv�UG�2%sp�0��c�A��gw���׊Oǝ[�Tڰ~�T�&ٜǾQ�<vQq�,Fj�C��7�S!Dx$�	��K#&K����HM�P����\����#��F��ڰ�N�̛e�A�1~;M��z���S	��r����G+M��:;
u�����o��T�Yw�ޑY��TV�	S�F���~�HO��}x.�|YQ{����ش#N��1i����k�_oxv�f��� S\��`���* �_�A�fa�JT�@gY��S�=O�oHh�����nh��7V/u�푴,{Q�Rص��G:���B�KA
u{������$�N5-27ߐ���<W��/`�Փ��á���<��M.=*��c�̕*�Z�:�ɥ�xr}(�8W>��;N���>}g�P�/NH�'�i��Fe�;<�̆'���qB<����V���'�Ƃ�ڇq���u9h�� �ً��n�R����l%�mנN��n�1]RJ^^n�;������.���4V���ⶤ��O����v�22���8��'9쿋�!�p��í~����ϡ	`�[N&������f0�MW�P�P��O��*.~Jf����eF(7d�RP�,�B�B�@$i�8VH}����Mb��V
~)9�yT�~Q��{1�0��|��A�1x_Ax$^к�%}�;Ni��Bs�"f�h�-�ȥB�%J(ߕY�;��=Cpt�A��HÇ7Ke��f�/��G��,�ۅǡ��z�1n��zp��V����1�ZW�(|�&���.tr�8)� �-W*Z�z����Y�������[�ǡ�BP(X"�;#{IA�4��Q�|�R��FćQ��տ�۠��:�MT�]��n�q���`72[y�����<��Jh桩�t�E�W�����&��8�����Qx�1rv�-Ļ��-�S�-� ��!F2p�{TA�5����!�@w��R�Վ����N�[�
�> `�����v<56�
��X֎nyo�lي�I���l�ǈ
l�:�!����n��1i/%�@��[��U�+�di�	��b��Q��+�����Mx�7��oy��A\��r���_�a�^�H˄ue��xӲ�K<ܶ����÷_u��r��<���+�R�K��TR���tC�zd�l�כ����`��ݨ!�ݵ�@�~�y�ˀvL?�����������8�g��ot�q�ষ���iY��g���C׻>�[��::��Y!�V�;���!y���=�#FS���� }�U�����_Q�qx8`�o��WV:�}��J�z�gd�-ʥ���<�7#L���؛�����]Z,�i�r���0� /G��G���|h���������W�>-[\L9T�qx8`�7��M>t���y?�k���+])y���-ə���MF�������t��|�8����G)q_���qx:`�=&[?���wկ�+P�%يqt9|t3�Vo�|϶��2���a4�a����ʐ�С>���j�uz��%J�K@���|��Uٺч�7}���1��ڧj]�$d���?��)��,����%��{D寣-XJ3��O������������}��׵e������6sɊetuJ���R�c�V�c�i���2ۯmo��V,�]�[�qx8`�7ko;|����VW�:�B�t��j3�0� ǎ[зՇ�]>�o�J�Q�`��,A�b�]�t�d��ě�T�ﱟ�ں03;I�[?�������QZZ|�O�J�@�
�F��e6HW�������H,[Y�M�&��5տ��}��"����0� G��f���ozF�|���Z�@E3b{����|���ѷÇ�&���p����h���ą�OK�r����w܌�'y�[���Я�g}z�1wa�2�1�Ѓ�r3�j{���z��ѩѧ��["ұ6��v��{��V�>�or�v��h��"�Z��$[1���=����=���7m+}���:Z��O]�	J7�\��wycZ�@@�z$��]����2�L�ݨl����sx�g�q���H�Я��mo�I��#t�)��i��ruq�.wa�S��҉`�
��H��[��P\�*�cOM��6J��.�gq���(s0Y�^�eq���9��IJJ�.X����2:�&e� '	m�W8��þ�	 g��(����Ӹ�Od�?Cjݓ�c�����i+s�V"�p�I����^�* �b�\�Փ�	���B�%,[Q��!�z�2��l5��'�k~���N4?�"���\���f4J���~{ގ΁4³�q��Ó����h)�����4�n=?���;&<��G�R�~'l��KN�k���si�"X.bxw��'}�KFμ�d�(�%#�ȁ������r�)�bf�����%��]θ8�M���D��rc��KD�����;60��o��"�_%.+�葔���5�:� e�����)����Ҿ`�,~����Vq���i�e���D�LPGYV��-\�M�3���	ڬnky
MX����O�ؽ:��4@����hI&{��� b�>/�h��|]��(�*:����b>�qy9.��c��(S��5(yo�$��<Y��kxa����Uz��B��HX������V�%��T�} �l@�c�m�(���c�V��-\��$o�1� G��f��.z֜�����gu�F�7m�:x:�7��r�R
ҁ�e���<���Ӳ� �ӡ��a�W@PT�	������lm{�	W�`Ug;��/L��u/p�}���8��+39�͡��'�<_��9'|
�1P�'�H��p���u���W��3O@��S*a�d�g�s�x���+L�s��R��wI߇A�j?�3E)�m�[A��Y0d��F7�O��s�B[�P��E�瘷�~���"d����ʜ��5�79J���
9���������
��l ��,���`Iy2^荫�&�17�+�(�)��y+�@�q�Xb�օ�c��Ҽ�#�ɺ�T���PD0h����1�VP�2(������0'����P�s�i�k��,K����tu��4M��b����i�-3LeC�ec���;�������X�E�»n�2��<�R�(�-�����
//���<_�{�c�إ�X�o&��J�잃v��.�=��C*"�bl�����3�;�M�]�],$w�Z���<�yq���%/�J���e�z���t��"��*y��pfy����j�0el��}��21�k�ף�t�����n��DW?'8����a�� ��6����Ug|B�1�1>'-��@���gD��YK�м�Q����%�zP@W_�jR�Q(�o�f
$�dzP ����lm��Ӊ�����.c�����qB��sw{�?���acV��𬄧�7�y���Z��T�p��T�{���%t�q�.)mRƊY(3|ש{l�K��+�&��@��
d���1�B�0��@����P����
�����I	�.��GI�6�Ywֳ���4��0zaq	�H�iƽB��3���tc�=!�\��L�y��`�
�nW=T�c�X�=WX��^��0��TPTYm�N�eX8Ͼ�p��sL��N�w2�y:^�g<��I���4��+=eX%�8�n�9&`{�1���Hz�K�0\7��8�%X�hJ7/8/�����[\�1x�0��xd3+3���濵�}��ݏ�g�����fx���:<O{�_-�>��/42�Ojd�/itUp��خr�����F�r�|�r�B�I9l�e9��O���\��B{U يe��i,&V�>���w��������%_�V���:�ru~��xR�ɀ'�ڧY�m���۾�Y�����ۣX��fd�-�s������[s���0����M�.#�VE�c>E���B��}���n�R��+.z�_���p�EV~��/�M������.?��t�����,���,����a��.���؀y�y��e�Cf�m���ʃ�B��?�Y�Ya4���e���ێ���t`̤5.}�3�����V��)���r_���/R��v;�Kj��tM�n��\�a,Ec�~�0�5�U9���ta.�%0��*m�d��AC��P�:�+s8�1����	h��uR�\Dx��X?T��'1�]�Jn��!���,P�VHS!TJ6�l�\n��+C~Q>x����}>��=��+�z�ǸZf������bL�X�s���<���#bo�G�t�A�� �=d�?]��ux�܎t���S����CC?����MwS��癿�{���C�C�\֜B�p�\��v��Aqjm��\�Е��=�v�<��(+fY[Z�+E;�h�d��Z��~pJV�T��oH��8�-�]�tQ5�Ԇ�c���B�xo�)]:��p;wNr;ǂ��:�zC/�7#��!XW�0�Kr�j��@������K�����'��h
���'u��ۀ�j�6=sfs�'�Z~�{��g���C��1����nV���IV|�G�U�z�>e\���?���Wrd��H�g6�$!]Ǐ��a�Zo�c��v�E��Б	��e� ���ͤ{ɽ�,����Ϛ���hoD���N����%?�X)c�ϝk�I삳u�g�\ۿ��>3������R_�Fbև���$���z��q'�D�!�\	a���޵.�T�%z��IKl�Y��]�u��ρw�]�]`xߩ�gb2+ ��i3,�!:�l��C���k�w�1���9�G ��N��;Y}��ˋ�9���K?��Y����<�C^�xΕ�W�m���e�߼�~�#/��1/1O�L^�Z��P��y��3���J�L�+b~\�BP��O���ca03�0�GNE��a% |�77˟?���w�F�:u�I���`�J.Un�]�T��Y��U�9����"���-�{������xqn�52.W�ww����NB'�F"���^z�4ڢo��!�j���i��[�KG1�@�� ����p�[����%�_)א7���"��KW��f4H5J��#t�I���w9H^6ls߰.R�����𪦮+٭*Ϩ~�Q���|큏�:��)����s�.x����@V�P#L��7�K	�ހ�Ӑ�F8�6��>��fm$���c�o�=���?5Yl��+�;�Uʏ�	�hY%E^[(f��p�H�~�^%�o麀?�@��t�U��H�]��/u%h�Z��0��� З뀹�/r���|����ʄ��FE���X�4(Ǿ��h*œ����|�E�^��R��j3D57�mk��+�N�=����=n��������r-����l��$L��(�Uҫ,��UL��I�z��Q�����@����@�A|���=���J�&��9yJ�MS~���8��H,�Ph�w.5>`Z�0�t���)k����џI�KSW��,U���R���������	ڴ���S��tk�n��i�'�>�cd�ԍ��=A�>cfT]�S�*G]��*��x[��ti�ܡ?�tU��؎QCO�Uգ���A(�k ���
��Ɗ��ќ�)}�����(U�7����Y`4c�M�f��6ű�'���]m4�gN1A��o�i�Fj	�:<#��$�ݓ˳I�:� t��V�c�`��@�P����9�.n���+ �s�*B�}��`��Ʊ�Mc(��x�P$��\�v�27��GJ�m	폃F�'��5I�#�h6��R��ԺH��Hc�6RНi�v�qEt?��8'RInX��q�_�9?"����AȀ]y~�yu䩃�)���g�e��(�8a� l� ^��:X���)8ujY$��>k;[y��Y�d]`ݚ;�}.�)�y��z�W��)��P��95��K��B��#�\}^�;>_��ؕ����Em��� 7]���'���Æ�:�^Cr�8�5,:[�J�"V)����=t(���0wqLf�N�j��������I���x�XRzwo0h�VC�}�<��v+Ui�}D�8�;A����������^�q�E�� o�f�\��_���<S큲�Ȓ(��/Py�RE~Sc�r��?��U�PS��E?�ˇ0��V����
V�������{_�`�!��]/�\3�|���g}�m
I�6C�q�0�z� _.��.*	o����Y��lc�I�O�
5c��
��dSO5�A[�ʺu"�kX2[��(Î��N�Ӱ��~��'��趨�)�2��-���\z3&�V)�wg2�d(�}�EU��J�Uo�9�|ڊ�B�A�Or=A栵��7�1�c�r2z5����C	s�{5�C�Z����o�ˏ����9
�d�����b�F���e�x��E��TA0>o��ʭ|�j���a�a&��nv�0^�~ҕ�U�����\t��(����'@����?��ls��]���*�f�^d�����2v�����U�ydk�xd5���y(��{��vݳZ􃇜��7*�S��Q�x�VT��ŭ�"��P-o0:��S]�.�� �?|����*�M��&��<�-�����z�+6�R� S�Z18Z5�B?�0�`�8��I����x/��]��Ԩ#QN@��'=�:{���?�4���B�&�p|�NL������4����Ti��w8�= `?e+m�l�@yr+#6r�L��Ȉ��@����ʍ��u_��j�jx �ۈԒO>�f>�+a�q]%�Jן{~)� ��]�zӿD�t�o�"�<���eϏ��L�����TP�C�������m�{@�^��-Cͤ0�ȕ��B*�ř�h�e�\-�W���{mZ�{IU!��a�?
��d��S�qԆ���oЦ�4�7S�Q�V� �V����*ut�]��K!��`C���3���{�m=l�p;�l"�:�1��՟ۖ?�5��Y@e������z���W�,~
��ȂNA%v�:��m�Sl�������R)��{ӝ�/�2���9)�^hW�Nv�{�|�B{J�75�5K��YQ��е��y����y��
��a��a-3x��|�O%����3�����4GN��
��|;e�������y�;}:}�
Τ�K��S�vo�Lg����i���$��P���$����!ƶ>�����P��Zර&U4���;G[A�f��x�%�c��L|���k_����Ĝ��]�����BB���Ӵf�y�����
���B����P�H�Ɠ�C���a�T�e����h� �g�l?-YRc�QƩ�fӕ��b`ɷ��,�J�~:q�N����0 C5�6�����ϣ�}У�["J����ɜ�؁�g6\���h
�<&
�5zSb��@)����H�$8��Ɓ����ȹ.>ΜU�����1�Ȃa0"ԕ�n��5���!�r���nx��c{�Z)�(�3�d���9� ���F��"É�׌��O�˧=>/G���*���g�k�1�(�p���j,�A��3��H�P9��}Ŏn�c�VPS�J��>�
]L�U�X'&�m毌QV�����ڏ���͟��w9�aU���e��|��Op1�1�e>�����M�,�;��(��<��dR{[ؘ'H�A|D�:�PS�\�����;_#��K����sGl~�s��v5R��惵�6$׫�4��|� mU�dU3]�ݔ��x�a�mM���S�ϡB�����
�����U~�akR�ejJJ�8~��@�O�j}��Ǩ6��oT����1]�
�G�	�Ce�?�!��P�b�vPSZ����l��"�J���N�6�uۻ�o����o�T�]�i���w0�ڜ�
\�*A9��u�B<�����M���}���S8����=���8�OZ����ӹש��,��շ؇�4�Gr����Y-�-9F߲a�=[���Ru˘�r�d����Mt��P}��mf��*j\=�I됏O!zFKj�KT#j!N���mق��SZ�]档�>bO��)�N��6@�5u~�+�Nr�e����zf��~)�D��@��/��}����lb����
���7<R�NSv��XprlR0k����t9x��DA��D�|��8��p<�+eR��S`�����Q=��q��JS���(+jZi��Ts�����Vh4z��\6��8a� �6n�b����w#Ϳ�~<[��E��(W�Y�8a�`����gp�g�x��˜�nV�?��YM���1Nx <���4 �9��l:3}��̹rV��#�(hC
/�4��i�Zq,��G��~{��a��~4n�r �9��L�DH �N��q�(!?�8a��z�SAƑ�h�6HZ5�nLu��fC'�tYڢu6(�p� ��?m��7�KwrV[L�f��i�ZƜ��u�g���[�V����V���W�4 <�����p��p+���@x�O���F����3C�kU�<�F�L�3�4��HQs��dڷN'��(�>[W�_A�+SW_��-�}h>"]Š4��π�-�'�W3��EW�u�hP��Jg���\��LMv��ǰL���U:s%ڵ�����վ �0C�ݚ��UK�{��~�s��	�?�U�$��yr�D=�Ί�:����<��ޏ��r��܎5Ǥ5�V��F��>�e��إ)�M3_ř��cЕ��F�q�My�xԜdw:�ve�`��	�Mݩ(����T]M��T]�*�*���+̈́v�+��\d6��\5��%���.����7%
�>�����H�>��*t�yfX(͗u����M�k_Z��#0 ���P^ѕT`�������{0���/;��6RP�gF]y��)����w4&uT�=(�������vM��kc��EC���dפGյ�&��U���7!%�j�6����s{^�N��=u�|�|>^v��M��q�:x�&��q�3���5x������Rx��/e�`�zGɡ,����e�e�:�
���T��Wa�nџ&��"v����G:7` e���D� Ǿ��J1��{��P���[Lg�,���G�:Pw@:F�]��)X�����nbc�q��F�<x��$��'E�*$�ϻ\�5ut����� �����6������Qu1i����7�E ���9W�v4V��Q�lo?�N�^�#h��Q�����/���ᣛ6�"�v�F�O<���(��Y�Q#$��,^P�S���}�p�&��j��w��:[���<=�\�K�I<m4ҵ>�~{��H9P�a���j@ދA�C�;UW~�x1�(i�)b��L?B�m�ъ���w��M@ս�pR�_Բh����&9܉���آ����������{t�/�=�J��`�l}��!�@ϫb�Ļ���F�A��8�t��G�k��$\8e�)�h���|[䰸��a����"�uH䰡q#�'r$�	n�"���ğHp��#1�����	C�{���*��F���d��C`b-�((�f����\��4�Is�`�[q��{��I�B��oy,^���UqQu�	*��3�lx`��QAXbM����8�b��@|�kl��D�ĩ��[�ճ�W^5���b��r��N�㼉X�U����>�8�?��D]Ԥ3����c��-:T���Q������B-ԾB���SpѺ�C���cT´5�� �i��o탌5	�(L��� RǑ�@�Q�Fy&�%6��3�Uӕ6h���&g;�����j���c��rp�[�~��^:-D�5��Be�Sr��:���	��^|z������)~�����Fsf����k�9�V����ۚ�x�����æ�� 3�O�xa��1Rg�bj���xH=�op@ )�Kf�%��j�� aZѣ��v���Av`]T���'�*n�PRU�J��+.+�����u�WO:^m�pjd�թ�H)�;��9\�+r�4)��?�u�U���x�u�&�,�����~�=�y>Vo
J�A[�يJ��zC�c�6�B�gR����J�I +��Tc�uAT�Ԯlx�����¶CaW����"-���gb���ۧ�0c��*НF������m���{>��*�{�}ޟb�$=U��,��5 ��)�Os�t��;��.�EGh=�诘����03	��E[�0v���e(�~-���B]y�4f(���|/�3Kut	Т/��]�Uju1�Ə'� ��~�_p` ��o��5��&���_��A���)k����	���W"FD6�T��N������!��P���<p>;�U���+G
>h�#�o��i�xO��3��C��#=�7����;�^���ؿv��z��	�;��cށK�:]y��GT���Y��^ni�Z4�c#_�=�uo^��w��O{�ݟ����$�{�����u�����#� �(]�-�l�����;��`<h�K�E�=�|ݒ�'.	��RW~lI6,�zRU	�f��Q���x�|z6�U\l�E��lv��ț����w��,����^�FmwA�gI�4�}���9S>�|�
$�Kf�Z��:�{���}��KX X��C��R���j�[W~J����/���Ji���l�S���?�6@:�A'�=�}q�	
Ug����)��О`��:�2�8� ��:��~�#���N����%�"�jW����e��c��I������R����U�O�O6����:S䃔�W�;����B��֭UI���ה���[僔�Wگ�Zu�6Uk�w��L�h�o �o�'t\y9�>ӜFЖ�fi\L>C�q���XzxC$�hv��
�������vp �q���7ŸO!_}�RX׷����V�`N��Z�߀�d����'���0��Im
2:Ӛ���o�}����)Ǩ���iM��o�{?�#1�q{��IeUY}��+Hx���+���&�jZ�t�+=����r��ԩ�F3Ɠ��1&�)��5��}g?/�9��;�V�Y�	��i^�J�@1^N�)��&h�:r5ي5�k����� �;hC����\�d_�j� �W0��H�*�=ߕ�هˎ�_�@+������1����A�Jc�<]�,Q&oG�:�x����|�f�\6CկO��-T��{Nejfȵ�S�4�n��������`��H
��.ۼ�:'_33,U�M����9��Z�Z�\���r��p���G�`�'��D�{���S��-r�]%	JY�+���1�]����|�S�i��4�eu�h�E�4��u��:W����$_�_C���L�쪎���
wA0E�����4x~�:9���<��犫�,=5l�f��:p�9�������:���4��<P��^;��;����e`�ޭ�|؋Q,���K�p����%�/�r���HW�K����D݃���P�Su��c|[�z��H����*��C���"���?-M�� 
�bYe�����׽{TV�'����PPmJ��t�b�#S��
�W�*}���"G y6*�m�[�R�-��O���r��%��\\6�/�$a����๞��������ʢ����*��g��R�:�tX; 0�A�8��
?�gu/�Y��J�?[�:�Z��KE��N5=(����Q��o��t��`+e�%˃?[��
�:��(��ʘ�ɓ���B��\����u����z��p��WRa��+1`��*@�Rg�ɾ�E:��o���� �y�y �ͅ���$��D�<��6Y�Bv=�S-,Ts�?��B��\u�Y�d�d}�(�~c�����?t�i�^��7&���}S!��F��$�9�1V��-�nw�������K p����_���c�I�^��O%(�����7qhp�!(����/���-x��36,^�7<-w����#�������o��<u�d�Xh!�d�%�{Rn�[DT�p������'� ��ُ2�����R�c��I��F���C�LK&4�M��9�-E~�"[2ÑO rcu8A�_E����ʐ��%��W�a�Q����=4��.;du�VA��4��>G���Ӈ&�g�A��d1%Y\nߐI�]D�`L��kP�Q�h[L�;���B�{8E���č���~r ���m+��~h'�y��m#����i�U#��W)G�AP�?'Ȧ�旨R7�� f�\A�����ו�K��}���G\(?q>H�bB"�b�Dą����s�i��M�$�p�E�<��� >{�{��c������9v\�Kv�P���@�;7F�QN�V����t���I�����Ļ���L�ig��]���U~Fi�-
���}��ʘ�?��k�
�����ἃK�o�+ �I�� ��Y�6Pߎ:� �c*@ǒxKb�uZ�J^:T�ҩ[t�����êh*��T.c*�4�?� �z"/޿�5��`�C�����1Z%�w��_ߢA�7���W-�����7�V��:�Y��X�14pAo��2��dg�Q����0�ȟFT��}�#��4҈FgE;�F]5ᙟ�j��'U����#3����{�[4�?yջ7y4��
�s��S���|��>��r/�*�t�\�> ��9o�.����
t�讴���20�Vx���҄"4�+��
�Y(+�j���61�\h��h� �}��}0t@��P�ogoP���S
E;%���D/�6�����1�K�jʩ̖�'�]U�yǨf�a�<�4�#���K������87:<�"K`�u˦b?��ܑ��e
�B��`�_��M�n���׻@�ʣ����GL52�vЄͥ�
C�^�0t��ɮͬ��q��l���jق�]�p�����_������ظc�@��5ЮH@�e7(r�� ���x�ߒ\�{�s�n6�f �t�LC�u+s�����N4O1nP��HC;}5�W�1gE_��!W��u�zt�s;�ҥQFU��J��Ka�A8]y��N�Z�HPA ����3h���>�F ��A8l6��$�v�M�2�-3�+�o�ow�h������z�o,0������Ltn���O�2����F���0�"�E�f�o���p��q����p�V�a7��3�c<����27$3�F=�t�c��a1�XN' ��q���/�c���#_���э[�����u7':0�ی1��&�ӓ�/#Xi�������t�����F梻���O�^f���8�<�2$QdtC�U#�¯V����T�#�	�n���T��%a��@�~ )�i]�'��MX�݌�g� aM���z�A���L����E�=��[6�%�-*]���Nc�Z:a���D�F�����"��ȿN�))�*$��<IV��c>�/��ܕ�����{Xv�`"���}Ÿ��@;��<����d�����4F�ʟ�;��0JEz�KF��z�?��B+���Lu�fl�\/M��m�x����d�w�_����W�+�W�������OYsT87!��և�K��;v���De���8���	sV�9����X�H�$�BX~�[B����Γ�5������@�7�ÝZԅ��uoh���)�o��:�"��x��A�����+�����4�,g,�m���N���醛{8��bFvG>��lCV�&~�E�%��E���Օ��=���<;R��M��1<,��Q�C<��/qL�_C�B��!TJ����׈�vc홺r��7�a ���+� ���>����l��w�gx^��$艍������FUT����F����*�r����� �`8� FU+(�#����1��?d��s��L��j-*�Na��"�=ԗv/�\��3N����hB��*%�Y9m�r��46�S�S5/S3�����e��@n~� Z7dţP7��B�ft�r_�H����;��$D61����PAu���<?�G����a�P�4�,muǀ.b��*��������T�?�֑_W:��طpVUW��hF� ߻��>���i#��lc��:=� ��@r��{���y$�c^cȡ�l?�TՊE/Cs� }��V��hb^p���}�{ʆģ�:�U�C��1��M�����\��u���		�Ȓ�5XR#5�ea;�d\w�I��g@�@�I�M,�s,�U�(�h<
?�7������R��W�W�^ǰ�c�w��C(v���Ea�s�n�e΂�����˜�۽�	"��$
��'2h
@��Ũ�OJ�!:� �p�-�Kj$T���t�ӿ�Fk�TJ}���x��z���_�g�{̰�X?0��X���-=�O(�vJ|�z�1��ޡ�Jhx��>4�u�;'� ͺq��ҳq�g�M�}�g���Yz>���K�D��SO�����Hzox���G�W���ʹ���(�i��똃��vìo�'0�o�Ͻ1ދ�V�w���8�м	�����O�`	�:�-ra�%��K,�SmT��q�������6�"n�[�c"6r��6~6�1� (i0��Q��9�X��dn	��
ZF�nS���0������ 4���A��0�C-i��_s�r�|V�X?���p~|�уv�8��}8~庾�ݳ��P9��lPۃe&$���{8+��qX�[t+�^�����v6�O��W���i��g�3"53�
����f-������o"���·��R�xI>!�=���,pc��X���^��EjA��3�o=J�z<b�ǝ6���H��|�5��=�纔�\��tRUH#��e5�R����g=��A-�Ҥ��PP��C�xNO�����B>N^ZAW�=�q��Q�qX����\Յ�XH0zw���A���O��^8��#��,�bIHL&&z�䡚�:T��j�3ʅ26��`(�r) ��F�J��`ӿX(��ǒ��ZW�ڜ��� �<�₌H�(�f��@��i��D{�y #�;)�$�$5��n� �aS�uP�ƌ����kw3���+<����)��T�1�Z����d2�~6g6���n�=�@�^����	��	qa[�!Ή����#~UPj꽟5\���X��?7����{m|�@�-x�c��Z�t��n{{�B�����d�#�j�zC"��إ���ga�x$Gʞq:�b�T��]C�dUO1�-U�$�1=�1��̃�ҼX��~8��㹶�iG�>�Cݳ #cY;n�r�H�<����z��$C�{co fk9]�n�sh�H'fI��+�Z��#]p]� &�S�rqv�\��d�N����ٓ�	���EM�V��ZG���S+뫚S�I/�~�Y�x�-�Xxzr�X�n~'a�����G�%/r� �a�a�����_&!-@ŝ@�*���1dsoS�,��;�P���#t:��\��~��@s�
��p��/c��7��p%�ʞ�7r�O��U�cuFk�uM+����5S��"J>�����16=E��`�fΜ�9�t4p��	�I�՝"�i�G}`<��8�i�P�+U��2�ZG�ԭqWϵC�5�\�/����߷_A��G�aW��*�8��3�z,�jƸdyi����U<�G"�B��q=|`$���~t9��:�#�E$R��2�^O�mc�U6�����*'=�i�g��)�q��0��'Z�J���;\��#��r:��E�O���RA�{�$5I��V��Us�AN�| 4��׍���m�3�1�S3�H��~~����O��qٜ2��u��.}~{3�̥oS�w�7�qs���~�������c+����ɰTm� ��D�O�n�}5^Z�n��#��#(D	��}�R,*�\Gx �!��[5~��.SX�<r��7���^��^��>���釰��r�w����'�	�m��'
Eca��; �1 �����������R�A@)Y� �x��A��=�@�K����d��ľ
���n�[�Fz��n���ś�J�i�G���=vi����L6x�m*�|8�C#��)�;E���p���h��鬥3ާ�����6����Tp�ԉ�oA�@�:-;,�a`E����1ud��Ng��9�J+׸�ΖzF�;�n�=��ʙZ<8XM�BQ�$H�C��|�uY�B���+K��I}�_����_�J?�6p'��3�xh��Fz$�S��<�+�=��<���D����ٕA7�իyR��O��0�������,$/ָ����|<�u�Z����{�tF��;=L!-�NӅ��4	c��T��ISg���^�4����9iz̓�����Ƀ��E�h��e�����G��c�x�v�����iZ��+;��ܙ�j,��4?���!0���>c�EG� O:���ս�	�7���1�F#��� �x@O�}���-�W���������tŵ;�3'��w���}\V����ʝ��Q��6n��ĔGa��Cb^�Qb�n�ۋ�;�h���:�=i{�����}�I�]����Է�-}&y�]Ē�%_F΄���,�I����m5'��ǋ.�L�'���w�m�0����:S��퐔&,�Q�\D�_�JPӟ��ˍS»���~��������r{������)ki�buo���_�Z�sB�W�����g�	b8���b�K��T{ѐ��fN�γ����VJԷ�������|xqbl��, dS�OBlm(]M*U��-m0���,Q��hM� ���~x"
��]9aH`��5#w�/�Q3��{w\�(�\ ���O�+���cƜ}F��𫿬=�5����@� ��j���X*����.�?^���3��O;!^P��`�(3̥֮���рO�\1qɪIk�ܻ6W����(�f)8WL�]F�{�7Th]��r=q܆Ѓ��hS�w��c���'�DC.��:���a�9$W��;��x���+�׈��y�]FVu��.c����X<�ޖ+�d\��\�6<�*!ڔ�e�yz��G��w}²�����{�?����OE-<�S�.���������X{���]�Cu���'�4��j�nAV��R� ��[��dj���re��x���9�k���6����G]��-;��{$�0�ٱm�djU����j=�m6�T�[{�۪�h��@��d6n#�zo݊�'~�g�⥎��(6e�$m��G`k��]^K��x��r�yu8�[@;��s�i�'MN����&�aՐ�iH���P��a�8g���_L	M�U��[`��,&�3��v:�i�h���	D���C#���C�ž��m�G����� �߽C��m��m��mG�m�ƶ#ж��m�ֶ#ض#Ķ�6[��h=�l������=�������K7���6(���ޠ�qX@�M�����gwH� �tX8�`�Eޟ�*�2,��§\cM}�AN�H�Rk��@SW�w���I����@�.ax��F��\��S]Z�~J�eb���d��1W$��@F�G4�~{�ĔV��C�m��(��e�b��*���z��<�e�o(�ŕP��m(?����2|3�q�L����_�o���h�J�d����4�Mq���K6gL¡""���т`��[C���q(��p0�K��������N�V^d�%x�W +nP1����&_#�"]
*v�Z|�2�tL&��.���Oα�f�#f��Ӱ�qkzZ+�j�^�չ�l�.�G;�d{(���a	a�d���ٻk���5���B�?a|�s����$�'	�`Qi���q�f��V���k@>��.8��Ǎb
p�l����өs������mjN.��2�:���#Q��9t[u_����PN�ޤ�c ��#hS��E�YYQO?ڦ�� �L^�܆�:.LA_�P���(m҄w9ʻ.|!��8���7�RI_�\/E���n����w��c�#N��̢w�O4� ���֘��ڦo]6�s 4�:�/�)j2zכ�M�,|�s?ȅ};���P�����E)���:>S�kZ����*�Z~Vm$�4SMGK�&��{���H����=��]}�ҤI��a _�M�Ԥ�.�=�Q�^���S�����g�!���]��"�����t9tJ�\đ���s��+��mċ�+��$��N�y�z�͑N���!��@���=��oPi��Û��� ���
���빬`^�5QA9��Fy{x{��\8Am ���w����ǟ]XaqA�kTTv}5--�@.�%5/�)+��w���@�>�K�ei孲��2A3E1�����BMkh)QIIq�wΙy�yv{����?��uؙ3gf��33���L�Da����\n$��$�{d�22�nuB>���HѺN�US�ПȖߗ�.L�ǀg/A���$0+�0%�ɶ���V�=t�/gw-��e�>4��'Q]�r��n����N���0��"�!^g�����g+�����Reْ�Y�7�0}>Vi�9~����ԓb��������.ڭ�r�o�[��t�A�[��g��9W������]=gL���@o͙7W��l���B�>n~U0b3|�s�?�{��I|�z�V���69�������:6$��u��;k+�jA�)�ZJ47�9��n�*{>L>@L��F��&�H���s��}��p�_��~h��)/Dk����Uu�&;�y��4�y��7,آm�w:a�2ϛ-N�Ӊ�9��I�T�,�%��!�ŞB.��rrk2��c#�uҔ�V1V���(�A�m��es$���B�m�G��G���v�&\٣1����.�6m�����=�a^1���Go��x�#��Q��[x��-�.�,��a��N�#<�T:��S����^�2#����!hQ5W"yլ�m�ǩ�l[�xm(�M`4�&�˗��:�h{����v�iOoag$F����<%\3��0 j6�yKhv{��A��;CE17�)���/o4��Gxs~�]������}/�N�����W
��r�O�&vh*��!�b�E]��֢bD���&P/��Pޠ�`�:>��5g�^:�������22��㇇���z��7���L�_n�^�J��ޕW��d�ڷ�oT���Z�M���QtvWA���s.���y�^���ޣ+�}E���ݔ'��࡞��ٺ��������fL�I/�֐iă�g�r���.�S����W����e���څ�f�N�o PG��@���J�ډc��]�㍴?ϴ��4U�a� �¹qͣ&/��}_j7.�9Qr�(���ܤ�w⡆(�����Ŏ�=����;�r'K��+���|D�O��w{?�B}X½.��3j�in��b��F�E��,����Kw+�:�SQ�)��V\�(�	��V��,ȩ�6P?d��E��3�7�VԎ��s�����˼9�w�y��ށwUeu�+Hp�	\���j��k�݉v=]���D�;�^>��=��/��y�V��+�x�"�H���%�~V^O֜3n?s�!G��\\��9��G=+��L���{��~�]��^���ǅ�@q�J(A�҂�����8��,�㨻�7�|SF8h�3?���SGh:�M:�9[l�g��T�i��\QϽ[-\7�?F2Jlt��#��kS�̂Ķv��"���!���5h>�N
MgN�(�0�Y�4hZ̺�i��O�`�Z�@��>ikk�A�y��Y�^t�(�w�K��P̿I[����3�b�Hْ�1o�A_��O��O`�N�9z��v$e�J$���D|�0���$���ib떇��]9݆�����@ʖݘD7��I��G�OD`&�)[���NNq+QT���[��k��zp]%�Q��X�U!k{ 8�m~Z/���S~��_R��"��<��}7�ã?Z�P*H�C�D&�R 9���C���tH2S�а�z����7fƀ�m�/����4ɼ.���"p�'p<�%�!�D[�L,�W�a��cC)7��J{�����������=]��4	��������@q�m�
�G��Mp�|p�w�M&a��]��ܸ��l��}��a�лL��4[���u�5���#��cx<��[�T���	&��=n���a/��u:hNgx!u�kG���g�q���v�Om"\5�hǫ$���#��-.��ױS����-$��iet�r��9;c�8嶣1�◂���f
k[��ళ��L��p"fG,9���&�!�B�PF��snR97�4y~}�����������?KɟɟE�TN?�I��u��q�g�wiOQ������,T_���������.#�'"���:%}�[҄ٙ	3lY���=�~[�����:����smz�Ӯ�!%+���}>
�VC�<�<s�}Z�^���1��g��ϱg���f�N�6sN�$��mp�1�>m�@�$G �0��ج�	��}"��=^�"�((K�p���֙�F��3m�H�.]��c5��\(������|�uql�~>�/=m��Ys�~*~�7��z&D��+ek\�ç��G�P	����4���e��4�CL�C򾝧�w:;��M#z�d�U�]gÍ�_�U��ۨX�/B�q=JG�,�_��rY���mk�}-v�1���~��"�/KtV?>扲Qc���S.q����סy�60)��o������E��䝓�\z���Tq�<*";Z�ፑ��%�]ނt���X+����,򄞗�>��y	t�8�lh(�<#6��z�j�l���i9~���C[��q+��d��H�W����r5z�=�'h�<$��0,ƴ�6H���`9Y:����3q*n�����F�#%"w��*�}���P�R�>��Y	���k�VZ�h�VZo���%<�_��$�&{�	�a8NL��!��������v���,rH�THX��y���t�Gc�e�0���$T��<1��9g)n�Ԛ6b{]2��
�{������.7Z������QcP~Zrh��il �.�eG�+كJ���Ph��i)Cʒf��iRO�~�>�a��?�7 �6)^���i)��4eȬ	�Dp%Hs��@G���u������yɝT�(�q �$y�7�����]`��YO�<�+���@�`�P�~<�rC�/�u��%WK�k��=�˝�wA x�^u�Gk�Lx��
�ޑ���u�;ʬ���ۑr;�Z�j�Y�ys�<m���'O����G�������+�04v�]%�,��d�*@����.A���E�_�O;�9�yx�b�����בd�h�F<Fc�@��(��Ţ�QgĊ[H&S�zlA�2-�;�NP%G={�9��?]t4�r�@��]�h�e�����!�@���0����DԳp#�h��k�\�����8��G)y��Df�Z�VΛ������0�hIa��Ɏ@�8���R:rP��L�-r�U��5�N�H���~ߑ����� ��u,o 6DϏ2��!S_�7��_7zVሜ���N�A�\�d~��U�`b��cΦ�Xal��u[�����G�#�i� �/�~c�$Bq�t>�֍l�'EC��e��r��%�=Fz�E�,�v��|gɎ_qQ�q"��t���59���k�q7C��¶��Ǡ-�D�H^0w����x��= ��w����'����&�ި�-(K ��h);��D+��C�������>���sK2)�%���|de��bN�e�m�H�Pd�Lt�߻0\޹��_��Q ���hr(�#��o_p)�lt��B��&��C��: ���>G����Ԍ��I����֕O�d���5�P�;�4�*������:��ҼX�Y~y�I����8V���^�W�ʥ�'1M�B������#Plq���t"�qԥOk�AΠY}!�c'x�ƒ��d�w8A��w�k�$M'x����j�r8>��$Z�B�O�#�E^yZX���	��)�7&����{W+M�4y�����1o��;���_�ӓw�T��_�2{�������E�������.����_V������Ĭ�e��T`�"f���/�����o	]
�F��g��)���v�bհ��U-l7J:J��u��rZ���MW���ή��;�NpnF܁�C"i{ݼyH���!nz�Nr��;�t�7�uRq�F�P�_�ǉ�j>9��@�4%X�p�et?�S�
6�/�bC�Ɍ�0�M8#�4�@�Bso��9�f�(�:A�f:)4�y:��C:P��t����q���
,�*�M�D�{�x-��H:od��I��+�@�����1:��fB
)x?�
�N��Z/��M��_��kNW�!۸j��d�a��r��EW���݅t;���������7��pb���(�̒��r�����
����r0͐@a<#�/7�\n���)����`����a�"��_\v5���]_t5@\K�zL�t7��`,��Y�?��̞��jy��f(�g��򘿨�1�;y���g��j�������t�����)�):�Ԓ�D����
q?�ƪ��t?�Վ��FN�D��{tڷ��ٟ?���(�%�R8޷�Cl�[ �g����r�xH�����d �wC��ǣy�q���1���P*ߋN[WV��^���P��+x����G1L�Įw@}�>��<�6���=1'ix����1�@��[��QMH�����]|J��-POT��+O���ƿ0q��*3f��NV����o�x�udz��b�6�)�\�9�w䟳�6�f�����*�D�qi�Ӵ�2y��Mk�E��.3η=лL��ٛ�wN��TM#ж����j�@_�u�n�

�o�����I��r�]�k�.X��Č	�{Qi$U���F�/,۴���4b��z��F�C%���6��s��Cc+�t��S��)�����W�7yl���[��H��K� K��}�G��w!�fDM����[p�/��H7�@b���I�"F�"Zz{:�Q{���
CQ���L3~i��i�kj����Av����\��)��{�N)������ZG�]����oa���|�����!��6EW'��M{�Ս�TYC���LڵR��^������&6�Wj���kk�ҡ���r/�=y��K-j5��5�q�y^|�M����{^k�CB�|�m'L�d~�]�,��~��5ߧ���_)������ ݽI��;*���H��z����tHj{��Q���ѨK~��Hh�{�/�!�"m;�ն�v�3��5��ԅ��Z�춶8�U�FV�r�Kqsfh'0I#=^�ȯʕA���o�g��N�C~T��J�ң=�;vF�D�������Vq�=@��R��A���1�����8�����ۭ��Xi�N�����m�?N�l�����׳�l��ϟ�E��_���6�T$�q���=�~�^�Ѭ���LA@T��c���9$����#����n	���N��w�[I��gΌc�	5N�]G����'�RX�f�C�\�i���Q��u�
l�1ɼ�� � J��Ͼ�U�e��T9Œ*�@��P�8�!��o�3�i�3�т=DV�r���E<m���"N�')FyW���@�MU�>2�R�����g�xmla�qE�{ٹ�r�v��u8v��l����Q!ޓdq̈́ǩᅆT<$TD<z��K�1�ZP��K��˄�x���7.�+���y�w~��ʥ��'F�%��������]c�*b��?h3�?��x��W���︼WC���qׄ
4� �Rv��U���D��UR�[���ʊ��3:�]1T�w��z��2����R��xa(�?���;�Ƃ����?����K?��2���(�Ȼb�d�����:ǚ7w7o~x�/Fk���'D�o�[�h?�{�m���U�\����6��ԆL�1�>ar�pa��E�A�׳���T�g���^��p%� �R�{����L�K��7н��zpW
�*pg
���> �E�>"���(���]��{����M	nS*w?��
�(p�p��$�;E�c�=V��w����"�n�|$�;w�H_���=½�CD����A�7���(�:pE:x�T�`)� �+����K��J��];�����W�d���p�!�p��6ᶁ{�Hg���4p�|&�w�$�O�т�<���"�(���!h��S�]"臀��p'�{����A�c�=V���;T���{����"}�NT%���;2���a���Q���Hp�����D`��Ƃ��tB�Ao�Ao��"hX�".T�������+ܸ��I�\E1q��!mΟ=����K�	[e�i�<��ΐ��irI$��A�/�BW_�t7�}��t�j7����Vtљ���SBN�D9]dֺ ]h*j��	�!��&Q%|��6��֓@�#���Nd��8"���N��o�?3�y�?����/�q	���mz5�J���gE�O���[����K�Dr�#h���>Ƅ�`0d�p=]+/i���ዔ��	���a\Y�����7��&~g��i�w����[`�.F�v�7'D��w��g�-�i�pz"�&�ۤq�
���]�*�#g��g�%e),L���8-l����9�!Ys��ǳ|\�沚�ϸ�ӡ��GWƼ^����U����W���M��`���-��/���������9�W5�	�l9����K��|�l^v��l����:�Wy���u��r�yR^o&/<ۓ�,O�|��r���i='h�n�g�6GP�ut*V��F͓��Ǧ�0���.�iFmY��p;�E&*5L�j��<4�� @L�
�������y��)˅�j�-�^�O~��k!�.��zb�ƹn<���sL��s\�>5!^9j�h��i^}�5w�Qש4�0s�+�ia%�r�R�z/��ڏ�/�L�W&��'��Xe������g%[x
7�������z�5�۠,Ӹ�8�t�8}�<�J��9��]�������ov���A�"�n l	b��w�nT�)�C�M*vb[�b�D���M�f"�aKU�,��v����X|���{Tl6b l��-@�N� �n�!�C�!��.G�2�V�/�f%����'��%��B�S��@�-ك�4%l6b�ۏ�����e�����������a��#�	�����_[O�hI%�=G��z�4Mʐ&Hv��伎0���f�6D�\�͘LaCg��7v�$�M�?E���i�?��8	����bg��aY<�Q3��7n�,N�+1k��4[��!�����?����`:�z���9s�6��l[�㞕����֏�$�#TTYQ/�9������&de�f̶O�����!<hb֐�ٳ�C}N�J��}´��Y�2 �,�E���K���Q���)K�H���^ Tr����2�|`9�b�����u�7
\��Xicv��fn>=����Z�ţG&K���#� �#uH0
`@�c1���H�\����zX R ��*�$ �5�'����\�k
/�ye(�laL�
��ĭ����x��}�?�o�?�۽~I��v��J��@i��7������~����,ͥ_�TJ�!RD>������϶͜.j�]��ѷ�㚹�3��kCZ�4+匑�R齩�pz)45����ٶ�I�"�;�
��5�����j4p��i����i�|ڤ�u��1�S�Ј����7y'7`�"�^
H�iϚH�����)��� 	�J���4�j
<��C+��i�!sݥ@�TGs�����RU>V��Y��gE�5n8cҔ���dye$5gc�)3&d=;l�_�;$ê��:er&&��';lVF���,L6�zH`�6Ֆ��+�w:������Ӕ�6�W�FS��P����NÒ)5��9e?�cR`3�Ǯ�b�&����|<��W��M�_6��(ڞ\ZsG��zX�M����X�����c��7��v��a}t��Æ�c��@��]�`�c���	a>�-"OI_�������ϴ��_�_����p��#��	l>����R�J|�+��xU=	^K�x�
D���5����I>�������>�:6k21����L5˭\Z�ß���o�_���"��%�'������]���n�z���- K0<g�m�	l>Yj��!��y����/��x�Pء�r4�1�8���y�H��5�r�${����o���<sMG��
l� 9k��M><V�����<[�`2p��i
��O`���Z���%޼��3����w��6̚�1}fֳ
��W`��Y�<[
�y����\�?#�gd̝��h��O`K��Tc�n�������3�O�=k�mb�#0���w����y[���"���&�	�}D�P��i��yހ yEzBS��֟pͩ�?5&\W�[���v�f/��v�{�k֯o�'_e�8��L=*]�tZ7<ˍZ�:��#��r8�sM.x��>�?v$���t&��	�c^7�
�Ϯ>�F�L��Y��������Og��������1'?��)oP������6����Wb�߁��j�+����8&�O-/O�	�4�`�c=iF�W`ɘ&ڢ�!�̥4����J�w��6��.��� y���a_P�뀧�Z�\E�:�x�M3u8�%myqk�MVʻd�i7|�I;�%^�W(��{��z���E}����~A�>{�C�7���?z��Fދ��<��{�k>*6T����Ͻ0�˶=�d{��i��ל���ezs��&K���󮃣��Mx����C�P�4��r�R��ְܵP��P��'���'���QXO}�R�iH�;��>��_�[Ԭ/Q�U��^�ڃTF��[=
�n���G�@�Z�Tg$��]=
Ӫk�T�@5�;���!�6�b�Ѥ���P��]z��T���ո]�ֵR�C�!Uw�X��Bg$��R,tnÄ��$IRVG�=ɑ��<�2�1�@y�Hz7��ZN��	U�	'�� ��,]}S��X
)���b�_��4�u���dU��*��%��k�lH6��+ ��7X�T)[{����=rU��-0��oq��w�Y�5��J��;����2q^������3�G��{;a���l��7^(cD4i���!.�x��f��~V��T��qZd�ִ��Y��w��
����k[�j�]`�Qi��@,�����Th�k�R����+�r�׸M�w����N�9Ӓl��)�)��;~���8c��\�m~{WR�!�!�t�O�u���� �;/I�>Β��}T��V�SJvc��0|�-�x�鐳#>��nt,�EK7�&��q����H;g7v@4��߀g����]�=�d���"]
�\,q%fk�U�9�<췌�w���r"9��1���ك���B2��Z������t\Ow�T�rG�Y"ſ������1�m��^���:Dh�Va���JTyRܝb������������\;���&*Տ���ː[
D��|�!�p-��|Fy�#�'��m#q��l��� �X�f���A
+:���}'n��1���Ӛ��Ic�0�s�6�5�%��fh30N��(� �^gS�=��G �x��$���-��K��WʥH��댷�n�����)IP
�|/~ݏE9Mi��)���S�P����v��P�26��0(�{T�����	�n�i���r��r�װ��y�Y<���5D��v����
<��?�_��Dz«�R�`m�P�oW}Z(s�a�*Q�-􄶅B#;��B�T��'~U���~���F6��1�{�"��1��m්>��:���9�)�u'*�)M���W=�L�e�=�\�λ�+�6iJ/x�G���OO/�9�y��\�=W��+~l?SK�"���`�6"����/AܚM���HG�:�]i�.!�0�q(`�R8�����
_v��s�#��>ֆoK��`�#ZN4�s`�?��`�cuƎk�R+t{=V���6�R|��
V3��W�T	%mE�Ӻ9M���h ��:�8k˟C��d{�Jk��z%�
]��]#s^r���h���hDSʉ&h��� �<��"�\?�F͓E��P��hsߣ��%t����	>��^�+c/�5W^rWp��^ó���pyLz�rM�O�(��E��9T���\^�Dy�C���=i�[�VO%��ɚ����i���z�����J�u��V�6�)"���aZ5�[H�c�)iUj��B�Uv�z����z�u9IIk�6-ݛ<�9��cڴ�͍cr��PfɺZCi��k�3�F4H�ȑ�O�Ud�}�\�V��M�m����'���4_����gk/PU���m͹�bV �\l�q���f5�������?(Ϳ��v>�<�5�����g�H�*w�_@A���������H����vB�0Д�C����?�{5ܼ�{��Q�z+Vz	`��� Lo�J�� ��`\+e����a>�_x`�� � ���:{��~ơh�,��!k�Nb��#KQ*g_A�)�nTe�<��/R#�s¬g2G6��5h5�}��n<�9j�,C�><$��4��!ocHWb��B��Rȧb�!ޢ�S�!�Jh����Dt��V*���#M�����#?T�zD�ɑ�(�AdG�	d �� &.D�RS �2b&fg��X�J|�Q  �ft������J6� [�A0�������M伌N�u�Nǜ��8G,��(�I~)@�G�*��x�ܶ�l��	|�ku|*��_i���5�������Vo��X�0	e�Rɦ@'��b�?�-���KY��I�yQc��*����������A�ɭ.|NA�Y#�\5�����������m��䗠���(c���1��(jA��K�%����e��I���D@�
#S���WVsc55�<ر��5%4
{5#FB����Ьv^n�;n��^De+�G��o��V��GtFk׎@|]�2^{ϼJϜ�.rx�$�-P���@=����kb��� � �|p����X�/@��.V�'5~�1��
�,@�� ��s�Ы��b��'Q�~���7@�.�����x?�^���ᾣ1F�s�˝����]�`V��L$��'������`"'��4V=��9�h�d}�t��"��83�;c5��lӰ������n�����{��+e�/}֟}��gQ"�)&Q9xU��|���'Q� x����y��ۆq}�f����݁��
�[#����!�7	��y:���jt�6�����{��=Զ�gB���.�
pW0��wb�� F<��J�ܑ�~��� ��� g��Ɗ��w�S5uJ��i����Q�][���?�5�CrRbU^$��;=$��D��ċ���PҦ�ċ� 9)�,��kp�$ya���N�U�fB��"�	��RS;��3s�����ae�Mo6���-���߁\��\;;�M�6�����^�Ô�ٵ����-p�����M�tf�Lc��bjL�D�F.]H�X�L�jk�A��᯿�Ng��ǝ5�H(FR��sf�㠯�1:�*:a��z�����9UUNY6d�sU<��}�;�,��~��9���J���l�x�IX��7x<?��9����/ĳʪ��<����>γ­�^]V+7���I,���Z�jQS^s�̋r$����a},�Ի�G��S�z���� 
�	�w�� rz�٠�tz^�ҟ�t�a���PW�����Jy�����>�'�Fx�J�R/{��F�[[���e�K,�Ieo����fN�;�}*w��Xn�� ���}b FL��>ګ��%������ڠ����}mA�ć�E��]�{�c�pm$��W*��߰�6�5/���x��?h�|���@�� ��}@_6��˶����,�s
�j��I��#�r���Xޢ��}��?͞w\����������XR�u�g�����@�m,�-�E��[~��5>���&�S�[�ls(��7`�ԽiS��v0Z����։�B��l�^)����g�$n�hrwG(�'��	2�A�L����A��*�v����:�0�l��Q"~���������	u��z��થ�0�d�)v�u׉�^<4AUlT�ǃ:*�{Ʀ��:*]B=���^Ps=�V��*��m���1W����zeo���,�������^�X��'3EOfl>��Pc��S��m�U�sU�*M��՗��
}�ח�}節��e����ڬ���yƧ���?q�y�G��Z�� � �J�x
��I�t��.�� �+ >(��W �P�m�q�i�/U�����}�dy�i�Q�~Mi5�T�w���ѝ�}�����x]�ꅖ|�4EB��7�ꄪ,+���¬�ʚ/T�ك[��r=����H��q�5���
���a/E�˯yP��Q���?�·���Z�6"v��rsm�]RQ�:U_.kF_~���oC���)�+�6m}�@
��6�4��;�SՏ�1�� ��� �>���J�����
.^�7�-�|�{�
�*��!S)TC/K�Xv��Ѕ]�T�>�:�p�Y�+��Z���d�n���*��`�J������Jj<M�y/2l����K��z�k­�=��nw����*�`|�zƷײ�"���b���u����	.�~J���O���R�۟�J� � F LX ��gMƘ��J��M����Wo^/5�K��]7[���Y>}�9���i5���Lr��F��/���R����]��Z���5���}*����Ͻ�tCT�5���|ְ�������x�� ��!����V��u�͉��r��`�o��~��KZ��8�Y���s��uw	���_��-|�ys�5�5��� �o���T�{)Qt��<v�P^�Oa���z�&mM�gk~Fy}^���j� A���M���	��/Fs�bO�[N[9};�ӻːw9����>��-����마�׸8>���E�0 � �(�0f3t���Y�#��O� p[ nx������B8�w��G�n
�ǳ��%�2CT����x���h���˨�է�"l`O6�~��}��5KK�o�X��nwx�Tc�
��
�ZO��ky��<&�n�RL)�9��g�7���/��ܜE�V~ކ�`-�3*HSʣ��O�w�Ha�Q6��^�2�K���i�.�p[q�� @<�X ��u�*����Z����A�� �\*A��Fkn^'tTR�ĽG%��qQ"�I_�1�����|��5^+8p�|X�ds~��5�k�vNR�v�B�\�#h������'}��hC���l/_�F�`�l�=F1�K6/Wu(�RU��<������$a�����&Ag1g���Ky0�4na���S'�խp���_��<ë�Ķ��Q[�t��3>���������z2����;#���4�T2u��B�]��(Z�>i���=�C��8�������>�"gO�kX����>+Z��q�=)v8|��	��۱��|(SҎ�_�6~k����o��p��e����� W� �������]�Ͼ��nc5���[>�N:BK���A����9jE�!x\���рK�6~�Y��ę(*I8�>`��i~��Ҝ�C�C0E%��;�Z�q B#r�r"7� Y샜+r��G��Q��ӢL��N�Tr2f��m�l�pN|�?T)��b4�w�%�VJ���=��e,�Q��#p��/�W�Z����/�!��m0��C	��� ����_�4��� ��X�
�ïhH��}���ǹ��2���m����p���u��~�RS����wM�{N����C��{���fo�K]셦Q[��~|�����q��U�}zgO����'s�HpFР���X_��!4(Y`؆y�Oť�c'x���:�7j��{�Ȥ�}�&s����� V>(���2��̓�\G�� � cf,ܡl!ޫ�|4q@�B���j����_Q�����{�3�@������FL@�����:��`�V�6�C�C�j��3qf�%r[=x@%�i:R���MZߡ�̈́��ivY,W�;��QvY�0;:��B�W�I����#��G$)�Ɇ��"�ɔD�H\�<�"��M8�˘����&�}r�0��{���nM������؁Bb��H�@��H����?;��C.�/��b{� RĶ����Q��o^Q�&�wj�(!� xKs�|�!<�]Gm�ޑ�(��.������'���H)�п�l����s;���[���^P���E�B������������X��P/������b�M � ~���@�X)��z7�v��M�GH �h�� y o��i��To� ��C*�z�}���^�Ώ��G�D7��R�" �6'��kN�omN�Ӝ�/jQ�?��r���=�ޱ7�:��Jj$I�t��	+�m�K��Bp��[E��:�v����Dv*:�*_��\:�ໞ��C%��04 ��Vi:���z� 0`)�G_ku���t�{8���w�܌V`�4�
�������7�K�ϛ��5+��ь��b(��O�O��o�x�VJ�Fj������yU��he�x��#(�{��aME��x�W�jQl��Z�5+bB X�{@���k����T�w����j��_�S���͎�S?mv�����m�k����͍�&HݓVsc?�_�d쯾�ٱ�F>�����o?���_=_3��
>�/�������/8n2�/��=�'m�2��c�%>���+m�p� `/�v � � ��&V�H��ߨ~���[ �:�&�# ��Վ���c �Sʵc�>�W�,���D_o��`p9��E��h"�r�0�b��k~<,����o��� �7Z�	r�H
MЁ��&|��Ը�p���FQ�v�(W"MR�S�.5������k����I�s�II�"5��J�m\j| -b|%�>hE w	x`(��T��~�R�#Ȁ[�5� �T
��������F�3�J�jF�<�i�J!o��W����W�h2���\��h"]4�;��M���%���y�Wp|cy��`�)qH��$���1%�˛�UyS*Bh ���=(�޴��V�
�P����X�%���|���'�/+�ċ|L�b�x�}(~8����e]�\�܈��R
���r|w����=��a� �ۭ�@� ���dF���ޞ[8,c? �y;��ۖA]az=�؎ ��H��:�҈���t}�?[{�[(��B�"��.<ݳVnX?��z9�.�M��K�q4�'R����c����A��M~�6=�KT���i�hN��_p�؋���%({<�9�r�=�M�� >���u��*1��}���j�_��Rs��]���s������WM�8��Ho�Wo���0�bw�º�=��d{�Ѱ���	�),d���}��p��^�	ƒ�j� �;�Ȱ�X�U�_W4�h>�.�k�\�4R�==IՏ!Հ�R�G�, X�@-@�0�:�!@p�tH�#��\�� % ��@%�5�f���L�t$S��}<9��-��>`���t�%�{o��<|����A�ܠ���{�i]6ww=./���h���|�
��.U{�����Hu
;�l�{��W)��S�P�/��
ƾ'
�P�D��� �M~5���4���
e+��B��S(�I���Dx���T
?�r�m����O(���hVs?�W��gE^��;0����gQ�%|
�_�J�C���`�G"��$I��S�[�zE�B�i(��;)�=
�)d�]/�� ��+�t��U*�n��0�\K�jw�=���tҌ��Ҡ��[��(�R|��R-��\E�G�I+��^��&����{nC�y�[�9��A�~�_������G ��X��#*M_p�6X�i��\�,Ԝ7I漩�'���<��!̍������f.��T^j��۸|g_vƂlS�g�!:ET�^BҘ�A%
�+H�Y/V�=m}{��mR�F�z��)��mdV�ۨ��!]%�s�2����x�4}�B���@�ދf=�N4��NH���Lnñ_���A��q�C�[���	)��*�հ��n<���ׁ�.�X�U�Q�T(��1�\�2�(�+��gE��a)�/#�/U�� �NI[�"v�)4�yӋf	kO�-Qh��(>ϫ��F��zQ#�Nc�ƙT�^ m{�P����ܽ@SZH����?I/�P���k=D���g-׈���Q��q;Q���w7m�
z6r� �BJ����{+�xg,�6&��������e(���_k��;{l�(����ԉ�5\Ln���Q'����nE�T5���P�`�Aw�J�٧�i
^�=��JQ����[��@Ɨ�[Saf�y�x��/Ư�\?�~QQ�D�@��ڿ��3ћ����/�Ұ�N8��|�̭}�j�����n��1����U��?~P��K�(L8UW�jǱeXuU����E�ϧ������N�����Uw]�0���ݡW��z!�ӣ���,�����fT�A\e� �n��7 ��X��8�I 9 o��@���玩~�����- 1 ㎑�b@)q�ॲ�2��ͪ�¦���dP��NB/g�a�����k/�C|u�������!�_����B=a�.��K3����LX�?!0�K)��$�6�p�ᭌ,�q�I��,i������	*��	ńMG>���:	���	���b�~\�u�:�zc�B��q��o/��C'hT��P{���FT%�4���Ba�x�F�X��E;�a�|��	M�Mx(���/��C��V���G�����7zEM	lj
Ǵ>��"��B1PQ(�r����Xi�I+���_  �N�J<~B��z£P��(wp��I�?SP]��	��U��PQ(6"E��kE\��jQ4�U(��N�6@�j��{Y�5���.�6I�o�AlbQ݅��A����lz�P0�>�Q�����:�[������OMobx���EuB�`����J�����P%�����:�Sm���c�)ɣ@@�	m�����2o�`9�.�6��z	���M�PX_����
��u�`g�R��q�9Z��}C��]�
�#��E��O�>�8!�w�e!�˸�pU!_Q�xY3�w��>H�,��.����ѳ�� �������8�-FO%�SKZ�0�vx�F8TH��|`���y�\D=���씷5���ڹyΏ\v^+A!tp���<!dg3�3��GpVG��s	���9W�V� 8�K<2����Șflu���뻪��L%F�����Q��K����yM�[��:׌�|��Ő��:��S�RO�d� �� ���t�t�wpvZ�#��x`4�\�e�QP�<�����4+*�~��'eT�5��ά��]��**�7+�r=�,i"*ޭ��EH�tQ��nETZ�`�����TD��8���%*��*�r�6;u|��������g�k�ط�#7����Z�{�&���m��͋=r�O���V$�žr� +UD���>r������'���=�֊4�[�#7_V�&ʺa�������柲����ᑛ8nT��~��Qn?+�8���/ ��+uH�x�'�f�O�_�Me"~�"��s�v!�Pd���M�|�"�.hVnnd�����������Q#��>rs=Z�H�M�}��ᑛ�,{T�"_X쑛�{�I�
<rS�[�eRDc�"��T��!&E.V/j*7��?C��cQ�YĎ�(�qբ&rs	�.X�{9��r�|�Vn�9�r�X�M��s.(��%����	�Yᑛ8gN� ��l�C3�?v�O�I�䢤[�e {A3w�.�ϝ�yL�-��fk���oyA3w^���o���@�𷬥���/s��#�Ѩ�_hd�5w~]��!86��?އ"��$�ħ�"�=���矢xr�5r��q�>�!Cm��&zW�m��h{��Խ:h4��{���Ot.3�t&C�e@�ι��(g��8+Rѝ�|�x�=J�`Z���^����b;�)�����{�.�9oƲ��R��T�{{=��'��J�O�Zq������z�|���?��O���J����/b�P�����}�٥f�m$f���_�l+�]|�ìA���H�(|��@�1V�r@�f��v�����ņ���:��֊@?�1#-�D�Ȗ�	�R����F�^�j����IO(�^�<~ȉ�G3�VI��{xx8��.�`rę�7S}xYI��-�2���Wx��k,�4��/m����A�4�g��1yhxR@�/��ީ����D��)m��B�|Du,e_�W⬎D#������(k��/�e\�{A)���8.P�;&pR�\��ר��U��C�{߳=ϒ��&ߠa�JkD��)����ȡhT�x��xz�Ƕ���X���8m������ж��-���&Ԯ�?���s��@�����/��ӟ�zE�n=��@7�

�0�Щfϳ:�9��t�V��k֜h��,L�Na)"^�S;��f%���\�Li�!�����}�m��jv��f���Üv��N~5��H[9S�7޳��Wg7e_��uN|x\��X�%�s�|0��ֶ6�lc��j0�ϓ�)1��p	Ɩ�_uY����ol��2�����K�q�z{@v�(=L�J�����S͛�Sp�wZF[��sLc����=RAα�D&a�J��b ��+~[�=�=��ys��{��$К'������z����ŏ;�ΙGX��G�oب�L��D9!TN�D����	��F�~>2�����x���*���x�q�4�s2!��8#��"�6������Z=���Q
�-fvz~3�Z#���c�� }{U�����|V�w���p�mF��A��#�\�y>*.I�q���T��"�k����J�AK��FE���l���&�����
MM���o	˽��Xf�_X�����Xi� @�c���.��m����7CF�ѣ�v������F��9�Q-ga�;�U���zow�SS��>r����}�K��!�ư�<̼_�g[*�N��ߐ��JwXKu�Ju	6��cU�$���R����du� ������_��X�۸s4��rZ�N�ς�_ 3����ک8�6\O�&�	�t��r��6D��u���ڬ���a=mԱ��^¥��~x�ӥ�[��zѳ�EH_`�	�3*G� ���P����)O��`����x@АW
�/9@O�N���+L8�s>�V֩+�4.as?�6�p���(�,�-��)rrL�1�wZ/|t5��В�Dm+^x���c��5aￋ��©�(�:鍒�[]�f�`s���`�C���Z6���o�@ �ʠ�ءF��&�t$v�%x+#�����g)�z�W�XnV����gz���\8����o�C��~O���0� F� �H�"���m.n��pC.j���t�>�CzV�����#Xy��P�w��vg������wd;����Xg[��|��yӐ���o:�>t�=�<|WҘa�M���7ya�8�X��זL�v7A5{�[�����k��`��KM[�x*[���y��n-�����e��yGK��U�#�����[s\P�fk�~����?QXS�=-\��N�T#ۅ�(k���y(r[k�/n�B ;�'=/0�%Td��c���er����p�8�f��_(ʖ�0o�D�8�N��K�$���*x�O�잷W<nv��
�"̀x�p��H�i2@�&,��b���ʫ�/̈́�j�y�AH���'�޼�G�f�F��AXV�4し�Pr�9Q��
���9��*��?��wjg��� \�;AԌ6,pO̔�4��M�x�f�0\���K�M�A&qf��[���|��#)֤&u1��]���|��^>���")��T2䬜S��>��v����N.7� [����Z��M�2i�ao-�om�h��{��"-�܁�ɀ�qd_D~���B:�9�H+	��($L���8���.ҹ^}�o)L�7W��ҫ.|3E�gF��� 3�����2f���\�������Ss5kBg��}q��F�&�^�����6j/X��:�e
����=2|(��#p���Kmw�#��	l���U�9�`б��1��.k�w����hI��p^���g.e�j�A��1H����x��6�����{ ��hFs3̛��ac\����ã�A���~�y
[�?��P�}��(�B(s�!
ey0�*���:�!�:DtB�B��LO� �
߳
�m��;r�:'��7o�H�X����f?қi��(5�xC���uR��fut��_i^V�w���1�V�֩��WIuN�֡�9�g:\���@��;1*�[��<�.Cz�i�'Ek��K-Wc�0����o�[����S�S[6z��ޝ����n����'陯_��LX0.�Vν&͋�d��h����@"��t��3O^1yZ�7b���Ih���C����z�_p�&U��J�����\gH���Eǥ�� x��d��^�o�F?o��T�^���tBGB�w��4����;_ob�~�|+S��k0A%b��ټ�n,�������h�#il�c!*���;������KQ��o���v��ј���};*��GC�B&=Ak�?�?z�rhf��rO�'�R�n�\�����6��qǸRǸm�q'�N9ƝU�΂���䆂�kd�:=3ޥ���L.#�]n���������p��1�q��x\C�OM��|~t��#J�<�6����ݺ�y��G���sz��M��!���0��^�����Ah]���s�2�h}�ʟ1r��_w7�H[p3��4
����:�$��$I�,�����Wx(��}�.�P���<�� ���w�#� ��eG���'�/P84�|P
߅x������X-�V���
OI��{O@S�Iawy��Bey�I�R��9�q*J�RG򄪰���Զ�,�Woa�۔���|BT����,��g.�y�#���{�]J������a��v�l��e�g�q���5yg:�"���p��k�:y�W�Kh�}?��m
޸x�=>���a�jf،1�Xkkg..�%���'k5�"�y�b�3w,roޜ~-�L#6�W�ʐ�F��������,��3tU��A�-��Z�3Jue��[[�"���2�m.�����#�ĕa,�7�>�q���rr��U���Y(+�K�1R��q�L��1������K�֤�dከ;���V� �sK��νI<\�ey����I�5�n�?z��m�v�<�J�Z��H� 9@�l5�=@�<��>��?�W8-b>�~g�W�':�`��HG��Ty��H/��u��d��A�y�&�-�sI�q�=�]H�D�?��0aȭ����DKԎ� $အ���:��^����^��f�3�S�������|�+��7�������:QVz�S4�$�aOb�7��(���.����U���[<	ٔ�����@��H*+�V�h��,�j��N�lWV
>�V��y��SfL��L
��V���g<=c��8Ö19#+��t\愬��	3����)3gڞN�6s��h{:͖5e�dpd� 7m��ـNΰeΜ����	�5���P���-5c�̬I�<�,넉��~�W����gg����fX�2s
Ƃ�)Y3'fL�geB9ΰ��K%���%(%��J�����ʃ>Kh|S�y=!^���^��X�zieX���7�0=����͏�N���~"�?JW�wT��y�&�H׈���^:��o��2lX.�2*M�2!*(�63+c��������9�B1�3���lz)P�j��+tP��^*�ίi�7�fl���p���>�8,�}�\X�����pTG>*����_��i�����)��w�w�a��qhq��0>T����gq*'�&�++��x�v�F9a�F����m�Ǵ���g��~@�z����I�c����e�r�,��p|e��!�ڭِ2���Gp�ȮT�h����y���r�͛C���?n�C���|�U���b�g��i���{���K�����Q�)�Ks���F������Ll�8aI�<Sc��!��`k�R6͋2�GJ�����ah�%o��@�Xݙ�J���kA�iЃ��@��s��S�
�����I:9�,K�(���<c`�R���у�������oY<6�}�,�����=�7�rY���@����*8MJ����͍�2F���!��B[�C>�7~��>��k
�|�h�G����Eu>�{���n�����I�e]Nqy��[őF�����v���<�v�tv�]�ڥ���6��ɇ��wzt8���Q���Ҡ~@�[slu��xP��z_<
j)B��� s���n[����!J==a�Gu�\�mO��u�}`�iw�$e�R��>[�biXa|D'�a9� �M�,9?Y|W���ţ::�K���uc���O�舎��_W�O����,�j�0�#�u38�+e�FU��!��pcϱI�����T�M����+�����4���^G94��(�������P����Bķ��t*��:�\<>b񰎹}ߐ�~��o�3wJ����z�Ϳl3�:�&N����^`�)�9�KN�
�lޱ���+s,��% i�IW���=#��G?7d?hk�u�n�X�^d�~.�b�	��]��x|��ź�k�� ���,=�̾	p�C��I��0��S?�̼�mh���6��A�-?�>��_�d�U/���ͧl���<ǘ�0�5ǜ�ʼ�_ww;`�{`�gb����p��Q�ĳr���kOU��ef`P43j٢����"�B�A�/�+5Y>C �1J4
)�'��m_�ۖ��fmk�[�G�fZJi�m���$�D���s�{�ޛ�����=�{��{��{��o:"աrm��n�F�7��i������G�ig���i�k�(�`�QREK�ѯ����4>ɇ��|���ߛ�e�!O���:�� �l���4�_���ٮ(?hd<�EEX �x�4�}&V8SƩ7������滴�����o4���6�][A��׵ۤ��Ҏ�$2B�B
���}% 99϶3��Q:I{�pY6_ʜ��eB�h�#f���n��0bqbĶ���7�ȓ7�#� 쓦�,w�.�!���r��XS�3n�ע�w|E �J���"��r���lʶJKög6!P�-�8?Z�̇ay�B��>�G��A�Ebi���UE-ǣr.��Un�����9�|�E���A�?��?D)>¿M~N�0��|�����+�������y�SS����� ���{g�4�6'gj	핓L��?��1l`��r�\>w��ƒ�w1�s$�u`C��1�'Yu8�{���t�7��8�4�|�� ���p�+�$��O2��#}$EI�����m��X�߻�{fm��{v{��C^B?7m�4�o��i���冖i�t�k�Y��	�����X�n���>D�G��/xRM0��	����s;�s{�g�g���\�P�J̵�����r-��߷��E�E��6� d�xB��u�wO����x�^)�m��;>ǈq��$����un7@ +�H�����8������,~Og��>�k�Kc�գ` <]J^g{��Kʉ��ZϠ7���;����A���	�e"��P��u��v���ؾir5�����oO0Ʋy|� �_���߆_��/Q~'��L���[k �@�����/?�-��O���I����H��k!���V�ۣ@����Z�ǒ��rͦ/��-E������j�������т�g@�!���`V�5��G��z�`&���'�������?t!� 0����J^W� ��IG.V��qD]爩3h۰�}*R����͓�0�~��x����\��Qt�܌�K�Z\��\+���3�ʵ�I'u��^��M��/�-b3H�Φ���^�f˯�_����H+G�.��ӂ�J�~�1l�l�>P�lh����d�n�T�ø��l�U0����u]sLg�|ԟS�.���K��<s�B�ޚT=�;6w��oXY���T;2 4�%�]�6�~u���k	��	h56Rή�~R��&��{�|��]t����~��Ѝ]j��9��8��k:�����{r�@3��o1ٜ�����c�޽㿄~�Hqկ�~��� k'�H�҉[X]��|%�>#>�̈́� �2��j��<!A;?�8q���V�?�U,e:��Emw���.�B��?������=Uh_���	�^�Kr���c}W���&9���K�Q�X� ��O
��~@�3u��;E�M��b�H
�H�����ߢ�}��<M�)�Q�����[��D��u�n����tU���p���p���-v|4��:(���m5}�����t��'�؟�h�ϋ|6��<~�{F:����E�p������ߟ�,�cY�f���d�#O�[�-lP:�Ep]W\�n���+��R&���3�1����W�/jEi��|���6��SC�� �5��z�^�k'\���}��'��iOB�}���A��ౙ��4��Y~�N�{�O�fn$����f3Wj6s�ts�y���j��������q)�*�J3m�8�,��f;jo��� gY�٦\����j�Zq�,�?�?�F����۠�-1�� �<l} ��/]�e0�@��Mp��p�hU��$'��e�e�&�?]~gR:�c![q��w9��P��F� e�C�����(#��
�����}�c�f���
� F���;��Ə	����8r�l�z��m0��#)P���$A%�Mٔ�$��w�Y��ݠ[3x����A����r�J�0_8
��+s0r9r�΢x�L\
h˗�v£5:7���)�%J����6x]U�^�e��*w�*+�ʼ�U垲B;�݋�,,vH:s8s'�{K�o�,�,��STVXTiϝ�EE^���4v� �a��,l��t���lz� �	��|!�eMKc�pu��e#s��\�f�5���i,���c�#Pf\NO���(��������L�`��4hC���Ԝq��7��D��<��~n@V02X���,)-ҡ5�V�Y�2�E������x�ڶ����M</0uN+��"ӊ
,̂l�`���w{P#��f����i	ƾ�1=g%�w�ʾ�x2y���ۍ������&\�Lχ#nў�)Ee�¶�3����l#�L�5g�6~���$4�]����J��y��$�s�9���^Q�iE���E¶�2�톳��Zg�����߈S�gFe�`$�m�g��)�U��x䚞�~�����Aff���
��ݔ�8�B�.��烿����%��%���/(���ݘ�A�5U$�x��\��[�89�@0N�n�DB�q��M�oz���o�-�3���+�����Z�
�u&�M��#N��4D�f؆=�ź>0�w�������6]w���20�o7g"�Ѓ�4�K6L����� �F�fì�7�������+��nlAAQ��w5`� �V(��{�0��}'��q�����u0;���ix>ܢ�\,���ϯ,J���;_��-Z|�i�S��P�o���++�S)���T��.	C��P�C��VU�,(�RA��z�xQ��.��5�4lY��4J%��,��.�ϩ,�++��W�,��(��� u����c>�|�-�W%���[�� ��x��j��}�p����L����N{�3�GHB+{<��I@�i�H]�ku{Jy�l�K�F���,�a��&6`a�c9x���JQ㊼�е�}aƊ6��P�1�|I��j(�B����Nv3vH8�~���,s�G|8� &�'����'��W@Y+�Kr3J*��.)��;����1���5�ݎO��)��Nz���R�?lh:m9�1e��:/������
�����D� &�M?���m,�n�j�b��t�W��xoŁ?�]�LF���.H�Z�]<�t��8,���y�0��^��Dj���SD��"�'�s/�i�H�"}_���y�-R�H�&��ENC4��bǙUY~�ʏaā:v��%B1���B� ��X�q�cC���'��K��+��z��BE�E��`�V7	Y@��ȅ��T�X�H��ѿc�IU,�x�e�{�y���'�O^K_��X�wx��-�ж�D;�оL�/G8�f�ᩮ�/�r��D����V�h��$ğ�P)ZT�\��KCE���MZ>��H�̒�*��1ay1��̊�%V�"'d�����(1���i"+�JѢ��#��Kn�`�PTUzO<~*�TK �$�
H���' J�eP���N��&��E�h?�� 'bZ�b�tJ��:�N��ۨ]}���_p�	&��7��}M�xP�a�U�逕�f���+�$�bTnP�l�w�$����X��`���p+z6�d�NQ��K�[��GȲs��*Ȭ	���%�ly�'/�D�ʊW�Mzѡ*�P��"�a�R�U�ё�G^lԉc.Mg�w�����NS'�4�t �à_z:M5s�n�p�52�3��m������b��]�u"-�*�6�4�R���.��[��k���)�Xn(!��L�.c�ͪ�R��P$Xq�n
V\&���6(�@�p�U����(vp�n���M���
��9u/b)o���R�>:���c�q@�
a.���`/#�F��*_j�����]��������mt+��|�*�N'��h$g��#��u7��X��;�z��Pr"\ѹ�E�U�;�U��`ji�͕ԄA�� J����r_eA�ÉJ�gv�w��񰧩j7V���8 }�z4���q~]'��+K��Ϳ�H����Z��\���z���.M?e�{�H�5�<sK:k�����j������<���T�JͲ�f��ஓ�Ldvv��|�_��\���q�� Ϗ�ւ����Â8��#���<8��l�45�`��nF��z`m̲�r�K��$:���<Q�� ��&X ��V𭱐e|��y�\%n� ޠ�z���(��(Ϳ{��?�4 ��'�H-��3�+�Ny�E�����}p��#����.�uѢQ\���@�35���%�1*������"ֳ��#9���Q_8����M�n��x"9CH㣣8�`ÈM0��y��1Z�N��3��2��׺+y��t�A�ր<8��;!��\k�Z׊m���t�O��.^�%���d.)�25��EY"(�J�;3�*
a���9��=�KbEm#2O��E&�bسWr���J.k�Wq�L��Wq�R����X��̏d))��L��p���x���J�r���{\�zr;j���^͒��`>d����%y�#�0$}�3�Dcf'�@��[ʊ��i���y썭����ȕ4�A*�P*X����@� �v[��e*t{dg�p��Z�p���|����p%sB��̒�B$����[� ��盽=���i�	b���PԠQ�`��й�'B*�m��]�l( �:<�L�m����x4��;O��4l%r�G#fu��e�-/A�.�x�[�_�-�İrبK�꘶;X�����q @�a��g��NN&��ى�q_@!�G��<kWU8�Wbba~e|U!�|z~��(�<I((0���(��MqU��B�W���G���8fC��0�h�m�I���S�Q��?��]��z�dtd
���;?�˶��\�i� ��0�Bi�T���f �5B����T��������'��K5L�ig�.�3��;�ʙC��V~�gct�tp6�n��]��w\˝���5�����{��]��=i�zO�~�0\� �׶O�Y���,���_@>�ݍH�zx�z?�=u���֚��V�.�#���ZW\��!��� ��� v,\�>U�,r�6 �ֺ9����ud
VƐ'�	~�$*S� � ��Lm���N������d�4B�+��L�<,N�|�bW1wd
��p�f\˕��kQ�c^����]��qz�e_Ǖyl�O��]��Sڟ�/���iX~ �f,^4��ٽ�d-�b=���F�#���t|>��O��rcz����(�g�o(=�]�����͔&��(�=;F�l���C�	C��Bx,������7�2K{��"�4��U�6FY�},���+](H�VT��B,}��J����Q��]'|��9d����B���e���w>kl��
]�֎a�J��B��m���_Ųw��;��*UR��4Y$:B,J�B����C�3��pJ�
�~�X�����$΂��}���$��`?J����_K3FT4������a^Nc�ƅX8��"����N^_m�0:}�P-��kI�;'���J)n�:�D3��&��v艮���~L�����B`5�*�~*<�U���ؔ�'#�ؠ�ꣶ�ĵCa�Ejд���'YcC�4*'IQn�iRx2��u}ǐ2wrh�I��d���+h{��>�CK�m�y	�6�UvMs��ev:��r#��2(���<�͓�<y�'���[��5�O
�����ci�
Ҿ,������Hw�������Bp�uH��9��U�y͘�v��L�Z���r� ��E,����^�2���hv����k�����P����A�]&��K R��(���˔� j�3�q`w�-�=�`z�Hg��Y�~тO�!t�@x��,��]�:r�GG2BRj�x�� <\È�BiI�+��@ l��q��V��,<>�����t.얲:N����^�N�4*�d��CP�i|:�q��;���7c�ǜ����F���6_7������r:k���6�w8�Ngk�s�;����/�����_��up��S�;6 ��p٠�l�g"�5�k�u��F��Df�c���{l 6�`4�Y���Y�B$���~P�
ؾ���[�#�!�l$�R�&Id��I�EP�x�-eU*�T��z�`i���8��!�����8���و�ܯ�R:��8���)̒&q�a)����^Ȣu�x��u�UQ�C������Rc)ꠅEz'B��U�>���K���>�����@V�c�U'��q>��,7�u1r�Yn��,�"�a6��v��Z�x�U������,.�yl �M�4��A��	;k�Tqf�a��"��jMz�6��B!����g�0blxL�y߇Ԍ�Ӯ�(\�=0/"����d���ǓGy�̓/y����-c�t���]�IB�(#ڃԾA	9��j͡
&!���`�bJ�(%-��~Z7N1�5���V�۲O�c�����hĮ^� ��A��̙��+�B��ݗ�-��4��5Ul�?D��HGM���niTO�t�H���i�H�ܰu3G0$��H��\��}���b-�Sh$��X NG3��a99$����B1S����P���"��|�0��F|�f4�����sraz���ohkI~!�5 :N�(׳C (��rBH'%�86�[�A���a]���a��0�1�w`�aϴ��V6g5_*1��\p�@�y��x�, �k�>���4 ��R�Џ(��@m'���:�~��>���\��t	w%��3�y��`�Z/��e�> #��OUõ�,�H:�o����t�tp���� ��T�Qς�����$rF��,����,ZX&���R^h������bV}D� 1�3��Ԍ2׮
$��(֒K��<!�����&��rT$�eX�z[���rJn�=m�ur�+�V�����l�=-�w@J��SNc�C肎.��#��n��]s��X-�b˞��_VXJ��6�Q�8Z:Ղ��PjcN�j"&��活�v��m���G���X�t���)� �Y`��@����I�w���HV�s���~38+	X���P�f��I��<3�m�t���n_��w�|q�h�	�¸ġ�Ȉ���pq���+�3y��L�{E�N�c�~L>��<�,)p'��NQۤ�B����&�)�q�`��0��J,T,$K���D��W8@�Q#�9��� X��"�M���s�v��m����i~��W�����-���j28�#���IE��+o�� �g����ר�K���\2d��d�la��t@.w$8d��CTL��pz{a2� Nn��a�?��5�
�aM?��6��Ʊ���2AI�r��}K
�j�`䣚�0�����?_���u�|$��eš� ��9]�#��=���2�"X�.f��|q�H�-�cs��X�\�abr��JH��깆�y>���C�
]�Ft�`}�P:x�e��}��[
1�)DD���꣢�\��[��CvG�����c'�2M�v#]�]n0r���k�'o��������7�����5�҃���c�&y$3�#�7n�Q
@{ָ��?�r�t�5�4�F�e7r.r�V$��lv���cݍz�w��'��η�lW����3�6�����CF���i�_�p�mFH�C�x��o �l��4����I�DjƱ��)G�S@�| ������ ��t��u�L�sBsDql�;��w/僑y����6�i�C����O�{��r_E������9���s�t�H���!��*s�Kυ0b6������k=1�����
J}�Ec0ؤ���X�(�����*���
c9.y�x�������P�OSm�Ǔ��G�A���	u�Aj>e�Q����̫�@�Ax�$����B2�̛b��+y�|yԒ|O���Bǒ|H�w��B��_ZUUs+}E�>��,���p(X�������R����J�oJ� >�rVp+�ɀ!�z3��@ͼ���	53�}(�i������I�N�,�_�}6`3��.._��gaaTq�{aIi!XM�.-)ӟ��- �D�T�! ����i��H�g���]�a��ӷ����Q
`�r$4��.r��.3�����*��z�d�a`��3��
�s���t6���HG��N�Ig{�M��_$#��Wq�~���i|(J���rc�b0d���7����5P�	����i��^���0:sby�M�
���ꉈRf tB� W�\�������*�M(�huD�a|6�/����R���eƱ��B����f���Z�Q� =�����U�u�r�[q�>HQz07�6l�aI�:�7�1m�9�E�@���^���*�(w5[-���\?�v�j��Siw8� �Fg���çAD�����b@��͒�H- �R�������v�y)I0W�?*�m��B����v�񔤠"����6�S��"�q<}���D�:ȣ�M�������v����,�,Q�5OD��0��Bh���.��Ə�������/#9���s;Q��56�̣��5�$�R[@�9|�����wLn��ϑ���vDj}�
t?̦�!��@n�!h5"H�� 8@+n|K ��.���� V3V��#�q��-ƶ�M5`;�rU�P?��ר�h���gd� s/2$�4T�vAr�>�x���m�4S��t���n͠J�И!�1Mfڼ��W��#6
f�}�Z�� ��@^aG#3��Y��*0��*,��ě ��4��胍-��=�bf��yrk����wD#u�fV"�oV
8��
+���!��;a�8vK�F���1����J5:sɢzn�.���c�OZ��/�{ ��NG��a-��`�]��e�c�YE/[�4WU���\t�����镚���Up?�>iJ�/�9�������cφ��.�F�����l���޸��: ��p�U�����g�Mq�Z�Xn�ᮦ�L:�'�<4T������N��,Z�ROE��,�n��}L1�S�l/6 k��0��BX�)��A�)eBIAnH�l�r�ޭ�w(S�;�x��o� ����R&X�e� Y���<'X���q�q���
�/�E����~��5��D�s� ��+�>��V\�;���:O5~v�|��Y���.��f-�c7����J~���J�߯J,�*��_<�)�^�^���T�.�["UD:���z�>/ҏD����4_��D�/�~.Ҙ[�(6���V���'���ߖ�E�Y�ǫ��|�l��4���2�����PU}��e�܊r/,*��\}�g��%��c�T�{81�� ���?y(N�A���_�A\�ւ���$S�Ň=ę:-/f�B�(x
���U�@s���N�/�c*z!{#���bDq�BLc���X�����2b��
-��/g��mq�ʯO�c5P�H�;��t�-D�,6ƍ�0�/�QRXt² Ƞl?n���>ؗN���?N����w�����o�Л6�m8_�@5K��P "�
$6g��j
h�"C��q #��ش�¸�t���r�F<.fe�}��(J�8��U�.9��㠆ج�!t�al� �6� f�9!ˍb�g��/4g54g��,&~�T��`��3U�����K!���3Ũ���PR�`��?S ���X�gщd�u�+AHU�5��$J)H�mQ�����s�,�����{O�;m<Z�]�3Tt1�dAY��WY�'ޗ�Z(l����S�+X�0��Ȯ<�JW��ab���V+&�����x!K�H��ٕ,�
1V�e�,+��,^�.q�Į��D
���a�x*��sn*�0T�KjF{خ*r4�y�)Xr2��RiO>�I�m���d�,��<���n�$-�$gi  ��i�E���*���z��2瓠%&���=Jء�� va�
�9�6[��X&t����ljaP+YA�#5[��JvP���ƶ23�d�`�[X�JEP� �Z���¾ze�х	�T?������O~��*w�����%'1R�3�JD:Q��xA�j�S�`G2ܸ��{���v'ҳ�e0k�H�·7�����rփz� �݈G�{��cM�y���pY���{' Xi�r��u;Ї��<�*7�Mq�&H_�k�׌q����>��mG���4�O+��7�0������7t��vj/k))%��X�R�����k�[ý�8�{�n9`���̫*���/-).)���+&��۹�x���7l�������\U�}����qO3Ez�H��1�N���+D��H�E:����"��H���</R�H�%�/D:���y"�G���W}<�eCi�C|j�.��2C�������w��D����d��n��(c�Z(������B��L*[q5ؼ|����0n��zg�Z�2�-v��E��/�=�Ku����X9����朔�e
��D�c��b�^��:���lL���Ca-�S��D��oC���(�'���7#b�^P �Ѭ*�����Π��A5��j����լ6��v����G��6�ꦰ�4w���l�{Q�zW��cU�/�C���2��{ƪ|�9Q��� �����U��UO�hU/a��U��f����[k(��2�3�-�E���M�9��9f�����L�]�Ci/��r�Q�͔K��vHl@9�x���1Gch�%�Z�kY�\uN�}�S���v�(k�SȪ��LU�α�J� ��,�w�KRœ?�'����0(���>���=��(L��D?�m"�^D��RfJg".�n���wlA�[ؐ�0�I��|�����xl ��A}��>���Eq5p{�j�����7hF�Q���g?
�sʂ���z�"V5_,�(�kc�h��2S9��!�Q�f�/�=��}����������\�����Q^����B��wb����7�
�WT�,�µ"t�
����w83��YP%l;x��@pUP��VU��"ܯVP�ע��MeQ�����]pU|Z�
F[��I{�O���h���!�!5s�����8�91�6��>ش2����%�%��
�r|��Ar+�˪JpG�nO]�Js����!|����;n J�;�?h{�cuI��%��FOm������n��������T�۹sg�S �b�&�u\�pݳ2����������?7M�s��oY����_3O2�]��#��(��WV�9\��q�����~c:kh�+��o�e,rӼu�;h^w ��7&��M�zn- ��eH�,p�R����py�~��.���V����DqY�����	�6��mΖ���@8�(���C]�ms1�,R}��T^e@�߽�Ϸй2�|g�{�	�t�Dx�g�%���Jgװytd��')����F��G4���}��F�	Q~�G.㦉�����#ʫ��G�^}O�D�A��܃�P\M�k�J�Wʚ��D�%��{��n�J�lϽb��j�5[�ZE�E�Y�V~R�*?*]���W�^���]W\�:�Kp�W3\;�'
�l\�`�_��GઆK����#Hz#;��������OC5�ro\zQqye�<�
󡂀k^$	Q�"�*D�d�%�!*�x��
|^څ]��?����C|�E[��^*�ʆxZ �nlI�Ic�����k�'�u�YS^�
az�j�7A���Y�=�����O�]�V��?9�:7D�ˉ��Ca
"TP�+�!Cs�P԰0p!�p$x����1`�f��y˕r����f#��\���8V|�?:M�)�7ޠ6���r�����|k~i~�È������>��*'����H�ܨ��뇧91F��EH��+J�������գ���,l<T����_�,�/(
|����dnYX�f�!<ԫv�`C��m!`i��_c��c<��T��h�c4^���#Sq8Ory��'O��=�t�$~&�Z����WsK{��$���)9�e��Pet�0Ef=����
��/�l������W(דm+:�3��,���Eh|II�����z�ߴf��?:x:{	��|��܌8�ha����\=p톋-v�DH_�˱�-Z��OR��ρ�T������ƞy?��,�~�����R;��Mϯ*)�U&���t5��[�7Oi��.-Ba(� Xꡧ������F�!��D��˨BҚ���u
G,���YpO�� N:�x!f�G�������7^�=��}d \���(]+O�ƞ�8��޶�o;~1���@i��ϝpm�+�L�pni�I�`��~�,�[hHE�	(�P�f��|x���ŕG&g�y#هr�7z-����򏡕��c��Z�Q4y-ڬ���!n�Ni�C�cia�������� ��q=��f]C5�ڐ�1|?`Un~�"o���mp��qņ �V7$~Au���S��Ӭ<�!��.�sײG�ȺX�[�+��W��
�9}-����qye���ĖASۄc�%�a�q���H�+8�M��D��?�*��\fVO.�6�U�ޠ�yAJ��!�ou��'�,�~,�a^�����:=���
4}^��#�^,|b.���--�Wsq>���Ϝj����u�7�;�Pp��<���0��_=��4�>�E��H;Dzޣ<�/�D�.ҋ�id.�
ar%�y2�[���Q�IV�k�D�5T��Y�	�"ӡ5feX�ITc:��\�7T�2�lϗ����Sغ���a�8�7�a�zc�࿆<<kD��ó����Yc��óW�aOї	T�uT�a�O��Ĝ>�~Ne�O��M��L�Xg;1��p�����O�W�8���S��u�j���*UOƱ�P��@�I兾�"������eE<�=��(
B���Wb^�{�78�ڔ�Q�L�ļ�"����[��SaZC�S���q��)ćv��žz�ː�u\��Z'�$�t�H;D:�	�A��t�H��Y�c��"�$R���?��U�����j�_Rb(u;X�����ؿ��~d��\0e�9!+��z�_
�wcؚgB�#�!�F*k}P)RT8��!��>����'U�C�n�(���5-�e?�D.��H���װ9��-uN��T�}�$R����Κg��:'Ae4kŚ��V���;q��v���'��c��;�T;I#�X�s�"Ռ`��Z��n¡�	!�n�jBZ�p��u�d��攫�k����3��6w�s�l~[R�7�-	^K���GkR2���_����*����Ǖ����xc��9�gX��q�};�wf͞{�Z�򤎩ІR��4�Q�@���Vy��(Rg�%�hݲ�����s[!�@�Q_L��-�����=����Pp����5̰�[hi�ܷm�D{+�xu�;��/W��� j�@���W^{b���L~�N�S��[ �@j�]�0�K>���J�=�Hº�N��hə.���c�S�[�y ҈02m���:ĳS��tŁ�v(�.� ��"�Jn[}��Li��P��J�@h��r�yp����򽃿�$7����2�l���J-R�2->����4�VO�/�� �TU�-y�J�C��L�}E4s�-R�Kn�[x�&���B�Te�?꽸`l���@��nK �A�S��⻔v+�Kn�=kV�?v�9 ����w�+-m��u\ipjJ��{S����-��0i�S��P��w�Q|�'߇c�[zG~�9o�#s��K(�\mI�� ���] )y;�����V{��o�w����"W�*
Pwxj�w(p��ӵ������^Ĥ��S3�G����6�*r>�\���|C �)��_��/��493Xڅ�����1Z��|�w������_®�җ�G3��U�^�<x�n���\j���p����\��V+��n�m��8t�u�m�;�l�/��u݊7
��?K�� &�Xe��nV��o�ٔ��*u�/J{ʚPwL�}~�Ʒ #���q�� �cv\��ҋs�f�I�]�И��Ȟ�#7[{��_Dji����ٺc�f���_���a�-u%Nqˆ0�α����q0������1I����"?�_���H��Ƀ�Fioy��pZܨ�1MO��`�h��=��3���x�e���͉sŸ��㓤ni\b�-�{U��Di�M��L������.��,n��(J�;�3��gv!CT�q�䛱�~��_МRe_�s$��A�m�7?|�����q�#[��Q��Uix[V���/(��}�h��X��@,ڟ3�ŭ:��Sykr��>����r��� T%��&x�r� ��Ȓg�=�����<-��;�j�&��  �U�� (6&�nއ�~�>����T��I���`�}�0�Q[�`���iH��z�g�D[U�G�rRQ�>N���)$rmQeQgr3���P��r�K�8��9��H(ѽ����$Oc^�#�e0y���rR�*����	�VM����b��5���([>e�ގ�����2׸�<l���[~D`U�����yr6tc��Hu�?A��`�MJs��p�����=�VO��2�C�޶������a�my�[
��o�-�IW��	�	h�z:}�Z�,|�)'�'��*�+�e��[)���\�,Up�
�<�W��8Iq;�����{z�	̰W^@<��5*$��A=�P^5���ʨi��B��Ӫˑ�*��	�ꛗ% ����YU�4�e�^;c���_��W���U���@@��k��+���
��+ϋ$��Ԁ�8�YW�%���pz� 9�C���C'=Z`������==���j��!޿�F��۞�}>�g� R�^;�욷p�?Tޯ[��|�TNJK��!nU��A��/?� ��"�،�|�Wn�`���e�M5n�K�j�¬ ��h�f�.�S��C�tP���Z��0Ԭ]v�B�z��#�8O?����6{��ϪL�"��Y��|Z����y
ӳeF�@�d!q�/@�=y�	yy��� s\�1G��l<��q~w�-�f^��(H����[>����y���X�y����y?�Ō#ܺQӨ8��
�������h�K�ϩ�������i��иf��F74IP���h$4�8$�Tj��ވl�Z�4�h�%���m��4�s���0���]�����M�Q���:Q���]�ůc�>�Z��]9R��Ϻy�^�z���ȏ�����`����Km<R//}F05�D���/���$Zt|��E���_�p��1%��g_&�������� ���Ί=Od#�Jd�s^�Xp6�'?�c��6_�>�&_�Cx>	��4·��Y`���]���m\��]����>�^hہm?�L�����~܅m����6���P�y�K�F��[J ��iC�_ڢ�o�EP#��m"��]�Eu��e ނ<m�����������>�~X�!?i�d�2���)���
��!�������ڨ�C��߻�:兗�����O#�RwT~�Ҭ�-�I���~�wSw���P��ȟd,h�1��1�}���� X=��q�$��/ih��X���n�+�`,��@����[�J�iِ�7��I6�L��3}爗�6|�m�F�l�����<V��%�v�|����nk/�e�줗��K�F���hn����'@8|�Y�O=r\�:�+�[��=����n"��/�E�vH�קf�\����
h��qN��Y���B����5P�H�r�"��֐�ō!�3p�R�Q�z��)�E����L<G��\`&�q���a�A��V9j\��@�!d��q��ނ&8��L�\6d�i�u�u;�7�o��l�ݍ�3
/X4�Z�ؠ ����@�l�7ɶ\@~�]��$/%��~{��6�c�l�X�$�٨w�[����.ne<��D�M�G��_4�Ojl�q{��K8�_��=�"��	6���߹���J_$�;06-$����Wk�~84T�o�\ж��'y�y苀A�|��%my?����Z�6Y7�li���ű��*�������w���4��M��R�Mڄ!gZ����?z�c�|?�mW�M�Ȯ]��g��@��	���,��B�xtj��H�U|?�mS��j��r=�������l�����m�<_:��
��d;��,w��������2L��8��j�S��H���	5�oCY+/CLeh���W(˂p�Sd�>�T;�o�(?��@�/���)ڿMt"�~�7�E�L�A�z՜�]�Vh�f��b��Hx�������X�'�|�=̝:ϱ,ź1k��{|�V:�6.u���
�}?%�}Y<5Ư��oI���~̵ʍ7���g�e�@�@�h���K��`g�_�����I��{�{�6yx�*��'7'����lQ�*����0��ޮR8�t."� �wJ��o�6Y��@���7��l���n�@"or��o���G\/"�$�l��5���"g7;E�aS�I
H�A�c�����.^7F��O�Qt��:��-���z�ޗQ���� un�Zp��/�v�0ɾn�L����z���#���Ҷ�Ŀ(���:A�ݓS�,{.�׽��#C�ݨ��P���N���Zu�^������!�Da6d] <�u�κ��6{?���v?�w����w;'�p���y]�%�_��|��u�}�끵�ao�S���z���&�k6?x=X�<�������ٸ�\�&q	��O[��VT ��v��o�'�6.q���Q&�-���8ɞ2ī����6��G ��o��AYH�`[���{�S��:�?
��.Mp����n�>z�k��?���11@�n�@��o��:ly�4�n�K������� E�^.̘��L"4��6�ʪ�Að�"�'�(����;����a�un�+���뛌��G�9"�B�K݋P�R��#TViY�kcK]w���~������u��Lg���V:[��S�N ��4�G�&Z(ԕ|��m�~�0�9s�2��'�]h��,̮U	�����n*�U����")s6�"��`��#�F�
34�H�h�X7V�O�w��o-�m{>��V2�X�Y�yoi�����~Q;T3J��(�}�� ��τZyjC{T�#�:q�'ѳ9X��{V{T�Fq3ӑ:�#�,�E���i(@#~8|��h-�*'4s�6e5��чi�D%�?� t���~
�����W� �޼W#��f��š��w�"E��[�O�(GU�\������G�\�R���a��˙������2X�[�3�xc&���ěl�y�mKf"�*��=`0Ϸ��e�9x�CW(����{�[�Y���?m:��6��@�{�I�_3����Q�ӽKƞ��	=g
�Q%�����5��y�Ǣ�7oԻI�hmub�7VF9��uiϟ��{/g���D��߂M-�٥#��M�wPִ���(�����77{N�]�􎀴� 5$����F7�Z��l=n��iEK�v�[8�mSK;�}��Gux'��[���~��f����E<Tn[��P�l\f�!�h��5�O���X��sq\^W�r�t\�u+�	-*z ���tD���i�a�Z
�����B\����k̓��il�<Y[.��^&�te�r��MiL~�۫ȗ?�c��ZP���@��&yg=��Bc2��l�n'�]�JX)���k�ZB��n��eb�\x���(����
��c<B�����=-�R|=�*i�kئ��9ʻZ��B��x0��T<q�/!�1�n�avK]���(��I�`/����VB�0��.��Jq����Z�8:.!�{-�I�:�k6�I#ٕ�a�ô�ټp���P�4�O��/��`6�7�����=�k��B���S%|�ݬ�����=ǹ���a�FN�X�]P��e�͜2M{�2�PyU�c�W���|�<VȪ]���U�����W\�&��r����R�tp�kϨ[�d�8h�ݎv2UM Pʶ�t���9V�o|\�_���Y�M+<-揓�C��hq��6�3�1�f?1�9�i��OWоQ���O�a����J �w��*�ģSW�8l��c���_���ޯ[��B�/�V��!�K�%H�w.����b���
4�Zo<@�@
�N�Z�E��V�k΂zg��đv����c(^?�K�DM���;��Cw������C~t�yA��}V���z�8ت�$m
���{8�'�Tew�JTv�h��W�����{�� [3�8�k"�D�Y�[���t�_�K��q�y����T@z��mS��1�> +��)ْf���\�o�����D��V�5�X��nڦ�Q;�R�+=r��$+�)�:�ۿ�%u�x�����_~�[E�F����ll�1n����j������Z��&����]?sA�sRIs��U�<�� �����\_� ����z���8o�_o�p�r��=`�3 2c��ǔ,�\�\�k�:���A�t� ���7�F/tx#2'��In&��j+d�'�|��6K�&�g�XR�C����H�2�6����iU
�9t�F�Ӿ�NrѠY�zנY�K�,�V�f��g�h���B�m�"�B��%�3P��H�׭���O���� ���/>�� �^\��D93����^?b�����A�����Oа���h�#��l���!�=Z��5�9�50-]�;�|�%1����j�k�F�-��9�G��-�C��%Z�"�:�.�u�g_�(���hU��L0�=]�m-_y��6��3�ׂx���{|	�\�#P ���g���u��d߫�n��c�s� ��C�@��M�t���.q3�a���$���EqrO���$��0�sl�{w����@/E︤��k�I�5�d�<��ɥ�cUh�y\#) X^أE����5n-<^* ��Q:}�p���9� L�}P�6t�E	�%ǣ��"G��R�#u�d�&�{(ڂ����pNF�wS��Z��s S~g�qg:q���y�GR�Vѻ������^��m܇s�ߠKF��K���%b��B����9�>�+|�E�^�_�뜩�؀弾K��W����E�P`�������m�Q'73R�0�m��hm��j��<㞼��<}z��5��N��]��˱�is1L��I]�&S�=�?���m d6�3c��������?q��m�*�*�?v�%�ѴJ��*�\>9p-��� ���@�w�XI�`z�5¡��=��C[���6f�`6��\/g���bz?�u�['�F���PJ��[���Kc��	�K�p.}�w�sr�:%��[�ve9_��uȥ������oPu�<�*����a��E����T�P��G��U��M	k��94*�ͮ�[P4�խK��z��r��C���^8�P:˓�h�Ѷ�F��ZYB��r���0/����-`�S����5�=RkK������nu�x~R�q<��`��V_�t�i$���`���F0{���1S>z�� �� ôA��MB�k+���=�+Q[�6z~�t��bY�����Wi�H�u1�X�]�y߸���|i�=s�u����kR�'D�=�5��ɓ��v��� n"�`�n�ɯ�|���8�GGm��CB���p��C"��ra��$��O<$J0�Շ$����`�14q�"��y[��v��w>�]��®n@W:0i�U��K�ĸ6��<���崈b�W�u�����F��	r���s�"��񨽁��?�����_�^��.�gG�ۣp�&�5d�Z��"��b�u��j:�ʍ5�&��'m�O�쟴���uK�s�������;��8i'��H��e;��*`��p���F�6�����نk�����6���ԝ%3�|m��u$�]{\��f4ָ��W��ё�΃����W��(O��o�왮�ͮ�{V4�h�<	/g��鍾'���Uʂ�p1�٭U^[mA���z`�V=�n�ԭ�.T�Ȃy]�_T~8	k1���ȑ���;����kv���r��/��U�+�Ke���>L��zY�z���<O<�4�VF��
Ş��b�8� ^�Wߺ���A@+�.eR��~������8����u2���^-�{Lg��!u	<�<�L��C����@��Fw�^�������q_�7T�a�1�&�Y�ʂ"!��MBZ!Nr�0���|ȅ#<Փj����mn屶��ē��y��<^�? d�����ø�GF�tq&���F=+Sl8m�t���.1���Vi.��k�Ig�X� iw��Q�u�-��F4~�e������O�d��hvO���Wa�mp��oյ�Ih1�r��垠vzp�]���<H�a�.�B�K�w�6�A}a���o�rX v�U_���w���8(W�A�>T��ݠ�ۿ���Ǧ�a=|�Y�6"-:{k�������-B)v��Q�o����;E=F�VnX��>DbB��G��>�!d!�ߌ��,Ho�(h)މk��\:u�߬���Kzi��{~�GΖv�-L�l�B�'K��9쇋OiߓЄ�'�ROdN�!���E��މ�ޘ�����V!�ѽ�G�~dѡ
�k����] A��*�y(���%i>7N��.I=�$bR�D��'F��]��;gѮ1�ܚ�4ʩ3�B���q���[���0����lY �7��8`@ʫ����yw����{����"���L�q#�=��Xo{\�#�=��ؠ����)��16�5Ɓ��4�aC�w�?��mF{[�!��;�%�}��qexK6X�P��w����"�V��S�?��������쏮���a���A��KQ�yX��y�c��i�����k�G�����.���'1������zS�PC�nn|���B�w�n���\vg4!���]5g�<ܦ�+R����Tw�p�i��ܭ8�Щ��Wt���ƃfw�}W����[u	�'�r�����T�A�A�q���u,�E�a��"�r4���V^��)��}�w��<���xZ20n�M�#���}z��ӟ������,P�kе��6u�n����u�g���k��!E�ׅ��"�ye�B�5>8�kǓ�:���}��߆�z+��q=R�᡽�X�͟p
����g�WI�&�a�2��'�?X7 +�E�Fr�<n)��b�\���xT�=�8��}�W��`FG� ��'uk[��sӧ���8�qh�8Q+?�ܼ�1>T�;�K�>��!�թ��YsO�B��w}��+��b�P6�x���"9;_K����@s���Iґvk]�O�#��:9����6i��]��|���}ƻ@�%t��xL�V��(����k��Z��V��V;�>�<�f �1�>[:Ҙ����T��jK`�*�y��U�^[�1ߑ l��@;HDk����X����ϸ4)���l�A��!��G%d"�/qE�_��?�8������%c蛸|c_q����L�ث�n�٣)Pr�R�����g�A��=���M�=w�.�c>?
,�8��ɟ�x�[.�.���� u7��[���a(�\�xJ�=J�f��Kאַ�YpIb��m�	
7@���n� �;a�[�)�ݫ��J�B�:�O�9$kq]J�-q"�{e0��|���Z|�HѦ�W2�
p0oeh��Q�w��<]�@!l��'����v=�N���}Jq�⪏4��\���Ylȭ���O���8^ǫ�gg�֣n[�/Z�$�]J����DQ�>�k�b�=��t�d���õ \�o��S�[�]�/�6[�S�6�cU�W�Z� ��la����L��W�0�R_?(�h�ܷg�,'��,K1ߑ�߃�8z^,��\쵓m��b)�����| �W�p�a?��~8x?��m��6lԆ��;�YU��q��6���i��3�vY�-��W��9�K�J��.�Üߪ�8���KN��Q�i��q��b:�~O"��j'=�W�������>ɠ����A�ڥÐ�݉~[R���N�L�)�?��Z8��a��n�Z�]���l�e�"��P���s�l\��E�Н룈c\q]�娥ZA��G)9#��Fk��(9)j�T^"�N'�e5�k����t�[�(tr'HUn����F�P�aV�2����u�[h���t?͎�:��F[�h�#�@�����e	��n�ڝ�߉�3:r���J ��=�F�����D���y�5�� 㗩��ˑfB�{�4@s�%��;��m�L��͟e���y�OLr�)�-IN����Y����ToR���9I��O�o��%H�3	\�aJ�((_W�ϖ�7V���%�P%��� ����/�Z�#h��R43ҵ��mt��_i�?�!m�r���Ĳ�]Kj�����J��pAF�JO�����ꏂ��b�ԫx�x�� DD��4��͉~����qf�)f�9�>�V[�;dy��Թ��9V�}R�{T�����)��,�}��h�;��#�U7���f=L 繓��h��a1�ט��c��?�����r�l���du4�ϴ�;�뀛݉~�ƛ���2n\7�ŝ��Qy[��u�Y��S���� �5�6ce�lW7lL[������o�����<��sn�L=R��7�C܈?����u�;R}�>+�ڴ����ѫ���5w��05�qN�E.�
����	�I�9l&�H2�a޸@@�۾zt�a�0Z?�:W��:y>Rg^�'٢}�B�L����|7g�Q|�6�k���^�i:��~�ް��?��x���U�"����"�ߨ)���x�t��k�.��I�tzo�qu�M��>��N�]�u?�O���Ӡzü4i���̻7�a��(��ι�{VC�Eĭ�	��z�֤G{�t;�U��=HȤ%[���o�@2k6�>��-_7�'hs -�UT�:���-7�I�5�CS�IN�TE4X������8ߋ�G�]ȓ��-���;���Q[yF��f d1���}�Y��gH1��h���7p�����l�����&lѦ���B�� ?�a��B���c��Q�b�������� -�+�E�����hW��L���ȡ�b�����`:v4�=DnX�Ĥ���������)Y呅h��sj�sJ:���E���1����%Y�&:���xs.-�z䇦e�6��#�HhS�9�א4k<t��2AR�F���s�?�G=^-t�#�x/ 3e_�w���Sc�_��P|���ʎ�k����%�o�d��X�l���m
��+u��:��dGi�|�qҥ�J?��<'
{$�8A�=�dlI�>C���NJ��˗���6s}�m�^=�����S=���v˲pinG�U��|2���������X{����q�3� �挊��[a�Z�g���+:
���B��3�)����>Rf���-�-ﵙ���Qj��ԧ�TZ���pҁ���s�g�^���[���˹���{���S�!��贶v�S�REw��_ �.
�j<Φ	�E~īw�r��r0K>9Up�Fƺz�xd5{b�E�5c���Gp�DQ�/rR�םX��������F��?"�Q�Ok�EO�Ώ�]*��E��:0�yh�A�R�Q>!�>7(�]��%6.���z/k���>��������:p�Ҟ몄خ�\C��mQ?��0�ZS��\̳�A)�Nf[�4(��@�ڊ?��Y�1\����J�@��<���EЌ@�)��л��/��|�|�;VF��Y2�v#�9{g;ù]���w��.�ב�L�-������Wj�T!�k���d9���%ŵ�)I%�Ax�:4��/��W�]�c��!�}��:�^)Y�N�����:�c����$�����<�Y�bC�~U��S����yf^�7IH�w۟F�7]��G���[�(������**�1��Wٝ�+�)�y��0���;�n��XQ��P�ׯP�ڠ�	��6!��/Nq�8�i�2ے_�YN��t�����f_K�_,\
��#k�t��>h-�q�;0�OQG�����˄%wO�S�Ԣ%�I��?�����k!����}��̡�Z��e�t/'0ZdV��x��<�?DrG�G�YB�pf�j}��;�K�P���O�z�D�$�}���c�ɩ��Nx��Y�����{�c��������&B��Z��������8c��P�E�w?���_$f�	�\#bE�y�
�G�yo� ��2��|b��彾�6*�a�'��p��s/©��^�֙���o}g�|�ɩp,����;��C͟j�)S�0���jֿ���Q߷�0�DOQ��r��Q��1�EB�J���1�L9,.6yG���6(S0;�Hj+�fq�ӶP��%B!;ЮB�X7�1���Y����}S��i�4�vN�8���ʅ�����}y�%%o��xW��A��V+���}d�l;O�l+gE�~BJ�hTn�E��N�jѹ��C�2,�>���a�F�2s8F�ڢ��!0��"fcY��#4��(
�/qWB�D�T�������Q*�t�B*�R!k���h,��\HNܶl��SGw�q!��^�C6�!CZ���3�2�O���9S���v��\l�v]�~�dME����[�wY�íw����++R���(X�_*�[ym�B3�b�%b�|��F�+��x����0�|U��O|�r���]�8���pYQ�������b��'Z:��!�eJ�v���ke�0Y�{�R�52{�ȩ��G�O�>Z<[�F&-�MG���K��7I뀃ӹ^��Y�]��V���¨`�_U�,��M����s,����M�p���⯇��oP����Aޠo&b���S��"q��C2�%���;��6i��>9L.zy<mǟ"Y]`M�T�����,r�>�q�q�I  Uo��z�r�՟(��W+UB��2�(4Nv�S?�D
Κ�����A�:ˁ���[�{�
��J�YN�k z�ÔwDR�X/�*\@>4j�(�[�WF4++{�.��l��ܾ2�4�c�/��Y���x�S�����2���huT�_0l��N�zgL �)1g<�7��!�CD���r�ԫ6dm/��f�ÍV���x����o�&��td��m��7֢�V�cG�'n�o�o0�>i�Ǉؗ�B�`"��lb�lV�%�����n�;˰�t��E�X�є}�q����"�a���v"t���r��o�����XA���;�|�&�I�1m�������Ht��7���$���Ї�{�ߧ�{�Z�]�wk���!��8}V���sC���dnbR�Z�c-��-'�����ċ�96���!���*�V9'�=��j��d��ߕT�JH�O��Ol*����z�U���B�ɒ�+�\5��𙨕)�ѽ�1�/M�dV��&h�pJ����1��C�
;&S	��jA��E)B�^�ͺ]�ͭ7o@�,������g��Ffד�(kv��w�e�+L�Y����JX[�dmT�x�ڨ�V�e;�o�P~��Y�s�-Xt��o/ݻHXeпv�}|n�����K�vXzr_f�b�t�<��8'���q<�n��¿+D��>W\����\�!�o����fټ�<yT%��P�[�R�kt#���;���������D�Uv���%�UϦ-@}�D����K3u���]��E��)yX"ۆ�k��Ò�J(���7{��J��F�L����d�QI>X2�XV�{ ��!%�I �}VP��m�˸���iH�o`�XQ&����E]9��'�����G*M�.��#]�$�.���d1̊�?�x'�Y��ǖ$��hLr�$X_�&7b�8��s
MjU�:#
��H��I
��Vk����1T��g�n�ݵ��~���������-wo�By�{a>pA�y�ԛU�ԗ��En Y���A�ekL�es�Ɩ�.|��w�`���H�\	o�9�"�C���wQ������8�VP��-��)$3a��~�������y���8�[9�-�a;1�ulNG�{(���S��񛧢�=�Gh�c��b|�����4���1�*����L�,�ٽ��"��U=$Ck��"�vx��Z�Yj��h$Iy��@�-���.-��m-g%�DᇄHנP!��	n�t��I�.��(~PI�����Q ��^���K��u��x�1Xn��zi���	5�n\����)��k�签+y���J�G���C&�'�	]�H�p��;_Ƅ+0�9-�o�P����i�Scy~���%������҇�pn��C��I��_��jH��
�jFv&�R��C�}GM�S꨷�}��D�H>�*��Ek�f�s�Kآ�S�$��1�*�������Z�>��+{#�-2��a�j�y�Q�V�5:��h`�V#�gi�'�5���sqz�~_�Я�9��y)�6���Cd!���R��bi���=]:�>�7�䠆�Y,ߢsO�F���2�h�@�r��s�)Č!�H�!���4��87߀�:C�:�>JX�]vsT�ux��S�@��y㹆uZ_6��4�2{-�^���7"P���%i`�Ǧ���n{g8]�4}f��&9O��M�d8�ZH�V��NT����9�2r��C�������3��pݿ$T(�5oI\�r�dP��^�����)/B�O�n��d��>�G;��,����Z�,IT�%L8$3I���.��b3�)�:��-G�4�2K����3���A����Ђ��:Q�X���]a푱������(}9�;-`����)y�!�g(�2GɚIV��e�H�#i��<���tu��y�2��>�ϰ�n�l��rJ��\(�Tv�+Yij�^���J�'����j�6Y
��݈�$�ia�FXP�@ ��!�s��Nъ��d���7ڑ�g�z�yOQ���.1�Ffgo"���eI�`�^#��S'�{��'�#5��^6��jts���5㽱/�`��W��4M>`Z8��rw�� l�ֳ&�4��Z���v���4�&�15����V ����y'��Y��ri��sR�;��A��%OK$w�� �R0冭P&,ՠ�����t����#3�ݴ$_���ռO��֯z��7��-��>���X5�x�e��)�3����vL�ˑ�%tK����_���Ucϡ�a}Ì.��������Ffh��e���l\8�߬$�r��$j<�z���K���B�2�Kx0������X$��d�/�e&�ھ�-Fzz�>j��z�CeQ��)�?h����>v����+1�[	�_���ބ��o�e}�	m�{0��<�q䰧�I \���$C*�ų���=����)�S���Km�g�d�w���w!��3!���_�/�I�>ƾ$�_�zc��$��U���U΍��Ȱ�������>�2�~}���_�N�9�-�2c�������(2������7����N�#cy���V���2��ɔE�}�E.��-m�M_ �N4\ _�6����� �mg�.��g�7�I�y��רNw6��~�N�T�˾��m,a�(a�,�*S/A�����`���L�=ʘ���&;)�aE���P,="
P �X~]�-�;N�ܺ'��@Y��i�W�\m�������Bq���k�9�QR35b�#D4��=>w֜����R�E"��<
���G���̎���� N$n��D��D����:����$$�p�N������'C�+�^Is���T�4J�ڲY~剙�LB��<�j��3�?���c��e�ni>�ֺ�����:SS�@�
�%OфAO�vK΋��nk�Xr��l�t8��a�"��d�F�B����&oV{)�<�>��ʶ����iv�=�
o��[i�N'�(��l72נ%�(vd��(ޝ�:8;~5s�qn�c�PU�� �2~8�����*�������ȓ��
��+��|ɗ<m���ԕ��Ҫ�F�-ã�,��%�r�⪅f��y;-�k9���l���'Kf��a����ʓ�>S��TH�V�6�8�T/V�Xg��z� \K{}���ό �fA���M�jx,nި*�����*����$ͤv׍�T@^�=轖Mތ���ԡAo|x��v	��E�a��Q��z�Z�hr�.uD�
��+��5��];��b`
�DlZ�)ou&Ѣ���a�⚌�*��-���V�g���zU��x1�PZE��3;Q�=3+K�Q�jؕ�bjXD+��$�6�DRޑ�z����%���g��v&<fx��s^4ybܬ�.�f��g[3HX*����Ӎ��3WH����v�mg�`�zGxȢg*o�7���j�u���ڙ=1$6���83���A�h���dfr���5�,J4#��m�3+^ޞ�6?�^��Ĩ���4}5��b����<z�ڣ����$Q̒�A�ud-p]�?aGq�EW�VB�D��8 ���pÝȭ��i��jᮀ6�U����^Kvw��4�6N���Z�n�к����x 2�O��:��$��a68}K{Jޱ*��� ��t�=�O��#h���M��&���0�^���^+��B�X!WɁ��:/�{'�hF�+�%���\Qا��������J?�������܂Uȿ�k��%3Ը� C�@,���I��:]c(�H��L~�?�q����Z��kY�3N�}���Z�РH�]>�^,'�#�R4���v�A)O����E�P�[1_+�g����h���c�ʠ�]�b=��������9^��-��`9��[�`X��+��q=�Dvc=��#�qO�zT$��!�����k�8IZr�o�kn��[�^�v֮0�O���d@�" ��r�/�`{�BB�����:�f�4xDr�d��Kk���o�w~������%�����P��H�t��^ã�0T� Ʊ�� �`��0-F�{3qr!n9,^bF�'PJ��x*���o�se�\�{"�"���Z�_�!�|�ů�%|m¯��+����aq9�֨g��oHcF�¶9F]�y��,i�T �Jz8Ώl)_�Rh��T�i�@�*I�M�5��fOl�~OG����P��΄_Ŷ'����-E*�8OA+o�)Q�J��� Z���)*�e(!nPK�n�X<�O��0�^r��o,���v�eCZUM�-�>�mG���im����A5����/�$���F�E�!S�bQT!zW����q��\��p���7^ E!�\>pa�͵[ry����s#�^�2]�������t�����В��w�+w���=�A�c?�;BN��>G;��N1�"m8%����l��o���~�vo�EN�;E��f�����C��u��x�U��0N�V<�<�E�ϭJ��U��F�z�p3� H����P�#��v��#P�r�Ć��HC,;����}_꯶uQ���1	 %n�pvuwS8K͎u��E��H�W�|E��߅�%����e	5�U�U-�A��hn�0]�U��Q(���VȄ`��J<
@{�m����zG�tu��x�=6�nt��++0��Z���I��A���h!�����"6�\i�l
�jeH�$���]T>T-K&ʇ�Տ� ����܈v|;O�4co7p�� p�"V�{\��l��l�r��9�t��t�-�f�X�e�>_biI����	tM��ٌ}�M��؞l�
Ǫy~�����v:�FЧ��E;+5�?Ȟ��Ao�jf{iY4s�`Uy�ڈ��`���{v�A	��gkXO�vG,��Z��b.C����k��n�"�v�p�qxD��5�������g{>:�2�)��R��S����=4:����}�C���0�����fՒ;�!8)�!��B���*��|��ܗ�"f� ����ܕ��W�$'�vD��-l��N�:8�O;9�u�<����&����.���P�t�a����N<����e��HG��v��bP��=�l�}!rF3���XU63�W/I&�ǌ�JW�ƭ߳� öS��Q'ET��Qm1�#�G���ex-c��oЁ�2H����`f��!B)��S��
YTz�:+�Q�(�ӏ2�/�(������1�B���'��O��1v:ƺ�8�����<&ބ`L�Nm�D��2��?ҠΒ	�(@�q�
��1�>���0�"m��J�=�CM�˂N�ڂ'o��s�����"a`�|B�Z9m(����c�U���R��"�%n����N��Uv%	s�I��j�s+�8�Fc�.nV���`�0ƻT�	�w����������ǌ�Ut�����1��|V��w%�ivn.�@�a��j�N��}��2����ed�ɜ��nG|1�֞���`��'��h�x!�
�A��NsX��������d���	ڂ��Y_�!���p���k��+���{�!��rW"���پ��-st~���W4��'����IR`"t:Ş���Z��$���� T0��i�e8\�>ƞE	U�1�J�%��/��D�D�LؙZ�����]��2���-�=�z�S8�}�L��Q$��Z��⛌�����0�/��1b14��^Q�4,�T_�Z
���3��F�[8,q��ɱ�Y#I���so7=����t/T� ĉ�T� L��}˪�5�{��!�S�t��^�S{>&�����&�����IC��>�/�o'��!���%�)�	�вu������j��5^����6}�`��,n5��;��b|�e1��-�q�ލ������ُ�ܝ�Wٽ���MQ���#��5��P�A�9L�C����P����%\� �0��B��HU��
cQ���W��Ke�7�п��̕��q�9É��㈴펭��/��	�����6�U�r�A]�Kܶ��b\���^�,���y"ي�I|�3�����}N�+U��D$��Ƚ0�8|�K*m��NX�����QC$�F���3��.��y2�e���y"(��T&[r�����9p,xb7��+�98Y��+L�p���U�����mo b���jd\m����ȼ��c !�̀F�5,�a@c�R�E�;�~jDac���PkS����X���-<�f/+c��_�j�9U@x�(G�(O�Z�FS2@�E��J�O��H���c��=<Y3�FY7H;IW���ih^5��]��h�m�dl杽�~���v�fh�s�BC���Q�ּ���ƍm��X�����R���(�ְU�R�"J�i�$ަ�`�>hِ�]LGm�l�+���+go��
L0@���&�)oRx?��W�l.68�J}9��N�i���n2�LH�C��ך�I���ƴ}�6��>�NKK�d�������5�_��Cܭ��-�n�6�]�xu�7���u�,KO�M�,y��W
D��N���4�F?�}�0�)\��i4f_��W��g{� V�Y9�X�ar�w ԧ*�k�栒��l �\*��H*~�Z|R�=� .ԏ��JU�D�'�g7�rT��MF�y�@c+�C3LDj���!E@"k����7 ~#�7U�0�~�����,�^���;�����W��+��񻲪��㌆6V��*B(1�78��b�*����!�"�Ky���n(lՓX�.�yTЃ"�@�V��1t���ͼ����R09���s!~�>g�� �.B{c)k7-r(F���L�@��9��t�x'?�ߎ����Z���4���h� �[��e���4h�u#���4�A������e E��o����~$�x�J��s�8|�!�`^~��'I \aV���� 8��T@�(v&�2�<w���]��R�(���:���k�Ų���&I+�<.�����a{�,Ch���`�W��\U^|j����AV�(+%A�0�F�K���+�^u߂����{_����K�Х k��庬�0F_��k��iD���W����v�8 o�~O~o�� ����3��=�S�s#�������Gį���޿�J�{3���&\�mhiD��Ff�R��oIj83�E~�S����I�65��1Q]z��)�$v�A��TC,�9D=�/�Tr	�2�O�h��5 ���GS�!��Aá��4��M���JK0"#��3"��#�bD�"j���K�`4��qO�hq���T\�v#���Ur;���ϖ��,�l8��{����@�����fW��5�#�n%����U��rܠ_NH���7o(�s7��>���@�_Cy:���N�����1��c/C�S5��[<�*:�ۯռ��m������1��\�\\�I�H�2]�����|�'K����;�*Y)�qƉ�G�(��� �<&�Aa�o4��s{�-�+}�k���\���[:��}�m�e+Y.��k�)y&�;��d���
�I�O�8��J�ڈ
E�*���-OF3���TG�ǆI��O����l.j�@ɚ��<-8#0tf�Ĺ��áP�¥��#xM���v:��� �/�~�� 2��chh����>��O��2s۫4f��=�fT�u�pN��X���5�`��4/F�}����"k�i�o���d���;9S����'e.*�ə�����}(dZM:}��YM6}�!]͞=��P��R	5$�0z�	LN̖ꃨ��i��[U^�����A�����H������]��<gۙf��G��e�s��.D_�eO2�?�&�z�"k��d�ga�D0���~�ܝy'?w������ox>�����F�o�#���/<f���q"Ko5P��l ��}\?\������#�K��?�3��CJ�� �=ߟ�����7��y\�~��~��sNNKO�E~�m�PQ�����qۑ|8l��[
K�ڊ�'y�G��n�(ID��(�����,mc�ކ�c*%`X�[��~�a����!�S"l@%���tkt2�g¥ f��#̇����ue̊�9v'�Q�1�B�0�47
���+!�����Ӷ��N�2�m
4��/*@��w6���ra��3H��׋���'����R��r�:h��f��o��^M?cJ����?����Zs�sg��%��:��F�)Aӵ���_��N0��ѯ2�H%>�,,�mE��P�͕�A)/�H>��C���p.ǭ7�dt
�P������	DINLa���'���`��0C��b�,{���_V��9�ו�Qhz�T@����\��ﮌ}X�����5������}������cQn9�v�,��o<8Af�f7����5�[�a�[V�:U����$M�l�mڊ�-�x{,T����p�VA�=[��P����YFi�;o��wN��N���p�i;���wy<�UC�ǰ{�Ȳ�V���m4y0�n?�7�����:���m���M�:��M�uo����x�rx;z!�����]�e�IcG.+��Y�������;� +�~�{EҋC^�U��5<�b�k�|?�a%;�_�{G��j��R˪�t��]���N�]�(�+z���N��˹RiX|���Q�FyO	s����AH��ZU6�$2��G� �}U���Փ�K=�<��?��� �c���̅�<-ݤ�ae=�t 2ߑ= ��P�C�0'v,>�i����"��Z���֮��w��-�꒧�����PVC�].�x�խ��_�^��ݱ���}����"t|�!���Q�͠X�q�R�ĝ+�#פ��1�!Р-�(?�w�<9l��#������#⡵�G�K��1���z����L�4��)P�Z�)U��~GɓD!��V7����S�@K�kO$�` �EO�^��"�a-�AMњv��ӓ-XF��ԡ)+ݛ`��>E�J\�h�K�8���2�5,c{[�+�w�ܾi(>��wŖ����9�۽M��n+�; �T�.�)����R��ց�H�E�܁���߹b,�z�f����.ka+�%����������\R��Q%&{Ҽ�^ qx�w��B��G,��8���0��p��^�� ��V|@\S,4f�`�� N$���QZp)��s� G��^lbU��]s��ʧ��_su��8��D�P����D黦��8](�ˉ��{�C�
����3m���S���)��v�r��^vW�H���6�]���zn��< &�@�)��3�� 5�O̩�x�G`\�pZ�ù�,�f�Nu��鎦_[�52����O~��Gu����/H���������.�v9��=eC�!JgU�TQw��xI���N2u"�8p�Di,Z�V8D��x�x����<����q��{rX��4�m�_�@��_/��1�O���۽��=��ⶣ��?!.0|�iU ���[��iw-����J���j��s�E���R)�W����M�Z
J@��W�j�vfٹ�$�(�k��e��@))ʊ��EY%I�Zo���]<���@�ǵ�-x�#� �āp�(2�bj�yE�0��KZ̫�qk�e,[A���-��o6^�S�k���q(o���#�y-6�E�օ%׈%%�fmz��$;Ť�p=@�����ƞ?d�d!v��Xԃ?�J�e|ܠ�>J�
�L��d��|t�2wCHX��b�$�װ��y����᜼���X=���t�D;�gvI6Ơ�~ òFS�H�6ԇ�� P���u�-�y� ��/�����̹��,�fK�=��{d�-�D����@\j�����i��q=��2�g
����h�t5a���A9UX�
�C8l����믞>[�,��WE�m�I�h{�=�`���6�8��a��A|�;䍀��'��B:#K't� K�Q���I(��� Y�I)����#�x�Ѷ��P��e�S�N��S{���閶�6����4�)ʫNuX���:KͰ m�cE_�Q/�*A�!Bw��Y��;���եo��A�"�مT�j�lFf�R'����;5�V땩�� ��[mn5?���	���i����Q��)<����]��9E^�xY�  fhH�������3��g���w��k��}� h�T'4�l�)� $䧻�3�x'�H�5�N��"�m��4����.�5���Z�8��5В���	���o���|����>0d܏�Z3x�ښ�M������}{[d=�3�j:z8�ig�)�jy��P�CՉ�宑<��3;	���d�ܦ	d�C+����Z�҇sI���\�g�X޸�c�qͰq��8Z�M�MЈ5%��_�Oʸ?/��������<�p�)Yl�m��2,�5h6��w��Wr����U[A�!{�ؔ��Z��5(��S�m�)/C�<�&uZ�ӑ��\�7H%�j������}�0�#G�m9{�:�k����5� �S��o�[���&חdV����;�J���7q�b���a�>���Tʭ��P=�}r3��͡^���v��utD�n@ͩ?��D�GdcI&��#4c!�ã�M �:/� 3�"��\�wS$n�	��C�!�!޶G��9�[�(�c���b��5opX¶C"�ۧ%R��5�m�C2�L��%�%I�h)�9�!]������w;�������ߠQ(V�;���(7�(^���t���s��W�k77{���vp��|�ݬPd�q��C�ʻ�xm�ςc���p�~��6�:�^���J�+�L�Fq~KFG�m6�~�[�9M8�ͣ�`ײ�vq'�����pa�D��ۖ�6�c�>����[��Z�6�$��JG�1 T2V��h^��;`���t��:O	�.6�V�.��\!2ߖ�a�ȼ]o�f��RmLg��f I��ҜTڛ�4���~/-��zٺ��*���=���p�������м��k���5j9u���T�Īj�����e�e�:n�ȸfF�1��Ǆ���z��}qֺ�1�Z4x4�cl=*��� �#�����3����������ʺT%��(�������}7 }����?{P.�UH��zB�B��Ʃ���7���V��[�*Am�v��~��z.�p��v:�.�[�xk�����m:��/>`��\�%��xC�W�x�W	���6�1ʦB[�m�.6�.�*4��yMX��|���$�(�vO��6w�7�!�e�:.�0�i��R�o}�ש`�q�OA9-q8�s�
��J��5���\.�=2�_���-Ŋ'M�yf����I�+�"(t{|#?�B�W^���@J�@o�Id���bk��ב�C�[�X�"������m\��.>�o���o	l��1�@���ocJ�p~rT||����N�"5��x�it�.�k*�=��O���W-���N3?v���\��B=iB(譼7�x��Ԡi��]�Z/�#��3��F�k�vt�ߎ��7q"��Ռ�ꎤ,�kd��񆍈�щ�Q�(q�TtȾ�u����W����a��`
��q�;O3���I=��z�!��(��~j�]]�k0uG�*���'cߵ�EfL�&U�n�lTU�0�D5y�S�V�8.�x��r�ؓ�Y�Է}ʱdok�{��)�VRF���������������0�
>pp��8�4|-��xt,�⒧���`b:�:�I4��h�jPj�@�t͉NTvc|Vm]]������*�i��)Z��mR�`nBU�j�pB6��k���hM3� ���'�1�V��Q�%�ZU�u�ɰ�z�9���@M���TM4�Ó��~o�����YE$C"�#�8�a5ok������+�{�m���#�����$s�,�,.�? eu-NP[��p�� g��>�b�E%�]B!�9B:�M�Tw�i9����{~[��:�v��#7"���{��n�.N�@_�5�tw�_q��s��tT�v�Yt���lPؾ�������W���۔�I��Qt�d�AF�����\�ZY��Qh6)"��b��,��W���AO-�`��!/dp�8�������/�k'8�����-}���c�5u�mUFi���cf�1pS �<��ڡ��d�MG���f��dc�s�U����ӕ�	c�sb��N��Efb�u�i �� [HP�$��]�-���y��]�.�nŨ�yTĽ��[���(+��K��[�=�Q?r)�gR_۶�u�
�d�bk�
�b�����d��O+^����^ @[�q����[�Z#v�e�w��Q� ��9t��\�����'1��xmJ��!.�!�����T/�o�]ca^���Fv��j!;T�:0��Eu�t`��fG&]	�ndGa�S?G�X����\
AM��{��"HQ�1V�"�/��a����-��D��D��f.gV#�o�%=�H#� �zV�Q"�Ï!v��e��"�w�f��P�S�l��V̲3�b*!{.)m����^���;8��`���sZ�s��`܆���8�*�5!sd���e�����Ճ�F��O7Z�}G�.6�B&�4�J.�s���^Q�v�j
[����z)��2��8̧��o�'�z�&O�f��`�A���ՅAtN�2z��^� �_��ۚ��:�?�tPePښ��d!ch�&=(��y�͑��8^�+S4��S��6z�hd#ｪz,6�؀�ҕ��&q�d�V�*�m
D)��po՟���kNy�lO��Y�٠,R�b�pOA��rV���V��a�fCϕ����V$^��C*=m���iC����^���iL�`G5��;n��w\�i�T����ts����A�� +��sF@�/`���d�o���E����H����p�\�[��.�4��5��k5����S�m[��l��V��K�i��K���Ͱ[n�"��37��4��;�{㐽^�Ӊ�n�_\��G�����2�
Ls�y���X(�C.$h���44�i|��Gb����cM�Q?�ǄϺ���&��&v��<��\v�2�E�"��߬ލjN%F�F�;���5��fA�ݿ�*�JB��n�֓ey+{&����6�އql{�β�!�	�e�9Ae�vD2@��K)��?�rҽ�$4Q���fC��\&��M�=>�2,h�Q>�Z�������^� ���d�7�=j�{Ft+�(y���HH埠(o���C?�2���D�VZ�UgK��f�U���~!X��Ό���?B��T��]?�AَˎD����mɿf�n�vtw��Qɒ)̗9����;��r`=�6fۙ���ա��zxo��]�w�ַ�n�GO��K�����SWI\���?�"��&���/��,�|��׭�U>>R��-�Q�� P��`� &/������qtE����ӷ�(�6��ԄHb�+�>,>�_p����q������0y�F��>`������>���
E�l$����uÒힸ�L�1��`jD[4_�'��(+y<�L�H#M�v��5��5��/��׭�$��6�-���䠥׺a�L�km;#?����H��lE����q4�P�/�>������ݐ<�^|ʻC	��%n����[�oT��
��}#3�vv��}`���7�Mއ�g�g�����>��Oeb���,����%����D�X��"�D��xU����WJ��;nm|
:�*�b�&@Ѽ��I�����{h�=�κf��!�9�^�� ,u�uE4<y���ղU�ф3�~���"a�P��c3R�����t$��m���8e4pL-Ys%���$Ά�TGL��'��aQY_a���\)O�\%{�--��,�-���;֕�&?����u�9��V�LN��_5Ojf�JN6v�|��?2�7�;���ކ07�R�8�H�A=��t�8��.�&�'Z�b�����D&�S�Ud&G��;A�ӎ|�ɺXM�|+-��6A��2�9C��r�P�'��=�
[ g�����ZR��Xj����W���m�}�y�Cz~�����3IW�+��x�><�!�����:��b<:��$_ퟨ�I�ד�ϙ�O�>g:d;ݳx��܅��3�-��}����;ˉ�o����Ҥ�dpn��㬬��zE�cHH��ER�g��j��ly ĭ��'��x"|�lc/����s9��/n�ޙ�>?���p�E�r��,ڇ�rC�>g�$q�o�G6�T+4�C���Y���V-������l)���yu��yK9ד�Z�RH�V�Yr{����)VbJ�:�̻�:Vj��SV.I��ˀ��)���fEQ�K���v񏅑%��M�2��G��u�������{�� 2���]k��c�9JW�1/�E� &�g���Ke��Ͻp��B*���%t�����C�a�$���*4�s�m9�\�G�J ?�A~��B80n�-$�������������h��_�oiW��>
�W\�;,�5߂�R��`�����!{�}�y,����@��1r6�g�י��с���\v���*J�sOCn���pC~jz������8b
�}�R�����Z�V>��}=����\�(�3��8�ۋ��I�"�|y��P�����h���W�vҁW��*)c�㙗�0Yg��(�+�c��x n��X�-�t��!J��:H��1�g:Y}Pm��q�4=D�D�J,�hvʕ)�o#\ֵ*��r��GgyG�;�7x�Xtz�Ri���y�l���&��6̹��s�V�=�O�&�kn_(@vttɒ�{��~7�h�e��gN<hXb_双,����:��)e�xUH�RF�VF3��r��M��ƣ:36��������K"�w�Ӥ�@��z�.^��7&) Fi�h~V����x]_T�L���2�t�)��̝O⚟�rP�2ݮ_-2s>�˒���/i/+����Ɛ����+*i)-�*�&�P�;U��?�j�R^4�n(*�"y��U����d�R���@F/�ռ�$}G��l���kڅ0Z����"�usAy=v�j������A{N�dV�u�\H%��/�8n�E��`q�eG��eU�9r���;�y{j���G�S��O[����&�/�����V�x�6����V�5��W�|w�2����Lnbh����g�����B����~����A��}l����ju�}_D�*��i@9����"�o.q��C�0�F5��N��>v@洅��
��Rl�EWL���%}��H������r�f\��@�����=E����P�K����Rih�(>Ց�(;\;H�Bh���b+�s�Nv�2~�l~Gd�;`��ྺ�O,w n"T.z��R�j��\lY����IP��0�|��MN�IsD��<�� m�>��a^�A��~G_�F�O�4�fzD�2^�*�Yd�*�H+��k{rS�B��A�吞`��|H��' �
���	�I���C�/M�	s ����yY�\���V���o.*��Z��12�_	+��ޓ�T}N���{��4��sB��wlj�7����]�V�i�ť�J\���n&@�S;N��*݌��v:DW��u��&���OB6I�6��.B�Yl>�H��W
�����_�@��-�^��
�]�S�W��ڎ���b�V7p��9j�B���{��a��~=�c-��5{���O����Ÿ�1�g]FN�t�Y�[�?�n�����
��W��9�f+���<`�=MQtt�@=l�G���W6@8�����Թ�2������B"��������sx4Do���~;Rv!h�E�ze�:�FlZJ��y�H5�� ��AI��T����U��D 8eZ��y��h��y�x�ϵ�F<���G�f��9��EZw*�w���VC�[#9D���Kk�8�@��᝻k=�4��;��F|Kŷ���m·.����o��p�Ėء����w��
�{~�����jV���ΰ����>U
�[��軗�eU�ڱ��a��XS�}�ڊW+�!�
����HC�%T��?��׳�pz��	��)p�OT4��ҧ��C��'jp�i����w�+��/s.����3o���XFtX��;���q=:�4�ˆ�Q���m�ZC���dO�ws��=Y�;!M��Bq���3g-塣s�p�/�H�3k�7W$�%b������dN��E�s_��y�֌yr��q﷕Pǈx�#&�^�8��X���?ǽp��EKZ��dy��-��Y���ų�OH1b�'���|H1t��Y�˴�0K�Ӽ�|���	fQ�G����wּ�������{��!��G���KR����L��U�%c�U���_�$}�
�H\�Û����ca���+�>�a��،ѳ�_6!����U �Y��"5�DB�c���\L"����!�g��So$�g~��|��ؠ��Y��x.�g&,�������ϟų�2��)��g���s�x�M<��S�����.�|F<��A+��'�����Sȟ�����g����@<�����y��Q�L.��;��)��R<ۮ��e���xF>��c��	�<+�]|��ϘluV� �}��}D�Ù����U���T��T4�f)z�:�f�����\(iѲ?��UJ�dV�?0w�0]����Z����4���6I41ױu�+=wA����6i��)������i�gI�6:$۰\��!|c����nK��c� ��8uc�+?7o�R���R��m2a�R�P3Q nBj�"�+��`�1K���n���p��s��4�ܯrc]#h�k�o��@�Bnq��A7�A6�^�AR�üXȈ�
�`JZ��C!g4�^�9�:�ȫ����M�w���Y�ӽ�_5WC�`�A�RXhm�eH���3zѬ9������<�u�cP��I�� J�����GS/z�9W�~��.1�D��� &��ోs����㘵�/[>~��%"�������u9PJz�!�c&~͆�k����9M
B�f����8g#��t爼&~�G�����s�*E÷z����>�@�	�/Z��/���W���icMl�r�f�]�����9o�C-c0gƂE�<�ҿ�s�Is![f�џoZF�c�����M�/�OD�����]�?40XG6��s,Z�0w���G%�=ơ�ϔ<�P�B�����t��d�P�4����f�'�M�?\׼��5{�{�q�����
<��s�6�ilZ�Y�����_:��^�h�o�b�Z㨳�ʖ���H�3$��T}K��?�gb��ϕ��9�d#H�-���Ͽ�EdHO������'3���u̐6>�BIא���R�ht(#��Z��{���0�hU,A{�_��Q׏��L<������?���p�0�$H�s�1�u8c���u5'8F
��-C�@��{_�G:1Z�ݑt<�6M
#�a�$�A$�<�?���?��������P�D�MS�Ջ�(�:�(�&�(CAD*�O�Q��lR�Fbi��dqx�x-Mf�]��U�u4J-(R��Ѧ ŉ��hU���v'k��0��w7��� λ^����xHA�`�W��`6��IV-֮�P��?qv6���LE��>�rEѯ��ӹ'���N��˹�?!��p�~O3����~��$��ZFF^��p�.�xe[�&��&o�6S�/h�Z�����^"q�`�X�p��{N�t�$�P+�idTh�y�8�C��m5��\�mY�WG���_� 5������Ǒ����ж���CܥU�TGu9Hyn���I>[������i�UQ�&�U�Atf�)��-���S5Y�9ϟ�oƂS��+ce'�ۗ���C�G(�j��yλZ�,=x��?�|h��~�Tw��9��"��}��e$�!٤�x��r���UWNFYɷ���=K�I��]}��k����M6�I���9�]̽z�.�����#0U�t��R�<^�F�ء�$y�b%�pK����{�;�V�a��5�6E(8�b�!e�#Q����?U�݉Vۈ-(@P�	v�w!U@n)>౬9�Ey�2����,�� �o�e~���_w�f�P2���f#����*֜�P-�sK��^���N���U��^%dvѭb>���^�@���D���X�.V�!y�C�z�)�;E��S<{$�s���������eH�.��O�\}|�oa��l淼qEW�n\E	�9k��E�s=��rF��7�����G����Ek�QA�r` ��`HO���i��tSNY͹��,*�,yz������5�$�>�\-P�!�&��/�2C��BU�Q��o����8�d���������R{��u�=v�7���\n��^b���I��Pc�k_Bk82E�]��������ډ�_�ξ}��ſ2�Q^���z��PuV�J��K}�R-�J�VKe(5u�1��<c����^�o�I����K�������鿗<g(-"d���(�>�����+�{���yo�Ђ�3���F��c�!g�`�
��_Q�E��x��25r���hExX<��>�+<'�֠�G�P�[=���W���~|E��5���r��C`��p<m�(�i���9�qw�}��`���Е%;Ϲؼ�Գ j�eEؤ	��!�|�Ĺ�}yV�PղXj V��S��ȇ�R��J���b����7�Dc,��l;�WV-{�2�6j���4x9�Z{���d����� �;��&wnC�t.<����w~We���)�s`7^��XG"zt�]%�x�Y�����K Z�FL�� Hn5w|�Tt<��n5������YS�EΊ7e�OWe���>�H|���_y�h�ˮ�OG�^��t�c?S�<=�{Z�ED`Z� �$��a�j�ѫ%���!�+G}�5����3|���N8rܢ�U7 c��=}�{�r:DZ)�����`H�����-O.V��A)��6i��לV�CԵ�:v�4JrJ���C-���?'�fH㥱�_�a-5N�4��k��_�s�!}�����J��t@���$Z��G����UX�� ��	.�+;!<޳��k���w �1 g�z���<��wLl.�W!XW7 ����!
�K��>9�����w���>�GO�A��9����9��s�Ĝ+:�s�R�s皚s�:�͹;��s�ɓ�{��Ϲ�7�9������+�s�h<��Ry�F *�t'd��uHO�E
�O9�.�o�K� �<�@�O�
;m�\6Y��QEh?'����j����
D����d��"Z�C�d��0y��a�R������5� =�ˠ���"JQ����C��$J�9ҠZ��?�6V`�5�i�0�����䉺|���2�ɺ��X��B���-��T��X�.�au!�Y��/@E��4p=+s�_��,���D�6	ڙCiq��l
/�o��P?���k!v0Ĳ9w�s��+8�[ȟ�5��9R��킍�y�@�Yq��ު�>n5� L�{��8�Ƭ������b'&<�u"�y�Aah��̎���ٿ��8c��
�Κ&�$t!�o�d6췭A+�U_#�S.g��Vt���b9'Do�����jK�6?O>fh8yR!l�%l��L3���f*�V��{@�Y7X��{)�X�q�n2l�3x��K���[�c�\z��I�Y�͢�6d��-�?���'��<��V�$��9��c���&>�m�}��w�EE�����Bݾ��R)�N�i��Hʇ���=Εr��"|�?>�n��%�S���g��~�nKIv�u<F ��¶�H�Dx�����4�ȇ�f{G�6��C�*(>x��W��L+{Jẉ��C9V('^-������Z�0'vƒ�o8��������(g{\��gp&^����Å(ٿ��F.��c����^���H�@X��W�CiYw[�<��X4{���k
����J��孲����KE��,��/IޤT�uU˜�%j�`z��`��ZS�,l�krt���;` ���?��ug<X��U�/���x�"��Yx�'�2��8�b�ϳ@1/(�C��E�j���*��&�TG��A��t���jaް�<����ba�'x�8;�N1�ֵf�"��a���<=�>�~����Y%��}{����2��|c��t��HҨ�S)O�T����IҖ'9I$�=��J��	��t�A�,���8�%.|��!�G�]��/P�l9�l��CP�����.�(��P%��� ��3Mp�s7����hX���Ͼ��p�:�Qs�����|��Ǿ� ���Ĉ-�1� 9)ӌ��Tc�m穕��txe��Lk�2;+x�X���J�V�Ub�Ӽ��X�_?2������F�SA�OS� L�QX�ϵ��D=s���!A��@5��� }�۸X���Va�a�)F?�X�ɵxS���0o����'�<�`Ꭱ��c�Ű>�N�%�����t �_�l�_`���c��l�o·���7��͓�o��}sq���x��{���+TI�G0������!&���!h��	��QY앸z����q����3�냤���������{����wWh�y����K׭�E��[B��'E���W`���#�ЮJ�~8�s�S,F#��糨g�z�����
,�X74;�3VM����$X�}{�w-|�s���`!����b{�\r��[�h&d$-yV��j�е�l1DrYje�Kb/Q�w�j١e����к�
+g���*�)<�����p�s�'Կ_����>b����A���w��������娅�o�!ؔ�s��-��.�~L���GW�OLRS'����hf��W����H� '&�Mр/}KcB����%�`t�p[l!��sNfO"��ü��35l�w����������?����ϓ�j��AN;����;�v�~ۆ��͟��?s�26�v��D�1}�1�y�^�;�Ѵ=?��{�f2KE_�����fh��n�*ԛ!g��ܶ[x���j�����/��p��8�{o��Ÿw�t�qת�VJ�5Q�XӴ��vN��c~�m�Ð.�*?�E���0�;�����R����m"��KX�l,�%���J6H�U��4��]���i�âpϼ�=ܺ�،��p�=�f�����s(I���' ?�B ��Zɬ���10�F��v����X�8�8� �]���z|���S�Wt��2��DcaH)�!qwZ!��N;elk�|ܗ�h�Fٶ�'=W�Pr������k��n�;�<�ƃ�+�uQ�՚���U�xd��.�KZ�v����[��5�b_�X�}�_�K�q�������B6�{ђ���ı��k#���Q=����u;��ꉼ"�E�����I<��s&�kvM�s|��sFV��lw����gVV� ����
�?s%Y���͛��%]���|�9K�4A������@�Y�Г�hA^�/���ᱤ<`��d¼�}z;���8�I���VV��������OD�� }n����E�z̚�9�Κ���"��7g�+����(*/J�X0�K��_�"�M[�w挦;���A8��7W;h�b��`�ED��+X�`�21u���O��H�7o�����+�K��y`/��>R<���]F,,�p��������w4�>4�)���������6呛`nu�f
4R'������)DÏ+��Hs_�"Y�E���4w/|g�85�>�yȩ�MmK��ZRȳ87�O�a�F����[�Y���6� -��H���R�4O*�fIwBL�!<B�C��χ�l�o� �uK�8B��̗�n�"������Ś�����߿��\4�����=_*u�j��U���/�7���]�JE�����������Q�����Qs��������ZQ��"\��rH����ʒ�zT�CH���TTdTTTԣ:&��GEF����Ϲ�\�������gݳǵ��{��Oe�S�q���ܤKhV?��%�����C�#�)L�*��P��&ռ��U�Wxǒ��2�T�ώ���I���п2��c_o��SZ�b׺o��[�+"(��u����Z�덥,��"��^�qI4�����iXK1OB�I*����������Y�J!+(�@J:I+t�8�����rF���<o};
�����&B�f�����}��t�>����˦+;8֭_�/-U��A�h����	UA�#,l��Lj��4�y����I�]�b�����c��}�O(o�J1�B�K�������XG��0�j�kJM�)�/�p���)5a��H�x�'���Y�-�p+|��7�ICE�۟b_��$�!��O�w�s��{u���:[��(�
3��
�������h��n�s�?f#��rP�X�_W>BY��n1�9G�W
��� b/r�K�����K�(Ñ�f.C�p`�Al;g't;�H�i�H!}�n!C���n!Bs�r#?͂���4�G�PP�ħ�KU�����2���A�²�X�Z��䤐\�g��)yB�����<�s�7�L��U���<,�TT��h0��BFkϺ�"t|�z߭^-�f>If������߭M|s���N��[ƞ�Rz��:͆�F�X��LcQ�m$�)��S�Ere2��7����� ��VRK�y"����},�G{��j���Yi1�}P|b�K���g�C���6K����ĳr����
���eSg�b��P�.�������/��E�QDn<嬡�W�D�ɻ��vB4������j_�N)� �j(��#�����r³��x�^M�/�O�]@[%�ĊN��p���cy�vJ?����u����c[�a��N6%C��?[z��.�A�g�K�"~�T��9�j�Jǻ��
x�����T�{���T^2�;v��賈c=�a50�P�%>|V���b�����z}[�hƅ!��1i���l�|һ{���-�e����^��l��m��ťD�?!�G��߷�n5�����Q_��ĥO:|T/�>Sճ����ݸ��P��N���d�������ǹ&d'�����ݎge���K
z ?���:^�N��ά���UZ�ѝ)�%��s��j�k'�AO҇;����󥕴I��'�d�l�n��h	O;��ă��fڕ@{,K�|����.K'�c](z�4��R<���Sw����p!������A��<�4G�P��O�K����H�Kfm����>}��v���=������C�"����p���Z�8�����eA|^(A��%��B`�ؑ )P�a�����q#��v
ɇK�*���M%�{��A5�q�n���!�p=�)��gm[�uݐ,=����>���_�������=�=��\��j#��ez�vi��mr\R(��i=��{X_?����	�I��X��"�d��f��n��Le߲���$H/z��
�%I��L�i���2��0��G��z�E�K��)m�Ϳ��1�H3~�Y:Oڧx�Ф�w*r	�Ͽ�/(���?�%��E6�� %��괻�������,�T�S��^�-[R��F���`�}͛&�����sl��6�S�~(O�c�����������}��
~���J�C�_�f�U1�8�RVv)��}�F��� }
S�����V��޿�w`Od�M�{���R㵿&oO�ơ�-��D��|U*'$�����)�o�HR=�����5dr9ƶs��H�w�#�n��k2�#fK3���L^Z��-/�.�����!Z'rZ�=��2b��Ap����Z��l���<�\5[z��i�w�+��t���F!R"o:i�:F��'Ɏ[
�b����"��j�T�GK�FKy�[Vw���O��/����f�ۥ$�.�%a}RSŤ��?����I�@�\ �~�c;��sm
�Cڅ�2ʘ[¶�[��n���7
��'&'Q�
�L�imgWEz�4ĮtP&������r�M�#�r�E9��P�hVF�<�.�~9No���ѫ���Ů3R*.�e��Q�A��%����XK-TQ�,r�v�/Hy��}��\�CJW"��/�ѵ[�
���ؘ�0�@*� e}l��z�~����֙�NrG?B�H3�0"�G�]�Y�<ͅT�0r����,KB*�X�C�WT��������yEi�A�JG��a,!GSr�t9��e�Ќ8T��%nf��jȫ�YU2�����WQ.e�)���l�[�t$O��Rͮ�m<�5*��"q�ȿ	~�Y��[z�Yy��E�&I|��@��g����|�X`,�1�Ηe��͙�
�'��I��5+��%�?��g hT��f[��)4*SU#�P6�ʾ��f35�}�21I����v���oy��&��f/�T;�O�a�L��6�������{�wk5~��1*3�?YLS�9�9�#�j�%լK�_�T�.�q]R�l��[΍�뫽_a�¥��h�S�Q6{�db#gl���@Il�v�OtdR5�5�oN&y�����Ժ=,v�t�Jh�A�,8���a(IIJ_�":UE�I7�"��"�y�=GE��"�Q�T�_�����plY�m�=�Bؖñ�?+��\S��`��ʹ�%FA�4�S���KA����(��)���1
j9�Jim�H��ޓ�7W�/���Q麿�5�E%	�����H�s<�z�	�{y;�[ԗ���k��&'⑇�Q�J`�er�#i4�ͬ�3jR�^ ���Ra��Y/�=K��G�͞C3T~�����%�����w��?�z�0�o�[ɛC�aI����#�FgK�p����ͻ�����k(��l�Ȼ���+f�Z��3�߼���ӷ���|W�"�2��p�y�-�Ɇ��i�7�s1P{P-*��V��~y8�"���N��9b���	��r�1�Iީ�d5���蠷�^[P�Ը��AZ�����*y`J�n�~�	R�h)�%��q�:�A��k�u��]Gn�޴��N�G���u��Ó��=5e���n�������٭'�g`��2O}���9:�K�N�;��J�I�Vwv)��3p2$�_M����S��
��^���A/\
L���c�t�$���P�/Zrp�����Ӷ]e�%/Cj~����ǩ��A~�Ȣ���{�Ηkl���0����j��>��[کr_ϗ�z�e�Gn�꾪;|� ?Ϫn�6�?6D	xk?��x�'���A�ym5d��vieK���R$��=^��ney���,.}U�C�x�����7���,p�]�������\�
b���,ZkF@-j9��"O����jj���@�2��3�4��:�"�2T�>�M>���2g⫴��4�� ���\���������[�vߦj��ό���Oe�Зo���̍��פF�"3�z���'��Ef�x�w��|�Z.�3.f1����煬��U�/$��Z�Y�V#S��F'��Y���k9T�)z_��8���l���5��t�0���,Ej�u� Vo����}s��'*h���F8�l��K�n��� ��s^�&��+z�	�-��~��>Y\��]�~�/EǓ��	A�L���'}R��i�qAp�k� ؛���կs����a�7x�%��h_I!���P�{7�[t'��/�p�r���5�Gw������R��'ӿ���G�u݌�uI����a.��x�s��7TX.9�n���][tr�����:�I���>e�����ԣ~�
+mz��1=ArV���M0���l���m4i�㐛(� J6�%k-��Q�&�'�d�<�<J��Md��~�-�h]�v��ە��(��'���yxV�)d$��$4�	ͳ2�*��)~�����ƇT'�s"5t#�c�((�����$W݌o��<�z��,ոy�9��(3��}m��<1,��cW+�GrU�<��<�B�}i�L��ܤ�&N����W���1���ӹ?���8x[��R�|������[��]��z��࣏��ݱ�7��[Xc���w�nQ���7�wm�6[�:-���iS�<�>�}�۪O�>B���6��oRvH��k�����C����%K�$K׺>�Mr�tm�T����Z,�j�������Hʀ�J7���BZN�߄�sv>Ƚ�'h�WS�E��!�6�5q�1�M듚��	��Yƪ9�L��(�S�uՏ�͝���c�;}J!�a}R�t���fce"��a6RQH��~�X�:�`𓎛�>��h%��z��AT_���"���<�ce�Wb+wP���&(��,���
$8��>��cw1�u7��C�A�1j�g{��fJ�y'��[�>��"��>���Vy�\ˈ�I5<��"袎N����G���$CH@\z?1�s���
|�FBT}m*�|���B��.�G��+9�4�Q�:�aZ��l�Z�VɈ�>dAo{�H�d���\�Bժ��-N�OZ�w��^�\��4r���vK�.�Fq���S���4�W�����#T���}���w���o��i����z_�ޭ�ҕ/R�.�6n���w٬�U�|��AX�.��lE�~v[e�{�^D�=0ޤ7�;���1X��G�=��`�)+a��������ln�Ɋ�V����^��G��x��A^��Iſ$���\1�F�ΤT��$��]�W~K=P�t����wD��{����&)�	��J��ޮ1���_��W��?� $y��:_��=�����+���!�����\�T�T6�K���_����5�����'ӗ����v�l�*st~t�J��b|���rRU6G����E����9Y:�4xe�B����6�G���)������mYr_�8x����t��cu�{��9����6�\��Y�$�$���N_�0��A%	1+?�[y�oȦk����q�=�yWd��%1+�CWv��T�6��9ҝGhƮ��U�{`�i'��؆u���b��yy;�l������cwp��N�v��'�v1ݙ0䅩��b�6	C^�.��Pl\S�ܡ�Vr�́2m�K�X�@,�`������[x�w���z1�����^�\�+�~7�qhh�%<k'eIY�R�+�r�G�(�V�x��L_�ƴl�X��3�7d��yboB���*�R]�TG��#"@O�l��_0C�E^��Ny�S��3Q��Z����j��Ɛ4�0�F��#�=��
f��S�G�߼" ��+���#
t�0��Kx'</e*/�	"Q�z�(��8� �ՠ�N?Ie�*�f$%dT�.?˨�D����$*믐�{�Xr��N��c~yCܑ��Ώ���#�	���eO��!'�SD\G���Z "�����(*���FQ�3�<�ioE�F�y">��J(�9����!o��!uE=��o��_�vVޡ�,��d]c1�||��Nc�����v�˾������;d�,�G�|��;��j�<.�d#aZ+�|4��V�k{���G_�����Bٮ��lĖ��|��,y�)�YN$�bX9��Bg-e��mE'B�_���"̐e_^t�i��@�!�d+������;X���/�\Ȱ�nY��\�(�Y��`�Lf�}l����?��&��L���섓w,y2���5�e)��m`(%����w����Uo�%REK";Г������
/.dD>�)�#��P��gHܲ5��N�x�1t��#l\��,e3b�>s�f|̓�r�}7A��~���c�s��q����+_�U*�IP���u�{x�ʞ-�Q(Z�����1���U.��˶R(��e̪�as�y���[��lǿ��x����9��)�>Y�C�t�wB���s*J]x9�vt,c���8K9鲔�"���B��)̟�9�c<N��>��|�H����W�������2���S��gQٽ���SJ^�'�V��J��׻����!��m�����(��Ol�'6��9
���?��WBsA���9w�mڭ����r�ܵ�]�/�}��Z�.��T�䅐����B�֯�)z���児kw�K�>v��1������r&���a!��|Jr��}Ȟ]���U�J����>K!����~I���U�(K!�������n�_|c�0d�7�RP^/�Q(�P�����<��H� *�Ny�M���Zʁ|�Q����}�.u��%\0줷�V��y�U��h��W��-�1�Ԡ�I��vZ�O!�y/'��W3R\�Iݣ&u��y�s>�~��C��u:�
�:s�</@ٓ�uuUΓqT�� V���V��,���W��Q!������E��q���yYGe��(�������W��m ���Eh/�h��ȫ��/<�p����6��?����y��rH���ڝ��U�1��>K�9�d����l��8�8�B+�v�6�~C��&|�ܫ��mD���ߗ��?T���K�[ZU�O/�Nճ>��p���S� ���4/}�L�#��
��#�������{�m�=����d������K�vyh��u�/��О�BVz�B��]^�i}i+�K~����(���G�@}C�O�#|�0�;�<i)��LeO"��K�e��{���f��OYB�{Y#�#����T�|�^�f���u���e8�}ѽ�'�:з���\J�CMD�]
�x�Lf��0�)��C�q�s�����XJ�8@]��pG2{�0�`����Mӛ$����S�3�'�!�YV�z�[��|����C{���z��>Z3�%����Ly�V�����-��^��4�i��Wۙ�W�)��髖��>^G<}w���A�ry�z_(zѱ��}ZE��!�zVp��o�|�]f+� ]6�!_����t�ݯ��N���({��X�S��;��9q7���KXM沽I�vB��z����0靅p�cʕg�2��C���,X<��9�-g�y�C��d������S�J�{{�8�I�?�i�U��j����~��o�*~O��ݷ���`�/��n`�l���o��:KҾ��	`9:�3��F�$���n6~��vv�Gs���4��0��O�ǭ�.
�X+�\?��.=.1w��;ZF|w���s��5C*�D�ck+�o-�S�B*�Ƒ4E}B���~G�kc;��hfh5]s�Jb���kNگ�&_ē5% ��;n����3:
̷�^��kl~�w�F�t.]"�Զ��S5yf��P)M+A�B���Y4�ɢ���x�ʽ{�_j�)�&y|y�j
Y��m1M!�U���q��;��������G0M��A��]Z�K'�zV�>�c�)g��~oI
.^��z�j�ʯ>K4��@ngtǥ�3,e~���vڛ�?®��z�{/w�"�=��,��R�g�@��!![[���uS̢5W
y^>�8W��x���tT2�. [���K�������wz��h�^���������I��Α�"�\i�st�o�?�=�m3u95򎌞�zQf��
y�=7\éۊ����|y��R_��Y�4d$�v2�r/����y��f�˥lƉ�
6���E=bIuO�]�U�%ͥ���u�����b[ ���0_�ѻ(��TZ���3n�/�ζ6"��A��J�DZ �Fv0kLϡ�ӜP۶7�/�p�O?���=[GG����
B�纤�C��uIl�q}R-�����{t�z�P�O:����h���y�yx&?7�Ϯ�WN��R�&��XH�������h�~F+D��Z�����QTl����Z�|����gt1*pr�ꉪ�7�Dm������Zm�m�`��?J�8%x		����#V�jȆ	~���<J�M>Qʻ�R�~@�8��bߧث)� ��v��X�����	�O�ڭ��_���羝%4��{`C��?����Җ}]]S/)�6����dVTء��h��nɴ��9?��(Rf�(�{��4�ATo���}�J�������;�qݔt�>�}7��+�^Ȧ���K��UGQ�)jq�j	������0�����S��kz�%��o��s�k�S��K-�G
��@|g�T2�+�}����'��-۳�F����
�j�<���u1�`qL�M��x,}S��U}�2V�����*�}�L2?{����i
�p�;=��u�)�xhޟ׈2B�䓒�����]7������lhOt�Y�d7�&X�˹�ߣ��z�,~�9�a��K�7��r=���S��^.��dt�ƻ�E-�&(7��ȣ��|��}:͘�r+�7)��{�j&(v��'�+b���̼b�)�k�Ť?[�,]!���^�;������W3�u�FZ�/��F��11��/4F(|$��-�?���?ٿ�i1j��.%R�#�1�B���Ez���#��x��E	�x����!�F�Y^�s󢅰� ?����ȏD<���K��N�u������[)�)��_)������|a%�B`Ui� ��Z���M�x�T����G�ϟ�6�v  �������g��'�	�'�	�'��U�m��8�?�Bp���Rŀ- ��l����rf� ���D�S����po��;����>�
qC{��<�e���l�R�]���x\�9��w{�ec�����o������_�-��*9,�������C�$@��M�������ϋ2����R����ں�|���{N�
�=�����B���v��*Bh 侄��#�� �>��VG�~��"�&@�A���Ľ�-[�{�!��/=Ͳ��6B�*x���������oD#�#��z/�IoG�#���#��OPN3h����,��<T��d�������
�[��+�-�M {A�P�2�w���wu�kGF�TޠQ<]5��D	�F�X;&J%�$��Ӵ�6�㸿
������ h��%$���7�~~�P�O���N_�y5޸bp����(!���w�5J��o,�~q���C9��Q��D�4'J��%WF	�Wy�l��뮇{G
�jD	A��0@�|!OW���Z��x�fD	�3��U��Š�$J��Ȋr��ݗ��n��E<_���k�Ե��u]�0�6�O�͛?��(��n��u����W����'�	��ß��P[U��q���?J�����z��a`g89���|M���e�d��ɑ����?enfvj�u��S����^�?-;�=Ow��@<�s����`�O��H�KY�N�;uVb<����������-MY���K��e��g�-��w�-橙Y(eڥ,��)�K�O�Iq�qZ��R���Н�,m^����| �?�M�N����-,���d����ᐕ[���7Ӟ�s����uh`PD��x`��!$,B8<p\ap8.iQg׶8�k.���uv�8����Pvt��C�<1����+�\����S�����(�L�9�=XR�rrD)h��f����m1���~p��T?P�0��.v��?�b\�rpor%̟S1/?R�6�:�*��pq��1�R��Ɛ�������%�9��
���"�r$��.�Yp��]��_�*�g��=������ջa)y���7,�����r�w>�i��J��{i�k��W�!��}��)R�oE��p�Н��"�u�F��m4Ŭ�7R(6�a�E|;y:/e����S�c�o�'n�7�g��g{Pש��=�^g�E��v ��4W�h�g4'W��D��|�u�`���_�J�WqX�uCE�qj��y(J��[�[׶�g�����I�" Ap$��K{��Ub�d����҈����jճ��W�3�qg�.�XG29�఑#+9r�"������wv-S}S���F�M�a
�g����@�sǠ�#0@v(;�Ɏ3N����c該#d��~��$;F�.;F�!;�����c���#l���,�";.&;&�SΖ��C7Rv��d���a-;�cd�}��p�+;"�ˎ(��qʎ�EBIRg��6��*����n_��7��x��ϿZ����;���P�C����;���P�C����;���P�C����;���P�C����;���P�C����;���P�C����;���P�C����;���P�C�����u�숹HvL�ʎ8����.�13Yv$PCuTz�p5T��&ǒ�P�
BUC��,7T;��o���HvXe� ��DiI�E�B�����*ğ�T���&�F� eR[E���Ȑ���{�G��\F�E��@��Iޭ}��R��Q�{霐�;l��B��*v��K����d�u'��Ŕ��*��  ��8�O{�ϡC2�ZI��:��fQh�N��(�?"�AA#(�"I�1�]qCJ�
�J�
��1�Ce��e6dU��K<~��*�(�n��[x|�o�l����y�x�\�N�I,^b�7�x�T�A����R��M!o]B�=����ث�)t/�FP��Q�>NA�)(�'\E	7R��:���P���G�#xh���z�<����F
�I��Rh�Hj�!�L��(�=��B�S�Z�У��{xI��=G�f���<c}��n}�(ߨ���׆��R3Y��
�p	0H[��q�sPJ���(M4������Ҵ�H�{��=�]Ǜ��8T��K���&�!0b���(�Ow` �k��ש����!�7��vR��Bk(�#�QD�_(�
}��N2 �L
�L����Z
�e��@����D#B���,
]�C7S�[:�B����;�*�ю:j�غ�ZJ�u1j�L�s������Cx�$&Dz?#2P�놮.��r��[J
�\KiҨ��q�0��P������6EIg���Y�3݋LQ{(��j�â�STE=@QϟM��)��.���{�#<�b��oI�#<mIʧ�B���#<�뺺.����	��~��c7�������'1D��p
�D�Q�ϡ�	摗�g���D�M�������zb�Z�.1�����w_7�Xm����
��jY !���=>\a�z##3̊x	M(�P��¤�h��JU�(�>J8�^��R�o}�Q�D������;���p�R�u+X��	].���F3g��"?Q�i��6�̵�p�P�¸Vi��+�M@e�PY�c�c�v{�⫩$�)r5�<��KUE�Y�f����FS�+�Q���չ�lj�.�[c�%bz4�͔5���;Li�iFb��)/����!�Y�
5u5Ow9�_�ui5u9�Y����4e���7��6�iu'E=�4�ʍJ�Dޥ4��F�#�0K]�_����רk��"��+ְ��UcI�S�SBT:�u
���J:�%8H��O�?�"Mң/�����<)�񱀅��j�	Z��l즾�����O�����}��ݕ���rvRh;�Jw�D��7<��Drٹ�sP+T�HHN�����K�u����{Gݿ��"���X��qc=�6���ʍա�T�PĨ!w�p���<vC��ݎ�ٙ�����R.;�\>����ܿ�o�\��&�ɷ�U�r��?ӧ�B=�s=���d�﷜BU_s򽅘ڒ\��x~[��� �c2�����~g�o��:�Pn���y����u����u�O���#�Qoe���'z'/��2����ӱP�"MƗ�(���;��V|y���T�\_���C��Ҕ[���~�n�(`4���M���899������T���t?�����Lv#�rצr/'?iU��i��C�(VF��6#�Քw�7~(��{��sC�r�u�F'�������WyYj��X��S���_ x�=�@�wD��1C~G��P��6�M��{X�}�=9)�������$q�'	�6�lU��m��z�� T����M�����_��6���R멌R��R/=J+-����[K�|�p�L�o�rnkwN�=�{���}���`_��{�8�D�_��e��Żk�����K����Nʹk��s���*%u���|������M'߳мM�2�����>8�{Ll�o��p��w���C����ɜ�>�$��.�q���~�����c���d��V�1�ZO,�'�a��͓�-I=�z��1ԇ�4����6��u�ǿ��sR���Z�^�mݽ?(֒چ�I˙=�D�ez��SU��0�������_�k�j��d�S��$��7ˊo�)-8v���~�:?BqA���* Հ:@����7!��}F����>�E�g�|��3��ś��/c�}�׳��>�p�O�;����'~~?�����_�O|q?�k����O��~�������~����o�'���x~���~�C�����O��~�����O|u?���Տ���#����'~k?���ć��~���8q|q?�m���x���~�s�8>���W�_x���SO���/�!�k"�P]�`6DA�! �^W���oվ��G�~�Z�ǟ|���߄�/��n�����J�gd�3�����?��Rܡ���N/�&�%2*:&v*���f�%�T�e5�"��x���g"��x��s�YxF�Y�g���
��xf�Y��Zx���Y�g j����ٌ�(<[	�xN�3`5���g��x^��$<��ӌ'71x�.<G�A~�n<mx�%�x<�)�
��4�%?��ǀ���x��?հ~<��&�ɏg8�a�鉡k=a
$�3������%�˕�������}mn�?�P��B�^
y�I���m����B�^
��.��P��!���Ө"^^xo�)E�^mE�����v+��H��"^�E��Ro���I/��k��6�l���F;sذ�=Æ�9rذS��>l����>r�ȓ(�l��5b����g�1rȐG1d�YC����򳯲G*���ס��+���ʠv��5�����#�sU{������nlV+iH1��Q+uخmB�6��̺�O�%�$�\��_/��/Hw�]��JM�r@�	�h�:�AvB �a�I `� ���d@* �VJ� [ e�r�.@�Ph 4Z � E�*�(+�QR�g��\,?ë0� �{	�z��@Bu��v?��ƃ����h���G�k�j��Z�O�
r���&E�)�KQP�"R�i�3�w>O��g��!�SI�)?���ژHaRl����(s�S��;a,���)c<��_g� ���%�$C�M�Q�`�8�g�~~�'�|�" 
8��S�&�{�NPx� ���N���8p�i� 
G^
?�ҟ�����	������������8�ӼE�x@9� ~�B�y 7`�Ph?F
�@ P�
� !Ơ�ƻ3`N�E@�0�	�w�%&Le��P�d0���B� ��-L���ÿ1Z�� M��;���m�B��p�~y9�(�A�x͒��i��!ϐ����x��G�������3b�T�c m��a���4�er���T��Q./&Q��Cr�����l)�r���-�a2"�S^Z�eJ ����Kc�"�B��O���V6�r.C�H#˻R�5�T��T"��V��(BXܣ�Yx�n��ʸ��D��r.��x��n�g�xf!���j��I.�r3H�k��qɀf�[�e�&��Q�۸�Kų��,�1�
i��߀�"zOć�O2q�p� �M��4��A�{ek<� �ew"o9цte�,�R�e���(�2������H��-�B�g"��6.�i?�D*zw<�O� #�Fo�ک��l%�p�-n���n�-��}w�?���#��+��� !\&� t ̬
�@X� !N�F���<�k�Z�
Ӽ|�P�݆����f�7�}p��U�0�� !a���YKF�UX;V�
+< lAX�*��v��}|��Z��3�~���?�+ ��<7 <�  �hHT�To�� �� � � 6 ��� Z���E=b s �B��f@�y@��
�p�`���H6����*��|OO����/�0;��� Y�r�f<� ��z���)�
� ���, ��� [� j ����3^
.X��<�*�f�3�j@=���r�0�L\H,��T ^|ht B�k��L@:��p�)@�>���xJ���j�-` �H��[�  _: A�Ѱ��t�9�e�R���]�Z�{�/�4��١�p�00� �[��f@9�Jk��������s��R
�zݔ�,��>{y�Լ������E�?+-2++g!�O����RR���fz��J[tYAZ��9)Yi��s�KsӲ/I[������OC�P���������qS:�^TN!�����̴B�\aIZ^vZ�7WV�;o����HC|悼����,z3��觘��ܑ�livVZ�����sxR�>uz~6��rb��%�9ٴaN`��������4%{a�H��)���g�d�x���Ҳ݉yi)���P\.�!!����4z�ĜY�̨�n���N�Q��=�S�˙GUrKL�G�d���HS�SLZz
p'M�O�^T�JW�؝���H����0255m#����Z�������6�'��\�LY�	MBc�U��
RRǧ����\k9KQ�x�l���I~;�ef�N���wS��06�;�0�Ή�ܔ�4/�	s�2݌Z���3ث��.L�u���R����'�df{Cb�S/M�3��YI�סh��)�����4FO��j���xv��i^���/&-+͝*3QK���H��R��,�y���	�Lp���d�3�J�*a5'׽�%f��Y羋��}�w��woW���(ޜ�����ۈ�rs��
���*!�Ku��ޛ�d�����F�Yi�.X����c{뛾r"1-oif6���`�B���>+-?� o!k�ٙ��S�xa�٩DB�|�,�K�<�������4gYZLf0��-�%���H�zI�]��Ֆ��������$}qމ8�+9��L����:��]�v�)���E�PHb�R�,�&y�de%��3�Xk����������d�/az47ea���t�|*)��������%�u@H�-2��l	�S�XL��Be!���.1Ir�HL���'!SsQٱ��2�r���p�uYU�f,�F%g���)ݗL�M)�/Iǥ�\7����+�c�B��+z�}���ŒI�&Ƈ�"[-����5����<���,p�*�7눅Q=��u��|)��U��A��Qu3�s�~u^^��<ċ�W��������S�P�n��ȕĜ%�<���YR�����Ͳ�[bd��|7K���!����a����E��,Op�]�>-;5�PJfEL�T�[h|�P��$��eѬk�:V	��]��&d?�����iy�2y�a�)�Q�陌٨�T��?zFJ6�_���$^iǉ�&� �L����F�$�e��6W�?Q? f�K�Ǜ��e�����c�`@�4<�c�O������`A蠥+�p�F�I�k�hvi�4-�M�V�&jS��ڵ�-��}�Z���f�O�`]�N�����RuY�U�-��t�F��u�����&�t}�~��X���^����>H-���D�h#�1N��Dq��,�3�\�P,׊���Vq��C���Z�^l�EIl;D�h6�0����a�3$�n2l4l3�26|l��lg�-���+���ƍ�Ǎ/_5~n��x�i��d�n�o�7�jz��逩�t�t�lg��e�n�g�4�W��4o3�1�l�35�Yζ���̳,��h)�l�l�<cy�Roi��tX���V�j�N�η^g�׺�Zk���fj��v�m���v�m��e[��c[�-�oO�g���B�*�Z{�}�}�}��̾�^n�a�e��W٫�5�Z�������j�8�;;np�w�9^t�s������8��wNs�8��9˜;�U�Fg��Wg�k���Jp-q��p=�z�U�jq�D��b��5�ݣ5�4�5+4wj��Th^�|�i���^�5k���m=Z]�����Eg�]�K��6�6�v�^�}��Nw�>T/�����3����Կ��D���������3���X�q�h��Tq�8G�ZL��e�
q��A�G|H|\|F�#�,��?���07�5\`�b0������9������2�c.7�dn67[ε\`�Z"-�,�,�Y��}�fi�tY[�Yìk��N�f�6k��y�~��,G���q��i�ǻ��]�@����Lw�p��|����{��5׵е�u�k������i�k�w\����M:S��<�٩���'�ڥڧ�����O��3���ĳ�1���ŏ�;�6�5��0e��7?f�e~��	��XL�X�,˽�,�X�e���}����h�e���g��_9~pp��<׹ݹ�y�k�k��RW�+�u�k�K`;Fhm�ƭ�-�>�yL�f��e��@�T�L��m�v��D��v����� ���l�r�=����|9z�*�Z}�~�~�~�~�~�~z��/�N1�1^cZk��t�iz̳�N� �+�Oڞ�U�\���:�;jM��;~�Ø	|�n��>p�O���}�/u��N�,6�@�\`r��G��c�3���72[�s��������m��-�%Ӓk�=���ʺ޺Ǻ�����:i{�6Ğd�l����l�X��9Ϲ����]g��;���Jq��z�U�ڎ���tpvq}K�6_`�s�A�X�	���ho�ޥ}P���Y�n��'��_����u]�n:��5�L�&�Ӻ_t�S���V�c��������k�~f���|�r��������,���@_��F�M���Lk̷�+--C�`W��γN�v�2fo2�6�7�i|�����Xe�o<d|�8�Tj��4��Yk��\f��R�� ���������Ŷm�N���Q�����t{��������3��u�-�[]_�hkv���qi.׼M0�0E��.�XL4<9{�q��l�3^j|��<Z�g��	&��i�5��\c}���u�퐭Öb���tLs�q\�Hwd;9�t|���9�u�K�JD�������D�Q�/6�t�2�Fͷ�v�:h��&p��B�C���H���G��A�)��t��M��t{tt�uu�wt�>׵�:�A��h}�~$�])��O�v�һ�E��Rp�}����J_���7��-�V}��S �!����b����R�,�-���Rq��E,��]b�X#։b��"���b�`2�F����n�1�ɆTC��m(2�2�6����_U�
u�C����jh7t�A��hc�q�Q4�㍋�7@�=i�a|��`�73M����V�v��LߡǄ������`����?1i�����7� ��ᖱL�-N�T�L��ՖtK6d�
���=��,�C���<dy���˗�o,?Z~���^`�b5Z�֩֙�9֫���l�2�
���c֯��mCm�l�m�t6�-�6�6�v�m�m�-�v���m�;m���=e{��5���綯m�ێ���a��v�}*xt�=՞�X�ȵc4�.h�{����do�Ll�w��!�ю0�$��;b�DG�#Ց�pC�W9�8�t�;B���˝9Ε�;��Bn��<��:�5���e�>�C�Z�V�Ӱ�^��k��	�&��^���Nۨm�6lѶB�wh;��.@���Bt#t�a���uF�ź+u���2ݫ���%?����Y�	q�~�~�~�^���#���W�� i7�wU���mЛg��h�T�ZH���JXC��
2���3�0�p�a��!�n�K�7��0���g<��l�|c�1�x�q��n��6�S���KL��rM�Le��rpL���Tc����75�j25C�J�VS��W�0��4�CY�\�Z�f�v�h�
pU���\˨��`n47A��;̃�_a��fK�%ޒ`I���l�oI�dX� �ݖBKd�z��~�+�&h�6K�%�h�[C�#`E�Bn�['Y5����Xk���M�M�2�.k���Z˪�Zom�6Z�����dm��h����x[�-Ֆa˲��ܶBX^ŶU���R�F�&�fXa/�^��lk�t�	� {�=�l����������v�F+�}���������]pC���5�B3�0�^L 7�?�:nq���-G�8ju�zG��ڱ�����6pil���N��Lt&�Iuf8���N7�"g�s�s��Թѹչù�Y�l�����pv:W�+��
v��F�*g�����f�R]n�*�/]�\�][`'�,w��pU��!?u���A��r� P3B�	ӄk&�N5f�]����a���I�x��)��ު�˱JS����b�P�i�4j�4�GH�V�����h#�	�y�d�|�*2�Y�\���"m�v��ڭ��a�ԡ���w�u��f�2t����C7�ݢۊ��]W�ۡ�ۥJW���5������'�o������H��=0� C_�l�2h ���� �����@4At� M=@�?�:�Z`-��Fh���[1z�'��Eb�� �[�0r	��e4F/a�LBaI]i�z`�[��C�&��.��6��>�7H����#��и�q�	�D�<c2�z�1Ø���۸�}���Xkl46[�����fl7v;��L�� S�)�n��"L�`f�
MŦU��JM!6������a��~ȃo`��G�����b7G�c�q�xs�9�!�<ߜ
�o$�H�z�D�̭���!:͂%�h	���\�ِ�#VY�ZJ--�0�ڂ�U��}�G��BO�`�FXc�q�xH�R�F��v[_��������#!����=n����2���
[���Vc���A4�mM�-�����Q����E����@v��@Ìq�sB�;V9�b̰v�.G�܏z��N��p:�9/tFB�\��չ�C��ί1�8��r�jO��b��a�n�!���m����n�:�/J3Us�f��T�]�}�����6XG�N�� m l�`m�v�vzY��]Er�ڨݤ��i��L�c��]�
m����Z����kO�Ӎ�];Yg�9t���$�U�4�R]��F�j�z�ݺae=�q�Kl����W�����c.��B}>�ѽ���+����4��,�d1��z��i6�O�=��8����1�|C�a9l�G�alt��,�~1�
��htg�׃��<~��68�'� �h�E�ǚ����ͷ�5U���2}=v�t��L��d����k��ͷ��1?	-���3�?0�
f���p�
� Y@U��,Z>vYN����o�[��I��ۺ�z+,�m�=�wtZlA�`[�m�m4�B�I6�M����"l1�8h�[�mt�|�RXBB��n{����o�_l��q�|b�۳a�l�?����O1��	����Ʊ\x��.�_���׻Q�/��a�$���b�V�t^�������q��1�u��8W��y�d�|h�W�+���U�*�Y�M��CT�j\M��\t,�	�����h
��\��f�g��oi��v�ge~�Նi�������o�6�"�i�T�2q��ۗ����?����N�EB\��W!,�;!�+ �ku���^�tͺ��q@��]ׁр��bD�1�6*��_�_���H��Ð�C�9��:XÿY��W��ls��9�O�	B2�5����C1��A����B�d��^3�3��ŝ|���x�������^3МT!Ƃ�̣���[^o���:Ǹh�8�zB��S�)ڡڞ�����������q��>��rf�1N7��0Z\j����i�EoqZ߰~j�����,{��3{��2�n�[�.�9�n�~B)�4����r5�����20��Y4��z����k�7��h<n�#�A���3LCM�M�LcM�M���'�o=c>�Q�T˕�K��WX��v��R�j��:[�� ۾�~��~�s��%�X�3���SYHG[��� �L�~��+0����vެ;:|��j��_�;�/�����֗��T�l6Xo�� �g_4�����r��l�6��ς�:��9�W�۬YwZ[����xd�c�C�p9�omr<�x�1��rN�h���zɗ��]V�t׳��]?��-�������#DiӴOjo���~�~�>V?G,�0�"N�7�%�΃��ڰ��a$FswCMW@�~c�`>���4[B�E�tO�K�]m��m���|�umB��e����{�c�#v��λ������8�ў��|׭�]��� ?vx�f�Z���4_h������;O���O���=��#!���ߠ�R�N��������<�ֿ���{�����*�F\�/�&�-����V�%Ɖ��W�a]/�#�s0��l�i���eX �d�q��%��:�ǰL�n<�y��a��U������Oأ��;���.��.!�O(���0;U{��ȋR��ס���&#tSt1�V��[�>�0��F���4��&�/�;�7�ӿ��\�=��M�K��5�6iLf��Lp�荽��'�<�|��e�Zr,�-�C�[��<�1���x�o�h�%h�y:.=�O.и4+4ςo��	�NК���sC}��}W���?��h�Nם�;W7A���tѺD�պź�Х��o�u��+�ؓw�o�ca!.7�e�=jr���_1�{��.x�W�X���h��Lw@��3�=Wd~����C6f�h)�}�,��[Z,���1�zc���Z�0NZ�q�nXF_��ni_bϳ߅���� �O�]t�W;�[;0ry��c��*g:�!��;w:���9�s~���������z� ��	q�c^�<�������˘ݝ�f`
�#�/nf�0�ѯi�D�Û�\L���@1��Ǆ2K\�l5���Y�f����Rf�oes3��@�3�b[Q��ZS��@f��f�
4KC+4OCk4S�a�es5Ő�4[��Y�d�W��ZH��i���Y�H ��	��B37�F�Q4�a���NV;��d����`�l4nb��vc9��a��1��.㩦�LcL1iM6�7��OSM��ԕ��ͦm����0z?��9l�� �������Z��<�|�9ݜm^n���L'��<o�,?@�$ZS��a<��쓛m�l�ٴ�4��C�7!c>�s��1��aq�ޥ�^NX�(p� [��q���#�'0�}����H�F��G�8~vt9�C`�r����8m���:/s�Ÿv�s)z��Ε����������s�~z��d�1�w��~.�n��e.�(4ASK�#Me�f[/vp�v�|�RXǥ����*.�E\k�Nۀ�g��O7��vL�-���#�2������>�}��ן�?_��Gc��_~rr?���l���<��8q��i�Q|����~�9'x�JpV�a#�fC8'�qN�P�=����A� E�-[�\e�6�`�Wg�76`��������M�dp��rMn�􊺍�v�F~�$�:0�6�`�7�j�Ho��Xo��F��l���יe�l�l��y̎�kdWf����SK�%�r��]�5׺�z'�v��^�{��-�`oG٦��Ȳ���l��}�����`����-�>�n��E��nǈ/��W�����в�в�����ױYF��jo��w�G�#��v�8F8D�QI�,���ɱٱ2��y9$%��`���=a ��p���q�9�	���u�����p~��
\����u��׫~�����F?�nf����j.Ӭ��Ӽ	�~:t��Hm��m Fp����kuź{�_���7���A�Z/ �.���+F������w�9Q�mO(�AQA�
�,3���l�Uʺ�!�dw#�$&Yª(6DEĂ�X��.�ذ!�])VPT�!�W��}�̤mX\�����]��s攧��s�L.��d
�e�f�	�����.���!����Xuѩ:��r��1��	�j�9�N��FķM�fh���;/�>�W�(���س�:�rc���vw�w$��1Я��ἅ��]��#1n�ٙL?��@��@�3����9��������"��Y�M�K�Ox�{��ͺ(�Ѐ������pŢȰ�.�T�R)������*K3�%��_�ߩ�]�ݭ[�XG�w��y���d[i�bS����q�t�+X�Hl
,��Q��9��8��9���&���Z�R�͐ Ź��m��\�7>�Z�z����E�+���7]Ҭ�v�7��]?�4|&�6�]ý�m��j����=ߏ���ga�>q00�D����-�~�u��G;� ���C�%
[s�X ��D�x�͝�[뀏��xh�S��+ ��u~�0��.rw�`��|8<� �D�#�)_%�QnQ:��Յ�]�⤦��N�N�ΰz��1�l������i~�j�u���]��4k��a��}�}���-����G��d�d��Z`�ӜAx�Y�_�v����J�5�!79oE<{�s�s	���W�L{���=Q$Y;��M��3x/�b��1D�gAO.�����_�߱����.�M���]���b��J����g O>%�''sd4�Sf��U.P�+ �$ov��L���~����o���鰙w�����wZ�>h}Ժº��,��5�W�o �n�~`�����K��֝���~��v����m[
k���+$�qX�#�c,��/:���4:o��vD<��u��Aף��U�g]/�ָ^u��zǵ��'��`y�v�����w��47ebޣ1~o��}�_Ͽ	������+�����'���DA:8�~i��`��|=|MG�X�����W�ӕ&��z����˔+����FH��=��#�r�D��*�:��F�݈~uY\����j.t]麆����3�$s�j�o���V�g��τ��/Bd�
���|6�������۾�u�f���jԾ����t��#��.�C�e�%���+��;�������/6^by���t�<Dvȗɷ�+�urO� +ouZK����z�u��e��!v�� �ˠG��7۷���s�rt��R�	�Ug�W��x����n@f�9/��<�|ɹ�y(�!xN6��c���gEx�0{���#]��D|ӝ;���y���ܹ@Q� E=��8��5���<c�	�o���ʻ-O�j)fB{��~����9��<0�`�K`[���!������au4 i>�8�9�u����i3t{<{9[�=�-���YR�]�8�-�D��(�.6�+ſD��Q�"u��Bq_G1�툣�Q/U�To��=��U?S�r��3@ۖv��2�OwÞ��Z����˗���ʹ͵-y������n����TL2	\�x��;�^��e��Ⱦ�������(�+���M3^P-�;b�َ��%��J^ʓ�&�B3p� �2	�������78�9oRy�չ��dYs*t�.����*�C<˵�uC���\k]���r���������1�cV�#{��CX%m�i;���z�6��}-���ٛ�������2'n��C���Ԭ���;�F�[�O�����B��R	����Q���M�w���_��U����Rno	Z�F����Z�ڗF�i���hU��v���9X�a��Fa������!u��t��D�7#�|Oܬ��E��?i|�2N�
D$��Kc��hDI"�ՈޢkB;�]�n��;�=徲Yf�
y"l�_�#.���[�%;(+@�')�4_~�r��Ry���&�Y���oSOR��>u�z	4�6���u����#�7ЪZGZO��[#�3��Zo��<k}(~�U'h��V-���l�lۮ��g{���o�N�C�C�#�'�OET����~�}%d_C�3y?�����rS��q\�̱���ǋ�N���,�����΁5�����D�_9����΀�.r-�嶥�~����ܵһ�����o��ufe��,ak ��؋٥�m�#�j�mv��3��P��I/�+�����`g�"��5�u�(��b~	p�c�*�y~���f9�r<�̘���j���dZ�'h��%�Z��v�I�",pBlh@�#\���DO��鎼߅�)+�Z�d͖����4c�9��4kr͛,�o׉�?�HGI��"I���ڱ��ҩR��f����m~Pzu;�h����W.�,ϔ���	?���x�G>X�X����0p� �� �/+�">ݡ���p�?�Lw����U�j�z������C�]o=�^���l����j�޶n�jg�j;2{�m�-l�m��X�6���t=��O�]}]�a�-��n��cҮ���8d��#͈Bw��������D�ݜ�8�t�<�iqڜ���5�)N�s�3�<�y��R�UΥ�����9�r���Hw�vr���:�es��NrMu�]��������V�h�\ Y�)w �e���A�_��o��!�q�����@������n���Vr/s��-�w��\/���"� �ֵ����s4��'���b������ӖW-X����u-d��S.�^�1�_����$����-�����׊o�ŏaM��*9�J�!}����yҝҽ��W�7�w�Վ#��c y^9 �-?/�!*+�N���)��E:�8���l��=��j_��jN�I���L�w��UY�ޫ>���~����A�Zl�b�XgZ��3����^EW)�>f}����}�	�X{�
lV 70I�v��r�Ͷ�l�m�!�;`w{ ����5v��s����
Y|��*��K��.���ň�Ou�aa9nq�r���<pt���r$q�s8��B,����/�!:а�W�k�kt��F�_�j��U��`u?�������OSՎY ��Nw+��Nc}���bv{7��]þ\�-�;ە��I��u��7ѽ�p�/Ww���]�� �/F�M��~��@�qt�i:]A���e�e��?�NB��c���A4x#����S�+�z�o��n��:.�|>%�۸K�[�%��I��ɍh�"i	P���*H�G���O�rxn���L%Wɓ䩈6�e�Ȯ����M�y����K1+��S�z�ġKi�V�V6@Jw)�ui�R�PoW����ԏ�/�����Zk��$�)��q�'w@�X�X��2������S�Z�sv��5>��b����������.L�=�~��s�`����!���z�^���]�Ž�s�U�j� ����s�-s>
����#�n/� ��:�� )]d���$��.fF;����l?}��='z��^E��}��&���P�I<�x��k殄�^~����1$�(}��v�&��h�yOHӈ��Bhs�� ��;�W���{Rǈ��ǹ���B7�_e .��`��WHwH�A��O���	~.�j|B~]~O6��c��J��H�������_Jط	�)�L���X��~GYa�&Z����>�z �j?�q6��}��l�!�}H�O��1ɮ�����;F8�n�7/:^q�w|����sb���(N{ޜk2���y��I�k�-�t7بש�9�+\���?��+�ak�������թ�h ��Y����fo`og�GL�4���h\B��ψG�^�����gH���z*D$��{�{�������;���O�C���2�A�����'|��2��<˵��,��k�	�%!/X���>Wq�p�p/8�A�X�F0�G�ӄϧ�Aq�x]�zD|A|�f����t(��p�%����HM�i�t}n�]�s�o� y�,�N��������
�y��������U!��H)#%��x+b�'�5��U�Q�EU��F���aCB��@"H�D�E}����:Z����α�b]o�mh��uH����<�zzپ��:�#�g��Yw_�G�g9.q,�]X����� �qΑ4ޝY�O��,s��|����Z�[�͈tw ��M�ݞ�t͈rY�_����u�ԣ�P�\߸�&���/�c����c=�����3��׈P��K��>.
T���.G�Cyި����t	������
 Y�Z��_dY	x�Z��,�����}\�N�SX)�'|!�)t���U���s�+ć�g��F�Y�/�,@?��(}7aT��{��O.��a�3>��̑/zڿ��"��q�M9A�V����y�b��[+�',�2up�j_k<C:�~� Y�!+9��}T{��*}��%���l��ް}a���Ȼ�������ܒB��-v�����GG/��RX�F����CN�r�	��"�C�nl�1A��[ k\o��h{jix�af�a�gUv$;��o�v�1ą[�������	�4n&w.wwl��4���c����p�A�$79����
�����������d醨o���u��N˛��-��4o������jd����0��;��YV�4Æ\.�(>D�c���ؑ>� B��ݨ$AV��e������y�/�=���9�e7ݣ:H�:�M�^�宻r<�(�J9U9^�z�e��I�(�QV��u,��r�����5�t'�7�O���ჼ�j�Y2|Z����C�֮��!����I��.���������mn/��Bw�^l��~�}��M����T�z9Q�\�8�q��c�| �����Y�Cdvd�V�K��`}>r~��lW�}ރh���ˉ���r����_F8��J�v
D�v{3�(�<�Xd'ݙw(7�+��qӹ8w	���k��߸N�a�NV���V>������Q_�4�J\���*��"�Z%=�v�m�R�Q�Iu�(�ʡ�9�8�w�<�Y �5�� bP�5�t)F���<܎�5�g�:�\v{�*�)F��<�kDL����{�{�;��ͻ�����"~9�,t�ď-���U��Y~�L���/���/�K!�7H�I]���?���p��%�f�h�y�<�uYDQ)A�Og�;����mp�@�������W os����#�2ʵ�u��$8�3]��� B�����#.~��h�~��<��*K�q�M��ϊ���$;��#d�Ie�26��u�5���c[h�b����Y�z����X�]���H�a�jG�����d�e�\����D��_���!��/$^&�-�'v�����O�t�(���ԋԇ�����V��r�;�m�>���b����²~i�X;);O��6�y�'.�S	3�64�
��#v _�_����jD���K�C�?��P�@��:�z��lg?�~�}��'{�u�q������93;�5R2�u�k���Վ�Z�@*���Q����򇥝P*� �(����� �f���a�����W�G<���Ѷ����*��	��ɬ�?=�QF/Ǳ���q"�E�x1����M��;�9q����)�<˹�y�������'6�p>T�p�k@�A�q�v@�I$L�0M~=��^zυ9r}
���A�FZ�-K,+,OY�X>�t�/\F��� !�xs�x�x������#�Fy��2��!j��S�ZGX�YC�J{f����c��"G{�f�Y�|�yY�ٞ��[���M���+�>Gdq�p�p��P,^+.�'�(O����~�u:}v�Qz(�*1u��Q�;;�:�zl�*�֟m��+�Oٿ�Ga7:�p�t^�|�����^d����g6^�'rop#�?i��_gy������@�3�\"~"�$v�����^�rPn�����˻�c�T�P�(���/���̶.�γݥG!�i��l/�^������d��C��6�v�7��i���?�������#F����+�.���UN��'�&�NqMs�]>����:��&۞>{7���`�zx{	>~<l����������������8(��lpx�F2\׈׋7���w"�{P|T\!���_���x�|�<L��8V�(�W�(���ј�$x'��a���Z�>8r����z�dX���<��`qO��k!y˄�@~�L��>��B�9٬��Hj�����z:�)���&x�	�sl�v�7�ɰS+l��.����aq���q��z�M�[w�~<�xԱ±�1Թ�������S՞�Q���6v�7�.��7�+���Q��-�Y3�U��N�ޖٖ!=�"�9Q'��L���_�}�A
�T"zyZbSK�Sէ�/`_Y���;m���"��Υ�����^���^ ��X����k;^>r�ȩg�'�c$7� �{��f��R�t�"*�����R���z��p�h��{ k��<�=T9>�	�ǲ=����>�藲��[Xt9�[��Jw���m�L<9ۃ����[^	�s'�0��j�U�-�[�#w�����X&[�����gNY+h��T��P���+/� ;�>~��D����u���-�pz��~{H��h�/�%-�n��~@Z.=�}]� },}o����Dw���_���y,�֧	�Ʌ�e���;�������i�������������V&+A��*��+�m�OJ{��z�:RP���֪�չ�Bħ�!�$�������Z`=Ϊ N�am��r���^�9.����x��bD��Yϱ>`[+��?l]�G؏�;�������B�R�mt7<�N����x��X���;B�9��t�`�M�M���p��4�9�9�t�ĸ��c��u�s��/gG�!�ca�Abb�I.����Z����ҵS���)����B�J�K�4�q	{=�f� ��=�ۍ�P	�r&�㓘�}n;�p�1</u?Q�u�c�������],�Y�Z*-->���-7Z��GD�����n�?���tWo�P/\Jws�7@�ݹG�5�dq.��4�#�TH�`���z%�]m�
o}+|�	�/"��&gW�?`Q{�9N���ؾ�GXfAb�9��!�k`�K)+�~�1�b�7�κ����D`�gm?�<���q� ���P������u�����_ 3���<�A�(�C�_ȏ�5���eqXΰ\����G�睄^����_L.�{��A8T,���t����O��RX����tb'���U�:�}�ت#���H����&�Qe%b��J7��á�Vg����ꥈ��o�X���X���P�1V3���tN�>���ί�?w5��p]����AkO�X����!7s�rr��S��������y�_ 2�&�#�p<�K���i��-�Dkȯ�"N�G�}�S�OY�w�Z�NW�C����:�*Ym�S�Gg"��׃�M��1 �W�OE�5�v��R���lw@����C��>��϶��"{'몀]��u��Y��,��A�=����ĭ�z!z�����v6|��<ļK��b�n�]zM�Z�^�H{�4L�!F1mD�#~�1��nPuF�[���ZE�I֓�'ڧAƀo�Yk�ry�����1ٱ�� �ߋ�w�f`�S]�\��^t�u}�Ȍ�s��{8�����ֳs�+���.gW�����v������Us3��ܣ�ța}�}2V&�4x-��r���Gb�����K�%�f;��@�����e�Ҥ���C��yS�P�
i:F���b�^mB����R]����𭯵��8����V�t����#>���	�/�����2ь�@0���X>wuB�p��LxZx^�Vh/c���s��2ˁc^w�߉G�/8��� ]���>�v�('+�x���Q���:�eqMf�����M���٭�$b:���Ybə��7����B~��6˳�a���N�)��1���W��E�/ ƺ�A��Oq�4X:	�a�4��Z�c1�g�o��z;��j�Z�W��S��c�氌�U��G�gT�8��Ϭ'�����\;.r=��-��=C�o��ޭ�O6q�2۟��)WlF2/[q�ș}i��i�b�|O���a�k�泙���y�lg�@�'ۛ������~������s����v{5{{�L��ax�|��g�xo��������N&�]��n���v�};@掭�|�]������2��f�@D�6���0}��,oWʶ/'�	��߁���=� joZ�ۼo��ׄ��SS��v�'�~��,߻�go�]����������������{Wy�����ߩ�W�'���}�DI��g[?ɵF�|��y���[�Sf�Jg�����d��ao���{����Œ�l������������j�%u��P�{�f�#u+b���1?{��XK����'�r?��+��M3�Oun�3���H�o���������1����y���?��^�g����������}Ko���O�_/����������������g{r'���|������F/�O~v>f"���b���Y��ߜ��e'�x���y�.Wҷ�<îa�`��߳��&���p�
;7�;���[���=�=ʭ���{v�mn�	l�7���s�n|/�y�/���y?�?v�*�FX������/`�M���C`���-�\X,���HN��t�t��F�.}'�#u��E�$��'ʵ�ir\�L�M�R>@�T(uЗ��J�ue��r�:H�NS/U�T_�l��v��I��ZH����OZ����~f����f����d�٢��l�ҧ/�u�D��>��o�;���i��o{/�0G)P�Y�K�q|�8�9 ��9�JY�Ϲ����с�4��_��<�����j6Ò��B����A���b��2�`)`%f�Ḃu��A۽�����m+�L��t�������+��Q��I�t�?Y��&oľZ�4z-}/�G�"�m�l��$&1ckЛ���93SՁ�W��y�}��0[;h�i��pO����߿�;��Gj�:��0���*��#��f�2��gs��wav�0�M���p4��;�
��X��86���sq���p�� ������kM��vֆ2w+���q7�G�س3W�q�cq�c��p<�0�p��.s�&���r\"�u��V�L�h׷渾+�u��3���qݜ�:����׫r\���z8���;h��v}Q���r\8G��s\+��.�RS��p�����Í�~;&�O�n�ܑ�?�|ԩ�����}zG��(�7�#35�����Ȓ���udf������)�tdN�Ji{|����$o`�B��M9tc�;S�{���%;dO8�a�L��ٽ�B%�G�N��å�_��^ʌc�2L%3��ČƱ�)Ǖ�ۍ�fʘ*\!׫	����Y�K���:��>G��_�Hk%�HY�)�aTn���e�L�	�_��g>��Ŀ�8b�̑Y���,�����Ʒ:\��x,����E�x_�ׇo!�	�=t<���q-��ф3/s-)U}�ofJ?�Ȅiߍ�鼼�@p%�oڻu�)��Q?��q}�Zi��/�_�(�f��O�)%8Fi)�i�~Gz��8'�3G�7�6�X��F!J�d/>f��Z/�9��%q|���#�Dt��g�(m߃:u�hs�ӹC�v��1����c�<�i33�(���E�N�z:������W7�mh3�����X �j�8�L�)Y7H)@��k�iQ;�F+M�)?�j~\'rEx�IU���c��k�-�زv�����-ѢvR�H�0�U�֙aC4�"�tӾ=T��)��t^���ڄtZA^f(�?��Fl���R"�{w�����Z�T��용d7$$����祽Է��*'Cu-l�ЍZjk���g^*3Q]r��f���'uS�)9ҟ���g�qO����bA�	�Cj�`�o��΢���M�u���Y$�Gg�R��f�{
0�zN�'�ہ���(:k7�M����bܩ��cog�ڿq��Y��R
#�H�u<z��[�]K�{D���dǏ6�I��Q�����������d���]K��T-�V��,�>3M�|�U�&�"�2�oN�eD�����%�2)m�~�O�TL�9v�E+���c����{;&M�������t����ur�Q�4R�A�SCi��%D���o|Gf֞z�&+��I}���}^���wkg��6��y��`ʵ�z��ĕ��r�RC�r3�R�V�[6�Il_��0��`���z:r(�V���zA���4�Ĝ@i�D�A���q�#f�R݀���kJ��כ�@i�ӿ謴ޛ(���c��p��>��~�YW�\Z�#�������~�JH8W��_�Mk�3���F>*MD�4�Ep�7}0�Z�4��f*��4$L�2H{�sݟ�F�#!��D-VKl�������bO]���c��%A�;���M�_m�I�B�G��Q�bH��ߢi��E5a��)%�t93,��C����B?�Y�ߍi##w��t�>�"�;ӕ�jX<�'��%��V�Ѳ.%j�Ko{]j���^�SCF��2�^�P&�W�E������:5�h���B;G㿽�{�>�h�� �L�v��.#��n�(�3[J"������4� B�$�v��h9�4�8�K����Gn�R�i�.�!*;���f*U{ӏ�Mg�>�R�J2�o�8<�S�tԘ��uY�5�1�P�R��n������{5�k��ݓ9�E;�c��B�I}b�<AK|�����&���}�GԢ��������_���#�0J�� ȧ',G��m$��!9�co�Ƣ��c=tl�y�L�t������7�f*=1��U�N�����#�y��{;$�O�Ɵ�o�0���a�ɇ|?���Tlg����y2�����RJDFV�Z4�R�ι!��IG����.�
ZhG*�Hz�T[�R�;���}G�D#���&Q^n�����mR#ȡYt8Wݽ��ne������fomB�}���=O��@�=��y;�6��Zfˢ��*�՝�}^ZW������-���L�xc3���M(1�Ѱ���Y��.�?�t�=���h��h��Z?}�Nxo3E�>�*$)�3����b��0g���T�#��ωU�������<����#�M�L'�h�����dΪe�05>7��C���&���eU�w8싘G�k#�H��
���"�?���f.�����1���5���XC�)f��}�;`��>o��{��]��q��Ӻw���c>��g9q+��ݻ��W�>�Ԉ7G�E�ٱ�]kFW�~O�Ph�����Z\��5�m\F��}�F���Ef�=��j_c(�+�>�w�]�+B���(i�uM�i
��ု���[��0�苌	y}�8��P�Uw�qϞ�E�f[q��Ǻ�<�$�&��2LU�j�)j-'x�:V�kI�Ը Z��'cY�4Lp{�aj��\�W��s{���5^V5LV��z|�a���pD�����b�՘F�<���`��U�U�E���TUA-2�q7���|��#��,�M�c�l��ȱ���G����y0���5��hsU���|����������1U��z�r�i��������1��?X���@�;�i(�
Ea���C�&�"!��i��hC(s���R��B�ڽki��N3�Oj�E�������<�%Š5�7��*ǳ��|�I�-orϞ�̞N�-Q�7*�Ea%��������$���˛q���'W/dNiC�s/-nI�D���"r^�IE�k�����ʏ�يDw�򸺺�/�]�ؒ��2�=ZeiJ�7��Xn)o�J�t\ڨWS%��))E�1咓��k�l�8.���RѢq䓧TBsEaGk	���B�Zf�J�ۆ�r��#�$������<%��ZB��J[��Bj#B����#t�b���VyNh=�K�J�9���$Z-ُ]Q�/%���<�zB����ێХ���ВZZ����dIw��6j9/��9�Lm#ӡJ-�;+�5�Bsrq�����S�G(��7łZ�FDV�r���\&�G"�)���Ȋ(�m�m%���m%�ejK��fD.U��$�,��Ȓ�f�\i#���G"���\(�En�$�����h#秖���Omg.J�#Ɋ`����6s|��7"K��@d�H� �Zk**d��h��)�&�-��o��n����l��+�1_$�$�9��\����,�h
z��������R3:[s:IG���bA2�������"�j�s�Z�F��r9K �/��0d/��}�-N�[�wZ��b�8?���V�N���ҽ� ��	�,0u_$�g��$�\��@y$�Fr�I�*�mh xA����*�G��zDQl+()Ζ��'�`����n?U�R8-g��" ���J�YQm3+�
m$����g�#��6A��V� �qR�[DQ����h3+`�oP V�d?��**\�Z���K�*X8�K�itN\M�R,q�E	:ˢ-�Fڢ1\V+d�ec(H6����R[��X$�m"�|yqk��e�-"[Q֚3��ʠ?F��$E�\IG&%�q=MKkFk͑�;�?×ޢ!��-���G�-���EC<����"Z��X���*��-ET[�o��TX������k�	��o*�
�E[hiy�(
�,�2���P�T�f6�D�ĖҾ�6T*)n�8��(��@D-��E��HD�
��e��_�('Wpm*����g�։h��B�Y���,������\�����f�g�VT�7D%�����Ҷ6����6T(R��T)�k+�	m�A�6[|�eo�,Q��&���~�NA*��V:��bq_�Sb[+�_چ�ɪm*���V��g
�$���M:KԊ�!�\[Kg	�/�)����b����8K2�_Hgi���JŖ�Ya�ˊK��,)+���q�m�wAn���`6�T��Z+�J)��l�Hqr>w�*���R��S�
NhE �ͬ�h�f�"�S�<�����S<�[�<�xr,�j�Y��)mg?�Ş<�V�'�Jme?+��w�����4�����3�|���)*�Y�NF%�mS-V�lKgE�#�+����y^�����Fm'�"[�:!ժB4kk�S�53�H˵�G�R�����PSt���ĳ��u�'PS��<`�D.��j��S��&�g<ɗ\��lr �ff��Q��$��ٝV���f5-&�%H6MK���K�L�H�0ePZii�	�+<�{-	�(�f,	Fۥ�@��k9cR��
Yg�bZ�d��h���f���r1�>�Ġ�R!���ΠT�>c��4����_��c>)��|��a>)��|R����47�Q����Tc~v2�K��9�LJs�����+��+R�[�Hin�"���
�%l���=3���|./����2���|./�����|!/���2_��|!/���2_��|��3��,�����47�Q*�f>)��|R����47�Q��f>)�g�+TVr���*9YDJKs��8�`)r�$)Ur�$)-�)�(�ٌ�=2��B��*��=�4��Ɠ���`<)�*�z��,���4�f�U9���L��4��K+*����A(�.�T7���"r�&J����2J�ܶ�9D�X�2��!�z���������/��c�\���ry>���/W�c�\���rE~Ɨ��c|IYƗ���a<J�0�y��<�/-���x�
i�=�y^�N��4����dH�y^�N��L2��y^�E��y9��|����$�����$���4����K����6No�4�ƥi|i.Gu�4���KK3�{���r���y./繼���r���y./�=p�</���r�</���r�</���r�</���8��n��z�B�m�IinkOJs[{R��ڣT�m�IinkOJs[{R���WX!��'���=J��֞����4��'���=J��֞�
YӢ{f�%/�-y�o��~K^�[�ߒ���������`�B#�Fi�R%�`Iy�C�+��=J��{�@h�0�=��ݞ�y�����]s�;�!���"��|�;�D�I�S��~C,��ǋܴ��P�~x@!�p���cj��c�̥�ƖU��7��\1��R��˫�ǕM(%�i��ʚ�Օ%�r?Wd.���	i	U�%t\�O��mp�F�;h�a�1_�1jv��U�^�&s](bn��
�_8�6���҆HM�?��k��U�;j���|^sm��Fi��C�PS}�Y5��p�G������e*i1*O(���7�̡x�1c<��k6��b�tG[�V?�����c}�$�e��t${�ջ�r�n�4����}f��6b$@]�H�������/���fw�g��x�D�զ��yB��䭕hG�F_X���uVd�E��M�pB��f��g
�6
�$��!��ڍ��H�Y{��?�}/4�Bf��&�h���z��Ew�a��h��AT�9���m�F�-')��AC��I��&����@ð/�!�ACig!�E#��LS,�	����/j��k}AL���3��1&�|J���<��o�����������&�TĜ*�v�l�%��j�F�+M�)/2E�]y�lP��L�
G|u�Hw��:J除��R����4�1���(�n�ͦ��t�ECu�8�(����ꆖ�DE#Zq������_�F��=�o9jw�Y�.����EB�(�4�����`��sD���:�۬х6V�>7�B���a?ќ�>�z0?B^ؚ>Ӥy�giv9JZ�T�����ͱ�p�|'�"3[(~�`��!��wИ�.����4��0��� �x����Bb+��yܺ�u�7�揪	�U����X��Jc���!�o��1�^qL6$Z��ԃ����P�¡���"�Y��,��P"Z��s�A�����h�7�\����yID�!-�1"Q&��7�=	��b��п�o�����,h�+��"��Y��6�)�|QH%��T�q�����3�[�Z�ե�x�9�l:Ո������ �kt�u5��*�t���/��Τ��x��}C>�ɣzun���	�� e���Bu	F����LΔ��f&:K�M�,�3&A�Jc�X��(�vBI�=(�5���kB��G�jat�`�*Lt�th���n��n�4�R�����boi�D�k} b�����6$�S@[�<w���_ z	���׺Tp�rW�B���Ns3�$�}I�ĢI��T��u/�mJm�'�{��[��h+�	%�L�9�5F����G���z<�\c8�d�H`�TR&,E�ShL�l�i�R�M�k��PG��A3��o�1��Y҇ID�~OS�)
mtGf�I"2���� ��<�JάrG�Q�XP�mN�ɢ�����36Tm�%�n��5f�hn�Hj} �=��qj/��E}�7A`�KOd�\/��)zFM_dIp�41q�k�4g��f��#�P���gN����	��0���0A ��/�h�����2C�a��QL��p�ԓ '��Ě��E|8���
y�����z�F:3b"ԇ6��Զ�d��7��Nb�!ԉ+��9��R��$,OXY
p[���3S�A�bI�J������Y27��1�I�b���Z�2��f��2�k4���� MpCuu������ڿ0�HL�FB�ux�C:jI�9��k�1zt�����3�-1N��<�T��&���&Ri�0�A�h4����E``����לY�r�E|
�t�\�@������h���:1p��L� N`8�"se��Da���&��kݻ�ݤ��0=���A:����a�Ld�P�?�9x�6��h�?F&��k��2n8����|QS�:���F+�$C��	<h��hH*]�4�c��F1AR�tf�"��Ǵw��4�pG�E~���M�	�Tۅ"3y�}2?SD�mt7'�V������$���Ah��&�0*8�h?��A��`Vs�9�Ta2d��0$�����Z"Y<�S�ɪ��!��� W�d�ddZd F�17b�R����3tS����m�K�:�M�PK�$�/	vHL��V"Df���A"ZtM�M�WBzI�$���D�i��u�I�6�A�
��VS(��dN,�k���MJ:�B]������)L@�@4�V����@���Ks�����W���2ABEM�"1��u��9�4Zy���`����7���� :6;F�L�K�D'�Z���Yt�A)�Q�ls{i ��1_Vj��&9�D#�ŢʯM��poșh$;Y����Z��Q�$���I��A�Vc�nc|I
')�"DѼ��Rmt�L%�7=�c��%���I�ֲ�P�0��n����t��:ui*AQ �3�Ah.�F�ל�G�$��t�s#@ߠ�I�<e7��hn"���+	�H�7��R�	W���|���$U�m��)�72_��<
�'gC#�h�z}AoS��4�$İZtf�0�`Q��L?���d�͝G�ҥM#H�ŀ��I�
5i&\s�I��I�RGKRa~�4�pi�m$Բ��h��,��게��Џ:�5�R�b	�����9�d�-�}��i#��-��DpRr#�h"��rA��b�b�$|��'���S�����'Q)m0e�A�44g���DRJ)g�� 夷�d���jS3�{9�HF��"!Z��&��p��P�ܒX��6��LD9�i�E\V�	F>����E"�	>�h A�F�v�����f]h����$75�	BD|�B�"hIv	V΀Qb�Rp�7D�bL��)�+�����@��w#IX%	I8i��d�O1 ]b�ʆ��-4�>z����חa�g���J��E��P#Y�%#q<���=8 )��PCof�&>�e�$���e�(�n�:g�y"P#Ҝ��8k��Ȓ�$
2t�r���Ta�M��G��BJb���1�.I�1t(I*��ט+k
�%�5�5M'V�5n�x�������+�k��S���U��Ǟb>�rl �_[3�M ͘��oJJ2�+4'�6Q3bOJ"�D2�'H8�r���B�z�ʱՕcG��);��<���tFX\R9�r�)Tf**Ǐ-�і؋iU���ф����	�U�j�5ϩ��H�#�C?M�Ӆ-dK��*
G�KӉ�A�H*nIc�����{�(P��f��Qj��!�?�j�Z_��y���ɖQ&5��%�=���Z��2W7j�	�� �&p)@S� ��D��X���R���>�x���&��r�z�e��=D��$]��R4FVO��b��]�,�G�2rvU�Lc�W ��O?�T��)7ݍ����8��X5O���?+�X��� �jz�A��)Y�қ4�/�ua�$#�V��G��.Yc�@)�V�I���L��� ~H��ccDd�&����7�$�u3�_Cᰛ��oo"C�s�M���uM�$@�^����^'��J�S_�B�����m!��v{g���b���®O�X���®��=�ԓ�6�t[�t�)�?��@�t�L_i˻`e�GOC(��ib1eM�&7��|�b���ё_����r��mk�b�k��F.J�f��9TГ@{'���Um�3!���@�h��	B�Q�8�W�0/A(JƔf�3�;<����B$��4W�_&F2i"�X)ZI.K�:��IỞx%q��N��D�5��4��i���!����z��ݑFjj<�����M�Hr�IO���"R&a���,l���m�1�1�f2�$%�;�"{)�/1*��cˈ�̶��WU�F�$+a��a,����ԝj��$n,�`p���~��� =�אp�Al3�����x�f�}��f�k���X0eZ�N�4��S�R�"�P��ĊzB��5� �F�Q�0�<1ʧ���r&Q�h3�����!����a
p[ J�y��zRR�δ�&(*�3�Ј�ð�X���Z_r]X�F%���ϟ��X�b���� d��3��h���X�L�H��w��@w)���pS��7�<�C�X��Fj�B�M	l�ť0uãy���X8�ֽ�8]�ܑ��6`�?�����%$(�Rs���*wZ��ZwL��=��=��|FK��@�A�[��wM�e���C���C����r��|i�M�	��
�7A���a탙��h�"	��-gD�h��EL{�a:���?����`����G���<���O�F�>����K~�)I�H����Ր�w�:Po�Y�C~��v������G�C�ߎ�N�]3b=�}���ۈW������X��4����U�3�hSf〭�Ƶ�L;S7Sg��܎aj�k�g�OO|��ȩ�~����G��%��q�Q<�\zbf��{jUz���I�&|Y֎��)�n�t>���/�wܫ���I��v������h�6��?{F��s�{�8�qR������H4��w:�ed8ֶ�7�(��P�v�67���Z�+9L�Z9d�l���>���)�=p�Ǜp�.���Qp�Y9��8�7��Op܄�W8��'���_)}��\\Uiዼ� ��ߢ�ѣ�˫ǖ��/O�)�ֿ6Fgy"1��fT�h���ʱ5㋵��k�����������
���,3�5E��������[&���-~ȶ�����]�3N�_w����a+�?�2~̖����X�����+��ǯ_���q����~�U��m���wl�o�v[��;���Wm���b[�����w���u���y��m�h����w}u������?|m[�����?o�׽�-.���뇜�-~��O����l��p[��c>�O��x����K*��׎����O��G�r����~[�v��%>��O�w\�->�9 �ڵd[|u�-����n[��v�ck1����ǡ��_���Q�J|ǧ7�b�����o�t��C�2��7�M؀v���~~>�	��P�T�t��+��/Y�L���^���>?g�3�SO{&���gh}e��Yo5\9���U������w��_q�����o��l�?�{c������1~�=��;��	���1�t���}�n�pЦ��6��߸!ޯݦ�w]7�'��~|����_��T�0���~�W�O�}���]�S�X��?w�a����^�l�(��症�|i^��5'_��wQx�a��gT������s�\��</���y�q<��E�n���{p^�q뼰�(�p���[\v�Z^}��p���Or^x�u��/��"�G����ڈ����O{����|!r�5�o�^Qck#����Cv�W1�s&�3狟fL�g���������Z��އ����^�M5���Øny�1=�Pv:�fL���{ΟLL��˼�\�s�r���#����x�Vқ�ͅ�t��6
n�3����1b��P��~q�<�י�ho����z��o�t�k���D�v�ô�^��m`�%���J|F��N�2|6����z�Z�s#��a��K�����wtf��9j�ɐp��6�kmv�f���Əc1��Ǹq���f�� ���Sό�Ye������A� 3��ap=���p�23Q/��j�8^S��BY�!�"��A�&�mm�(#��3�Lg��gN��6#�Ŀ(���zŝq�	MͫH(5���y�D��q]k�	�"�����'�ߐ�W_dL��3Ώ{�1݃�z|�+��zy���鉕��/㼴�.��c�Lz���Dڳ3�cv#)M|�Gj���:���4e�n�;&Eڙ��������T�Ġ����}�b���}j���a��=b�o�ȆG����?.�?~�|�K��ƻ?|`�g��_?��n���I�zo*�������|��;ל��_��󯑮�,�q᫓�>h�����[���,�w~�ESV}3�uO����Wˎ�/^��?�[�a2�6cz�]�4�e���g0>��|,�c4�#v�8s����5Uw�D��x��e��"R��53u�^�̋��/sޭ��s��ң��{�/q��%�2�˜�	#L����kSI�8���J���C'	�}bT�8'��zI�vSQ[�_f?�_��d2=�����tᗹ&ӥo�����wc�����tyL���K��H�r��P����L��D�}s�6^��ͷ��6Jg�Lk��wr�Q��3��l����9��!�,D;����3�ݖ휆�}�foG��}���*Rho�V՜����.5)V�"���ԾQ��f�)�I��;�:gI��� ����$����eH9Q����6���~��7h���h=׼���R�u�����/1�c�g�7i�e��
:�wz�o�8&�~7z
�zZ?����1c>�t�i���v#��߈�
��z�M���1-���[��X
t�Z�CϧQ~�+���ٖ��u�xJ�Fj5�e���Ǵ3��cj��d:gc*�L�O[��>�M;��90��L'2�1�L}���'E�ҹlF�~���0�I����s�GC.'�_���Y�L_���̱��>��%F/�5�Gy/������OƁ�)e�34���Ɵ�0��vV�2 �Jʫ�Rz+��+�R���?��7��6&�>g�R8q��5�T�R��vH�FM�wi���z��]D��i���T��m.ˑ�6�<v9[�Z{W���m�l�p~��8��lo2���1��c:�w�T�cꈹ�7�LG���}˘:mbL'�ʘ�mfL��\�zO�����i)>[�mZ�kt�g��M�ǁ=�)����d{����%;_=O�L�4=]^I��w5ּ�9�3��4��ǏƧ��.��B�j���/Ï�hTFt�	=E��>��o%u�����ô,�F���S�/�R?�	��h*�k��J��>)î�w���|#U<�m���h��F�k�(������ڄdK��M;��3��l�u��2�;=���E�g}9i�絊�˟�����Lo}ϡ�47گ_x�'�[�"㓊��@�R��dj�g>��܈i^�D��P�G!z�?8�̿��)7l�=���?�L��&�-�L?�8�H��w/�i}�e�,ǽ�L����ێ&䨚���Xc:r�P��q%Hu'H-L��e�5�ũ�Τ�j�-+B�[Gр/O;5��=#�\�S]˼'�Ǎ����JZ��;�T��ҟ�����X�h/иF�����do��W��iN'��ĠA���Um2��=]�*�}��d�����L&3>�	�Ȑa��D�:l�����Ͽ��N=Y�V:��`��cM�a�������*��
�@m^o��5�i$��� :voOt�c�th���{��6o-��?����0����FI�|�h!w~$D�~-ͪe�r�y:�7��;�d��kc�24}��6'x��4���r|��� |߿bJ�1n���2�kL�� �e�c�1ym
Lי|�(;��S[������u�<���M�6b���M/�s��4Aω�Jƕ��˞��̿vy$9v�G��:d����xW׌�n�^���V��ᦴ�tW��t>�&SX2�ç�ؐ�M����L��sU��0��)�	�U M��_f�jZ�^�Q�d�� |��Y��'��L�1.R���|~�R�G����e��+��˪�R�T��,��'g��Y�T���e2=��h������jm�֫��*oS�?&?��K,2��C�##ϲ??�����uR�|k˞�R�~��F]�|�/�e�v�	l�s����y�~�ֆ	��O�'�#���ǻ��S�t���������j����V���<���c�W���zuuf����t-�*��T��1�j� &�w\ 8�KmY4-��I���Π13U�O�N�aN�g:��h����>�� �T��c�٥�[L��=�;
���FYֻ�Ԙ#�7�e�����sV��g�^fM�����Y���n�琉���{�>t���+��j����5�/~8}3ק�+Ǽ�����w�5��o�}�����G���ڶ�ۆ_P�6���G����Y��ѓ�|��{�(c����v�T�o����F\~��/O��`@�~z���v��e��t���ã3��Q�q��W�|��'�v�p+o�Zy���/�{��?o޾Vn�l��{'����;��=��ߝ����q�������syݨ����'>9���7}������/�z�Q}�Ƅ![�rq��,i(^2젇�?uhu��6���s#n��ܟ6�q�6������HXXZ��'_�����/��9zq���_۹薺!�|t֔[+/}{Pd����;��ۧ�6ͷ��@xT�_�=���}*&�uٍ,�|���w������O<V~�[�G]���v�?�L{�!�̴^qp�������7������k�l@�������G�p�����|qhem�{�>{�';O\�N���W�=���?��ݖ��^����c�~;}�I��s����⌛�Zw��˶��<x�/���)��5K܇���U�?���Lp���i����������g�u��x|��<���&�1]���L� $H����h�	b��%12	��H�1ci�Q�1�-���j�{i����jW�ƾ��A)"��s�$3��>����K2����s�=�}���Xm��[�7��|f������gp`��E�v=���_�4j��ףG��?>4�믯\?~����1c�R�=��������}���Ϟ۵�7n����W<z���O>y�����k����O?�{))��%iiL��o;���>��g�z�#Z�|uJ��ܽ뒲o_/C���>����˗�߻ySsa���>qb��f͢��vи�y.���V�v����c�����Õ�J��zy��ue=<J�)_�e�iӖ��p�����z��������6���/Y�j���e�766�R�i˪U��5ꇟ^}���+|ڻw�������1$���~饷N_��>���V�9�ϣ���r���m�~�Z�Ѐ����jLZ�v��\;���źwo��[��LjӦ�����,����~��ԃ�o<t荝��Ӱ�W_]���A�Y�;�\q|XPP�r�����jfݻ������h���+t�CB��]���_|q񓨨[�V�z4-44�Ļ��������t�1�[�߼s��M��N��������ԩf����/�lU޺Uv�##�������ӧ^�
-�_��򖸸�->���]��kZ�R�v���]��߼)Sf�ٮ]������:h�_�T���ʸq�^Qy���z�:��ԩ�]j�֧a�)���}]z��9aa�e\���6����'d��3�6��^�X�t�o33�g�;��+1ƶm#}J���~�n��������a��K˷m����Gu��v�y�����ق��~�R�'M���W,�wwժU�?G�\��Z�=v,����#ݾ��܉#~�&&���۷=��w������s�~�]��F�7��_�ݘ8qv��uGl�4��������O���W�j�<}z�d4~ܾF����qz��ͧ�X,���y'�ܘ1�&�o�i�u;��ռ��%����˖-�mȐU�-Z�}�����/�*͚�ޢ��~m�U�_ٲ_N�?�:;7�B���U�\Б��7~y����s�A��n�d��!ի��}����de�}�@������4���ٳo�Ι�n��+sK��Ӫ�)S)a��?�_��lf�N�ft���E�ּڤɄ�^^��Z�f�}��ܸ��+�� �	 , � @ `3 � � �  W �K   �  �  � - �  � |�l ` P �
 � < � � w�� �6 � � H ^ : . @/ `  p h h � �q @4 � � z 	 @, �  X	 x � �� @K `	 � �  � ��� �2 � 4 �  ?  �� @     o ��� �G � �  p�7  5 �� �5 `  � z  g �� � t �   ��� �N �8 � �  � w `: p � �
 \ n � �4 � �[ `  � g�t � �  U �� �H �' � �  ^ � �  � �6 � � � t � �   � �B �0 0  L � R �� �� ��� ` p � � ��   � d � � �% ` 0
 � � � � h X �W �� @ `= 0 � �  � �� �� � P � � d ~ �1 `6 0 H �  7�  
 � L > j ��S �,   � t v  _ ' � � ( � � �{ �! �= � P � h T  ~ � �� � � � ~ j �  @7 � L � � r�i @% �O � � �  l �   �r �^   � h � L &  o � o  ��� @  � ^  � �� �� �x �7 ` � H � ��� � �[ �( �	 �= �1 �) � � ��� � @= �% � � � � � ��� �X � � � � � �6 � � > J  �  �< 0 �  d ��   P H  U �� �( �U ` �  �  ~ ^ . / 3�h �0 ��   � �� �    � l �  ��� @? �  p � �
 x  t " �    � �   `* � B �� � @ �
  � � � ��; �& �g �O �& � � �[ � `? �	 T  � q �G @ � � X L � � �  �2 0  L z � �Z @C ` 0  �    �  � 2�s �+ @[ � � p �  �m �� �7 �P �= ` p	 � � � Z # + p � � F  1 �m �o   x � �  � �� @S � � �	 � H �i � �  z  �  � 0 h � � � �+ � � �  -  = � 0 H � � �� @. � (  N s�� � �: �6 �   �  �� � `% ` �  [�+ @' �  t  M  / ` � � T  �wA��B�_��ρ��A�����=�����.�� �c ����_����]����f������@�� �?���G��!�� �����!��!�/A�/��7A����o�������;��)����(��Ð�� �/@��?�!�����R��@��V��� �_��/�_�*��Y��������S!����/�_��s������ ��� ��)��x�����ɐ��!�OC��B�W�����1� ��P������ ���?
�o���?	�>��B��5�����!�wB������?�1��0��r���@�gA��A�?��_�?�.���O �A�O��/���&��������A�O����� ��e�����[!��C��A�׃�������l�����@����σ��7������@�_��O���������>������!��@�g@���� �5��&������B�gB��C�!�} �߇������� ���3�g����m ��A����/��1���(��?!�Ր�k!�?��������[��!���������4������!�[C��!��A����%�����C��!��e �� ��A�O������;��]���m������A�������-�}�����ِ�� �kA�������?�	��/�����!�����A���
���$�������3!�A�π�	��U����oA��?�q��պ)��T�t{������K�7�����]?�����#sf�����u{]>�������Zt��n�wϬ}�[�_�������A���o��2���ְ�V����]����������|3{A��ݒҤ������i��]L�̉��N���_�7��2����~�1��J{��|��O����w�J�E=U�6~¹�o|7�����4��	7�{W����3#���V�����^;��˅�5����u��x��n�묝o-�����o�[{�g?��&�z�⌁��o�z�O�����F��+���߽Ėc������G�4o���[}W�x��+��d�J�\m:���b�.w�<�;�}�w�}xڽ���%����9�>�ucw*��~t�`�����u�؜��9���O.��F���l��W��'��rr���;ye�ά��ZU%��Jy�ѵ����|3�դȇem�R[Ǵ��X��M��/�u2�0��K�9\�eӶ��^_���/���x����MK��kȩ�O^��c��*/|�k��/��:׹|�J�ʖ,S�_KƷM~����_��߬���ɣ��E�7��:��]u����l�2,x�S�[:�4~o�]�~��g�p��kǛ����k��>�:sW����u��ll��ݽW�e��rd�e/�8�C�2�z_��~�P�+��r�/�����5+��ysv��ѡJLr������v�Ȍ������G��n����?{�L�?�ϭ��ۭ�6n���n��e��-�3%lh��¶y'6HM�܍����;�M�2���Gk�������͢`o����ǯ������zK���w�����^����`T�W�+Sjn:���W���_KNv�����K}i��?�}���;�n����->�f���*o�o���whM���7�v�x�ϻS���Vz/���X;��&b�W}.}�vv��u{&ή�޸Ɔ����Kc�vS�i1����qJwl����^}?�H�,�t�����9�Vz��?�gnv��/�__?dO�������um��G�����~>&��h�5�����~5�l��>�d����[�1�hߺN���V��U��=iӅ��B�Yletl�z����3'~��q|L�����r앟Ǆ�h<�A�I D ���� �M �k � �/ � � � � �� �4 �] � �: � 8 �  ��U �. �/ ` � �	 4 ~ ^ �  � �D � �4 �3 P	  � � 3 �� � 8 � ��� @? �2 �6 � � \  � @C � p  � � ?  � �F �� � `% � 8 �  � � + �W   � �
 p � �{ @; �;   X �  F 6 � � � �  l f ��L �+ � � 8�S �p �   x  �  ��� @< P 8 � � ^ � ` � �  T J ��� @5 �4 �- � � H z �� �r ` � h � N  �5 �7 �   �d   ( � z  � �� �! ` � � � v  U � �? @ � < Z � @= �S � P X  �   � �  ��/��` `5 0
 x (	 � � � @ 0 �  W �� � �( � �= �  � �V �� � � � � � / V   � � . U� �T �  � � � ��  � 0 x � ��� @ �  � :  � �� �� �  � � L � ��8  	 � , @G `, p � �  �  F � � H  > b�7  - � p � #�� @O �8 � � � ^ � e�4 � �  > � q �� �� @   �	  v f ` �  � � � � ��f @ 0 �  | �    �! 0 � ~ \ �w��� �6 �- @ � | $ 3   �' �_ � p �   � @_ �< � \ � � � �; �; P � X�A �Q � x  d ��e @' �   � �  / �: ��? � � �   � 8 � N � } �� �� �_ �� �{ �N    � T ~  � �J @   � � � x  ��� @= �  L ^ v y �M � �
 � � u �v �+ �J �e   � \ * �  � @< 0 �  4 � � �a � �4 0 8 � � K���} @ P �  � � �   M �� �"   x � L � �� �b ` p 8 H � �% P � �  � � � �M �o �! � � � � 9 � �   p � �� @ �7 � 0 �j �   �
  <    � � . k�� �8 �  �
 � | � 2�[ � �9 
 l � � � � � � � 3���� � �������_�-�0���o �{@�@��?���/������ ��A������������:����W�_����� ��B������?�����}��-��7 ��@�'C�����#�����k!�7B�?����?��]������!����O����?�����!�gA����_������;���!�oA�GB�'@��C�������������B��������������C��Ӑ����A����w���_���3����k �= ��������2�.�?�I��W ��C���������%�)�����:�����@���_�����W!��!�/@��A��@����/��/���=������!�WA�߅���� ��/��ϐ� ��C�w��� �?�?����w����� �OA����� ����K��r��]!����_��_��m�����s �B�������� �C�� �!��@��@�σ�o
�?�9��p��ѐ�!�wC�{C�K������!�GA�_��O������M�� ������7��K��� �B���o�o��σ�?���#��T��J���!�;C�������'�:���R�5��}����?B�����?�1�+�����ِ� ��C������c�����~��� ��!�� ��B�O�������֐�� �+B�o��o �o��o����?�����1��p��C�s���������A����E���k���1����+�3�w��M������������W����G��������]������s�u����30��Ocv@�Ƽ�ޓ='3f���X�P��铙m��2W�g������������/�EЧ1{�W���c�B_�<����~�����~�9sf����>������f���"�ߘ�Я3o`�A�Lo�쁾�9�8}8�5s�@�]za�O�,�k����Y�e��0���d&A�����0}8��&�'�_0�a������z[�8�j�0;`�B�J�l�����$�a�_f7�g�11ka���Y	}9}5}?3f�蓙k�#ӣ3�a.�l����s�%�b�顙�0a~�l�� 3fN̔�O1{`�����~��
�*f@���0a��,��3�E��这�1�a�,�9s�������ӣ3'a�Ƭ�y�f)�L��1�a�܁�s1��c��0�a.�L���,fG̶��03c^Ǽ��ft����������A����E���k���1����+�3�w��M������������W����G��������]������s�u����30��Ocv@�Ƽ�ޓ='3f���X�P��铙m��2W�g������������/�EЧ1{�W���c�B_�<����~�����~�9sf����>������f���"�ߘ�Я3o`�A�Lo�쁾�9�8}8�5s�@�]za�O�,�k����Y�e��0���d&A�����0}8��&�'�_0�a������z[�8�j�0;`�B�J�l�����$�a�_f7�g�11ka���Y	}9}5}?3f�蓙k�#ӣ3�a.�l����s�%�b�顙�0a~�l�� 3fN̔�O1{`�����~��
�*f@���0a��,��3�E��这�1�a�,�9s�������ӣ3'a�Ƭ�y�f)�L��1�a�܁�s1��c��0�a.�L���,fG̶��03c^Ǽ��ft����������A����E���k���1����+�3�w��M������������W����G��������]������s�u����30��Ocv@�Ƽ�ޓ='3f���X�P��铙m��2W�g������������/�EЧ1{�W���c�B_�<����~�����~�9sf����>������f���"�ߘ�Я3o`�A�Lo�쁾�9�8}8�5s�@�]za�O�,�k����Y�e��0���d&A�����0}8��&�'�_0�a������z[�8�j�0;`�B�J�l�����$�a�_f7�g�11ka���Y	}9}5}?3f�蓙k�#ӣ3�a.�l����s�%�b�顙�0a~�l�� 3fN̔�O1{`�����~��
�*f@���0a��,��3�E��这�1�a�,�9s�������ӣ3'a�Ƭ�y�f)�L��1�a�܁�s1��c��0�a.�L���,fG̶��03c^Ǽ��ft� @�HHA�IoID�|�^�������^����ޑ���>�~�ޙބ^�����~����~�ދ�~�ޑ������ޅ^�~�~���>�^�����9�
�4f�o��=�a�s2�`6A�K�E�\�~�>��}/s{FAoM�NoJ_�܀~���Y}�zez~�?�(�e�3��I������7�C0G`��\�����o�ϘA0_`�A�,�����:�f�����蛙cЏӇ�_3���ߥ��d�¼���^���^���zKf���A���Ӈ3/`n�|��3��/�0��e�ì�� ��(����̆�{�}0K���ev�|��fÓ��З�W��3#a��|�>��=2=:��"�&这�07`^�,�����
��̶�0#a��L����� ��י�0�b���Y3�/̒�90�a^������Q̂�C0Wa����?=:s�h�z�0_a��̄Y�� ��/1c~�<��	3�r�4�0�bv�l��33�u�K�Q1aF�j�
3{Z\���v~۴A�
��*�%p��˰����^�^�	;M�=�a����+�~����j��F���Q�On�qO�{]��K���?�b����a�ުUGU�$ޱƿt��UE��ު�X�5�kTK�Xy˴*Djq/���]�9���ÚZ�̀��D��X.U�Tl�?k��o��=�E?@�/������ٸb�}�����~�▗��߃�'�[x��{��"�.��,��9Eթ�=�׉�')G�wJOzJ���6�OiH�:��n���4�Ž���}����^[�T�8��;�&OA�t��1ʽ���.n���]�]���CŚ��<����_�k�����DD>��_c�v�{����Sٟ	ff�|g}_�\�Q�����t�_������S>��w��z��{�?P���|6D-��s��;\��9\�����ُAA[󸚔��#�=�#�x��B�q��3{?�?��8fc0և;T�A��':b$PR~Գ���Ӣ�/{~���_+cH)��Z�+����ۇ�><�()^<�����[�}��q�6~G�_��Y./��c�w����K���{�Y��i	��h'��2<^c�m��\�޲B.w�J�z�*��O��<���7=𯗸�9Np�o�� ��,I���ϳt.��Ew�Mg1�D?C��W�t�g�8�}���z���Oxwo1���|b�����B�6}�������|��������ۻ��<Z�����=��<˼����y�|��%�ܿ�go�_������ŕ����E=�>8����Ͼ���O����e{�����7F��ׄV*zO�糖�x�<�_?�����Z�������q�<��E�K�O��ߎO*��=~�r�fw�޵��w,r�(�m����~�G�ݽ~���q�:ܞeH�y�bU�^y���[�$���R����g_�����0����޿�_+~/k�M�]}���G� k��?�տ��w���5���p�Z����V��O��d4��0dԨ�㬳�d�ḙ�p>���<�k�s<A�i��x����P��'=��y��-� ����]��?[{<�s����cO������dT�y?��h~���?Fa�[$�1��*����7aJ��S��_S҉y&^��������S�P�u���C+�ٟo����i���w�R}h���}w~{��/j�[/��?�Շ~.:�8�A-���`����'iȨq�쏇{~�+�B���J�=�	~�y��l��C�o~�v�)k6�.�0�	d��{Nq�����c����p��)�}��e���4T��e�E�{��m\w�؝�޾~_����蜛�k�F�z�>�SE��@��m<O��[NT����ܨ��l+�հoK�u�݌�g�Z�$]8D�qu�?��Y5�#2Z99�WN���Qi�����c��ۥh�o=$N(��B�����$F<)�O��Z�rZU?���S^*�9T���g-���ዕW�:.��h%�Ԋ�*v}�	�tO�S��V�+y|}*��ʓ��vQ����]%���س��'k^�zѢ����O^�ѷU�>��Q�\~���~��҉W��n�����g[��5���{�O_}���ū.J�9����g�1J�]멝�X��ZE���!��sn���y��XTힷ�'T��U޳����������ψ��syOk{ٻv���Ě}��ݛ�ʈ5溽Do�?ʹ�3ցG<B8i������%�%_���Yn��M��<9���*���x���E|�|�.��U�����J��n�����V���{�^Dg�G�f�3��3p�Sl��C��v,���[M�]��~�Ӳ��X����}y^�χS�����_�&�3��f�����?�t'��=��?����oR�}��;�/������n�za�����,�m�j"T�}/S��_��g���sގ�c�����/��V��rf���֜�a��������\y�s�����:�/���gU�U/�����$����)>Gv�ʳl�Ųq��o�y�}y��<)���?F�i�>;������_m�o���<����q��E�׋�7q��SO�f�J��g;ٜ�}(����w"^l�`�?%~�BYnk������G+5,�c�s_��;R��y`�:�3xQ9ēʑ�]�Y@7U�o&
P5p�Vâ��M��7�2F�^*f;����v;t�	���8_�r|�Z]�Z���͔�0�o�t�
����{��9����5����5w��*nn�%����ǯ*.���|%���Jx�v�{��RE�3��UԚ�_7`O
G�^n��Ϟhڿ9�qD��a���7/<yl?ޮ}�W�����ׅ�3#L%��c	����y���:��Pr�^����B-Q�Q��k-� ��� ���h�����������Һ&���bL��W�=$)^>O;�;a���	���9|�1a��;�^��C��C��*
�彨\��>�� ��ݾ����휓N�.���g�^n��7nG����	���s�ϑ
�ki}E^�G��Q��w]�Ϻ����v����	#�:B�0Ө׌�G���v�������b�u�Q|���돯��n��k	a��X�����D9��)��p~�ȋ��l��ݡ���[�q��jċ�r��ٿ�2.��_a�j�����g&�M궺℉-5҉�/���Eɩ����S-1��	\����u�|����C��,��D;s���3�Y�Y��q����Ϻ��<}���}9��|��7n�o�%�������+�J�m��@�oY{�����fџ�(��Ί��{�P�8��Gş��î��o.�_��|N��;��k!�����z����ٯV9�֫pI���쳞�Z�g�{6���}�ޤ��[��ύ����Ԏ��gW���9�P�.�qO��V����I�1%��S�ߌߝ^S�����uli3G�ſ�*��[�ܙ���sQ���1e�߫�{���z/^�P���r9���o{u�f�����=Ӌ�|���y]�p�E4�5����rQ���㟫��zYE�}jX�`�"˺�;kG�F�Ck|��)�q��p���(���9^�
�_����>Pp��h�xD���\t�W���UO��*.�����Y�4z�$^��khb�kƈ!�����Td{=O.��|��lQ�F��)8nϻ?ō�����}x�=����ɵx��uU�l�q��~�;}�XK�g�쇇�bP':K�����(�^��5�>]����^��=ژ�0d��G��,QD!�:���.�C�{~���#�e~�Z��x���$�w��3{z�.K�z��=)}�e�lQ���8�	�GRԥ�����]jg��O�?ŏ���[����-����$�~�|������䂲d���k�=t��΢�Г��4Ǳ��R�'��z1~�K�Z5�2��Y������>��q�ꢎi�^��E袶��~��*ի͜�ig^��y�(#���w��$;&�ۓ�s,и�YV��Wu���ۖ.�ۻ�k7wQ�*tn�I㷀�v�U�}�����?��_���ra�����z�Yڞ��%=On�P�7r;o��>-XJZ��`�|�\>o�,G�=�	��O��$�\7�ۗ�">y]ܯ̣�RJ��4��	��$Z\%=F%�5)P���
��D�K{�i�=q����+��z��4����Z���UE��׳~÷Q��*fY�x���I�@8�c����%s+x���I~1c��N���3cB{/�W�f��\���E�����+�����E�7 �EݰY�I��(�#�x�$AC{�ܠXz�|�n.�(W�sQ��WW���܎���<�:7S�xy�z�=���4�����5����d��_����e��ݰ�u#�5�Uj}�_��a�NG��W����fI��W�uU����Ȯ}�U/�_�1.��_�D��;�Kt������m���=�w=�O��ڈ�c������E��1lл��[�T*�͔�<�5�Gg�m^N����=��la�,�r@��R�ݳ���B�[$��4�>�޾��%6�TT����+�5�p7s8~z�ý�����ۃ��e-����1��R��J��ը��1�1�m�;h��J,d��R'b0�|CQ�UI.j�o^Z��u��Wjڔum6���J�1m{�����'�������b����}�+ŪiƲ:���k��$kRm����w,��ht�(M��Ai�-z��M��.�onoɈ+��(b��9�T��<jA;�ڼ蘠�j^7��f^7O��&~�?g�������)�G#��y�	�Q��IT��|�Qe鼯J��k�}k*���3R�*��QE��M|�m�lb��y����\�J��>�53S��\�`(����:Q�h��\���i^3fO���ں�u�c������9�3�·o�-ʜ-�&�(��N7�;�GKj��`*c�+�|�O����Sk�L�����ǭ��F+?�bf�?�����6��� /|�XN���1Vy՞C�J����󷤊�w=�C+�E��㻢D�:�˿ۈi,g�%� �ض��XB��7=�;��>m��h��8\�j�8��_Li���^���nJ���~���
��݌�;�X2%�Gy7"/h?�LL{�y;tY���f򱙼m&O��lt�A�|>�U������N�X���X���Ic�Uy�8�\-&�㨖����y:n��ͷ����&�Q�f�r� `��<NQ������tvâXK��R��V[��o5ή�n�it��w�+�-�nfup$���V�wM���I�}X3.�2@��i�73@�ʰ�h>��!(Q��p`DTt�^,�ݻ'����q>��X�Z&4���g���wby�Y��ƒ���MW��+�	�b�c��6/.v�'�X"<��R�5��I��/�A��ׇY�����=@������~+���F��z����{���̚��H���g���&J����l0h��l-8ZpѪEۙ��cm1��L��d�[�o,��k���5������)�'6��r�2u����Ѥ�Q�l���A�4*���X"��j=u����rb96��iJ��[R��Q~��\���!�itA�ÏrL.��;N�O����L�륇��2-7�an��hC�j/`�p`gKÉ��ˆ���5�O����Kt��^��:�R	�f/�*~^?������7�sW�M�,anQGL_���{�\�魩�(���� �˶��YSo�!��Jm �u�`��9Z�Dd�7�c�o���2?`�#�Q����w��a#�^���G�v�G����M��1�F���c��0�y3�'����Ul��� L{_����s�0Mj���2�Se�b4��6�>(&[����Daa���#�:����<6:;��(K��X�tj��e�]ה�h��\k?��KUO��ز��a-	eW�GY�N:nZ���ۛ��́�	n6S�<�����g�����fM>q�kl��Y{բ�į۽��:�c4�6�>���D���E�k��f1�a^��=d>k*-�����]�aB����amژ�-����2�%�k}�a)�j��3�TrX�j��u��#Z�G�����?��+�>;.vXJ[�i�</p+��YS?Š54re�i��㓨����ļM��Sq��x�MN�J�l���ZF����։����b�@�t��nT5+��}���rN�(�d�ޔz�`��Qe�KX##��DEQi�%z!����Fw����:1�"�Z�P� [�/��QM�������d3U���+�$f��b��(�<�G��i9J�7�vQ��[�t���6_�i�,���(��� ��C0�q�M���j0ai�P�g��P ִ���Tw��)֢�6k������,Z?�j*���=��3�]�)s�9�V��~�UD_�A�d�������A��+���(���+��(������D7w��c~�������P�I�2��e�k*���-��ReO��rFe1+���1!uM�|�AM���+(j6�%7�1�0�T����>�)��J�3�>��|ӰX6��<./4�Ҋ)YnY�Ǻ[n:ui���Z�Y��Zp�Ԫ'�%E8�\hu���r/e����S�����[��l�������fj#�"��X��l���S�)�f��������	{y�Dմ�'b�mk�����)n���q��a���N��8y�-b�b����c'Fb!���ɽѦ��x��G�Z#��<7�i��R�U�#���u5U��JpƔ*�*�,V��<K��'����V��� 鞆r�ȣl�-�VP��Y#�\L
S�F5k���ƒ�j���������ynv��e)8r�'����c�K�
��M��D�C��[dr�N��l�L��葕=-Cg�����/��#�?�9{�P8>�Z�/E�3��w^���it�<#o!�sʻ�=k�8�ů�#ƸmY����|BV�~��L��3��ɕ��(>���l���y���sz���[؝ s�2E���C*����Kg5�6�-�����vp�\�:K�Q�1J�4i�Q�C��B��X����ԇEz�.�ݕ(�h6�{�=$`Bϙ0�)ɗT�N��u)���O�o�hw��x����vM,�O����
�o�l�BQ��vͩ�M�l�(6���tО6��槛���4|��X7��=��i,%��tQR[�	���S�4�<l������Gf%ͮ�fl����yư��X߈W��X�?�L���[봀h���p���JccU�FeL�R6��ʎ߇=��/��.�2�Xv�&�-�o���D�U����*SkִLc��-�L ��o�mΦ.�˙����/��ke �P�j���}&�v�c���^"g�m�V��]
�,-����<T��o���f�:�ւQ��Ko�:�V�kt2_(�fڼ��:s�Q�4t�U{#^|g�vKčxs���I�ryP��o���,V�5I����2|��rk{�\W¶�4���Ƣ����q#ϙ�L�v5յ���(�Ae�o���U�]-��h�
]���6��{�Tu��9�A�Ilu}�[)���4æ����햎!��ʁ�'hϰ��J��Q-��~<�>*��k}G����c݃����]4~�Y�=-����JZ�i\O?H�L٦NIk�G����5U?4Z�?�+;`o�Ux�v�J�m�ޒ�N�F��:�R������C��Q�������D�&���᷽U�䷊�n�k�]W`5@Ѕ���R?C ��-z�Jv]h��\�<߇KfG%j�����B+����s:���F���sʢ���Z��VqA��RI�V�))�ێb;�X�.���cAy�noEOC(k��{�#��c�=�1��6OeS#KTH��u���&���[�J���7���P`��w�y���i�!&/�l���f���X�k}��a�\T��.�m��/Qz�V3��Zy������b[�F^	��a��s��X��U!�<;:ƪ�8nSě��s�!� �o(�����XN��� � j�[z�\�"(���,36N1y8�!N�o��������*Ӈ?}u�Y�'���v]�s��1�W�x�Z��U"D���Z�j��>~��a��j�@��m�`��j5�F���shٌ_�vjt���pU<��(�?K���2J�*�̜z��/O�%G�a>��
z���l�y���ů=�>���{:��9�V9��8��tj�D5���d��Y��ڛ�r�*d�Ob#y�H-�e,�K�vF�c��R"T5-���u��}����l��Z9��.F�����R�1>�1��b�z��Kʁ4R&�/ߦ<K�㰾�X���~e}��VF�mW���o�>CG��t77M��l���b_��
�)�n��w�C�v�V��v#;#<�jY����<��n��^jJ��Zk����<�.go��-�lT���PPK�hϴ��i�4�t�&�.s�g\F���Y9�s�RҼu� �\�Weg�)r�	�1R�d68j�n�ŋ���i�9�5H���e�B�P�3B5��G֎vM��_ň�~<��<�O��]Rl���KI�V1��i���/{�a֕�䜬<���e7nT;�z�w}����r�
�Dj��2������-;�⑨�g��/я<Q���J?*��l,�:'}�R��8�-�lv5˶���g��\k�K��X��X��W6�]�ׁ~����5�?J׻�h�kGS�A���m[P����p(���'�r����GJ�&k�#����@U�G�d��o��c|3Q�nd��zs��v�C�9����0���a��a��rSz��6�?(zD���[y�[�zN��hv��Ts3�=�M�H�]S��[�l�q�_l�}��rg�Q;YBQ�Q�1����~�5s-�>��NI�B9���[�5sb�^3�fj��-ț�T6�'�#���-&ok��.:i�}��J�4�G�a1��yI.zr"�0�t\I���J��2W��Sܞ�7�
�Y�N�U��E��J�S�'��Ҳ�0��3���L+�n����{�@y��+{�Z�b�[�nSٔ]���D�����Ai�&������.�4���cS���b,|�X2��k�
:��h9Z�P75����U:)+�%����#���<K{��|���]#ua��&)�]/'��{�qS^Co�j�䅯9mY[���Р}e<m��i'yY]�k�����KA9:�)O�~K4��YM4{%�m�~m�Ş�BK9�g�Ҁ<,�/�7JZTf��P9�t>K���ňҹ��Ans`��ASxK�q��.�7�D���`G͘ս1w����{�G�Y�!��uRr��:8�k���&�vͮ\D��+�0�`�c�J�������ֻu!��K�
�=�%bx Sҽ�7~R*�С�E-�b+0�D+u��^Ẉy�⑚����<�哚��Լ���y���=�P^�2�Me����z[�܂�[Z�u�>����������hI� Ɨ�W�9B#��=v��?���2�/hO�m|���&��R%�-?��Tǔmn����+Y�f��S���u��7z�4�{�Gm�{���;myz͜�3K?�D�vc�h����Go�nv75*� ��F[q�N�(��BZ(q[���ŕᣔ1�g4ZJ�� Ғ[��t	�ُi� k�[�%��<���mv7wr��O_}5�d��:��r��ٻ�U3k�1W��b��ŚK���R��(bE�t-����fy����ݳUm�aqs[�������!�̎]A�1��z��Dg��U�Y�ve^`���5�5�p�S��Ч���ݪpBol4�57��6���=>U���a����-���2o�6�Jt�����Ɔ���`��o�f*^<�d�]A���V��:5�	Is�(J�j�����{���|@X����
��j���tOkd�TI���F�H��Y*���1n�魑�S�S꘧4�������i�Ek�(^ =Fh����St^���ҏx�H:�V�|�;
��w�v�mJ�Y��-^0���e�Er<��$�L%������新Ɩ�<�F���L�Yn�P��M�#�E���NS�c)u����K��ߘ1�н���جJk
�'Xb+Pn�-��
T�`��a�JB���ڰ�ܷB�m(WC��
MVG��Q�XB��nR�?�����Efͼ�$[Q��U|��*�X��:Ty�\�i�U����$����.Wp�cY@�ŋO����WPr�`u�
�+�ñ�m�:��D�~�W��cUYTV�'V�籪:�����sS�	���U�+�v�4��c\-s�_�9κ�0]Ƭ�U�a^*��H�e{�|��Tq��4&(����x��!�Au�Kl�չ������Lg��1��~�9�+���c�)�5����
�?J��0�&�:4ؗ�uK�CPdZc�,��/����xF)5����˝*�;*F�9R��� i�m���Ύ�uHR�N:2R����߷�)��q�ˀ�~_:2є�CƦ�J=��C6�zQ�,�O
�.SiL�-yY��{�&��I`1~钣������"���Z�6R_dv��͵�a(�ƶنݐ�����ER��)��'���M�0��/���&{�M������۴C���"� [v���i�j+�*�[(� oq�خIӃ��_�:�*�o�f̳/���T��+���Ԍ������|�M��P�ʢ2�e	[^��8�2,@���au<�VS���iٮ\kf�hp΀����� �H�՚�L�Y�5Jg�]{�Y�˔+/X�16�hs�����̅1J�r�(9��&Y
��p���̪��E�sx��D��a�*('��cu<E��ܖJ[�6�`i�2��"[[Ƈ(W��M�a粇�G-�ʚ�r��O$K���+�<�ĊkX+��'-Zϔ ύb�1�ʠ�Y`e?�#��	�F�d�($$��I��6"/J�&:iE��9v����u�6�j� ݔ��^�]�l�ȋј���{�A[�=YuO��Q�[�x,'��]vkx�����Q�S������y:�M�-��S�:���8֭�R����ٵD��z�e�������
�p�V�\/��Q<E?�=�<(�<�׏H����� 1V�.�r��G��A���cm��iq���R��YbPjS�x9X������x�>^3g30��D���ZO��h�t�7���0}�.�ڣ�����J��53e��o�D��4�h�c�#��Ɗ��!ܖr1CX������M%��_TU6�۫�TşU��Qi��Dej������Ma��l�Saq��e�ԡ;w�p�SG�Ql�[�ab��"��}�7:���:�=x[{��,�ňK��we�y"w/��ԭ��jZcy�NV%pnd�=e�2���^��>���RLd[]y���C����T�y�Ao̯�.���q��%>�w���a��j��eT͋��DQQ�Φ]�Z2��b�/�}ܨ�^a7�-�F���Q�w4�>¨�t�K?����W�]:;ob��y���{S�T�ͥ߿lw�,�����}�E��2�!%�M'����m:/��&.�{Eό0:]NL�� ��G��w5��YS�>�O꺬p�)χ��R�e��FK��ݡ���R��նO�.�vV6̇�V�s��ܢ����ĈX�>�︤�Z��,"�'��KT�N�1Th�6�>��'6�L���P���o���<�t^+)�H?��"K���maJk�q�EU���Y��%5�;��$�ƜS㲂�fEa m&׷�R_߿x����lwl���Q�^E�kz)kǐ�*�4Ό�Ć�W��V�������ݲ�
9D�GV���7��f���6�頍�����=��KO�Ii�=��b{��%/Г6\(ԓ�^x���慢{ұ8����B�=���ړ�]x����ҋ�$���=�5)�')��f�b�X?cs8D�K5�������2�#a~f�]���$]������q�c�̱>q,b�bq�u��}@rc�ɦ��l�t�1�;]^�q��H�����C_��-�����'����ܷ�R�>�ܷk.*�̏pù�C�����ް�����߰�؍@�5��,w�Y��Y$��s�۸�.4n��w�Db/K����ۻ��_C��~��8:\B[�qh!���yp�IG����G$�?*��x�*��P^�@Ğy@�?c�*'@�4 1P ����Y�(�a�34������3�G�o�=�-����q:�W�|���Kt���Kfŉ*���݆J��Dl��]�>�t^-��(��M��s���:�QAg�|��5ʗb��i�b횺�5�֗��"4�R�.�Ŋ]�5�_�*ba}�t�#ٚ(���F�ņ�P�*N"���xtk:4z�h�8����Q� ew���P��_*�\N)y+����r!���:Dsΰ;���L$�v�V2x�:Nיo�1�Sl�r�����_��Ze�2��]ć����r}~o���N�0��>�/��N������d����>�c��S8��t!��$k�/��2z�K��iI.f����<c#%�)@��GW��Au��)���4G�\����y=�!��9%�)t���	�ۃo�O'�:�DK�]�s��7Jl�c���F�������U~��a�Z��҅Go��)�r>�}Qc�������.�X��;>D��?AR�&èhLG�%�r��m<¥]݆�W�N�m}��G�^#����Kc�̓4ٍ���9^3��'��G<��	Q����z�&)	Lp0f1�J����t$�u(�򛢱� d�Y�"D��͋Zq^��M�-�v�*g�A��SR����YN���2t�����a���b��qxU�<io:@����a(Ǹ�M��| �7<>Pcv��Rϋ�y#��r�=y��o�1G�6�ry�Ci=���q��+�:�M�ŦB�MM8��۟��1�\щ�h�a(l�{�]�R�%�v�J:�P�ܦ��$�K�V6m�ݢ�m�78Ȗ�s��.bo��og��0�E\�7\�o�����f��Fz�Ԏ1�q�L�yլ|�!\����auRr]��Sr]�/�
�9����g���BEL������V�3+>?�˵D�Ť�WG	:���=�$�}�/;���o��~�}��ۭ8�^��)����V����N�>�� ��R/�/�dC���%\)	~*^�n�N%-k����O�n"��ɯAh�$��S��Ks9���n�s"ۻ�wP�&���"��~yd/����Gk���h��ܻ�y�z���k�lqSYkm�X���6���V��P'Z���0-��Nف<c�'����i��' ��J-�=���13�Yq��<t�8x)�#$�\!犻N���h��p��	�u��Ļ,G�$����Z�)�B,a�+��Q�f,�p��|����.J�8l-/Ǿ����Λ)��aN�&�rm7ԭ�%@��D��5�gb����)n�t,x�x�q�O���l�b(V��J��-J-y�ŗ;��t˚��_���-��S�ވC�#��QqN�Kb�;�}������"�Ǳ>h׊��Dw�fť���`�e:o�g��A��Qs�Ovyp����0���i*'��A��my�1�{0�|�])��՝��:�u�P]��'��d*����-��Í �����ԡ�gP����\���a��b��1�5�+��N��l֌u�R5���g�=ċ��%�]��S���<���9��kN�8�����#~w�����},������>�q�ǥ���>�>Ⰿ]���������QN=4�X�w]MhW1��!x-͸Źՠ���,xP��n�5���o��/~�3�����g��<A`���O����l�Q��Y���M򳟋�Rpy�_��xCo���9+�ӀZ>.��Y�z~$���k.k��1�C�]������,o{͞h��o�$~�9�Ytj�D���ݠ�����"��6ԲW�lV�~�p�Doi���N��5�������j+�,��H��X��X��ް��}=�,�0g�s
,g�����ӊZS'��7�N7V�h�|��b�a�*g���R��敺x����~�\����M�dx�C9i�m�M���/�0	,�ew�I�'^��;��(�������A>�A6�^��~�EO�������*���6�O.��]�ᓵ؊*spv�v�sEMJm�u������]��`��u(D��)��Qb��ћ1�'�+�4*cx���ﮢ����,^s��Ӕ�0�����E�fG"$�.)�槕�_���4���UVw?`wo5�Q�A�F�&pVδ�ڣ�T��a��	s^z�u�� x;w�N�+΂m�$� O�y��SS��cD��܋�����7^��j�w����@�gm���q�#?
'�1�b��������;{�P⊀��h^ f�-_ ֚���+��K8yѦN�eb$gFXщ�K�f�wlkkX�9,Ԍ���؞�X�9��9��9v�9v�96�9�k��b*�m^��4/,~Ƌ��pP�u���_m�4��14��� ����}�j�w���=O!X}C�(� -C9�-#���^"B�W�8��.��6=�p��q6��K�Nځa��\XgP�uPId�m�����7VI�u7� NLޖX֍��=0�RrK��c���<O1#���&��Tߡ۬�fe��o�gq�aS�s�u=���x���t���V.�\�)��AVy��'�(VŃr�)4^��x|k�?�|��+Ӫ�]�i�|oW�&��O�U*�� ��������l>�"�k�E�A�R�L,q�醦��@���a1�ɹ��R0�Д)u��R�ݳ*�`O`B��MW��$�y�g��a_��e�gK�7��uy��������L�s]ueN�Rn�ZE�m�;̊���3��W�)�:5���Of��\,��$��(�_�-?$	���`�\q <��SˍΖ�k���ycg��5�M�`'���\=�O/��)o�k��H$�������,v`[Wz���r,69�A�re�jqK	�y�K4^�h����-�[�)�:W�)��ԭ�b���T7a';Ir���\��ex�q�O�ge��X��i��+_�-5U�y�&����cb���r�e�#�:]&"���`�1�:�VXwL���E�a���X�͠��F��cI���E��aL{˴�6�L~��쁍�xn2j��<�8�����K�q
A]�%��o�$�'f�U���4��4[����6��l+������V��}:ԾO�b�,7��DP�E\X������QU��g�!��8�Q�F	1:��JB|��`��^�;��E��e�I(��C��W�+Z[��Z@�����P��B��h�0i!J�|k�}��s�h�����>{o83��:{����k��W��k��dK�m��;O]�x�'��1w��l��+�����*[�m�j),R�ڰho{�`z��������p����"@CI�A�ӧi�ޡ�W���X�WiH>Ίa�K<Ag���T��F<Y:�n�ݶ�ߌ���JMU7-��:���K�8�+��`�[q�(�n�;Dg���U��3D�UO��"� ����)��4k��V�x�6�� ��S�!�r��5e�P]hSV�g��o"C�:���v� ͸�ְ���_��
O����"#��؅Qm�Ĳ��|��b��
:n5��&LgR��v4o������L9�'��7�3q���C�L\�T�>�CM����G�����:hI��ͭڛ�G�V��$�kc?!)�}���<��,?c�E�H���s��Xش�ܒ�+e�q�w1����ȍ\�F�iL�>�d�h���d�N�:�t� �uI_��P�~�n�� u��9��:���W-���*5R ���4z4�烙��c4<��q����v�dv�N��v�tT�j�B_k:�#��j�h�j�jYcqf�`����p�P��b���.)����c�,�-+�b޴��b�A��X��Cn�����aȕ{��ɪ`#�DM��}�ƣj�S�u��{��׾�y�$���"�o�(�1�A�T�nM�n��f�J�͚
2ʈ�|Vg8������E�'Gr��"�NC���m8"4KsT�a.�0��=�g���+��~�xo�`�b��u�
ګ
)��������j���MD�O3k�5|}��+���%�#,s?
���8�w�O�me�#�Ҭ#i.�BN��LV�oEӲ9"�%�@J������+���w3��C1'̝M���8��/�	;�GR�*:�^�E�W�������U�z��*L���{��4.L*T��tt�S,VQ��҅��><F�]�T��J�z��g\��x7ΘY)f۪i��[��5��%�JD�t��s$�d�k5`@���&W�t���l�+4~(0~p>쭍5�fR�Zm�b�T�W�Y�;��Z�jt:<�q�����t��)#k�0riYR�c���R����� ����_d�����r���0v�o�
��o�������9�a��4��t��O��t%�
VTX�>�b�����4Dޛc��i@oA�,q�fĞ9fC�G7i�ͧҟҊo�Ux��V��J!�����d湄��<����p����@6��n�[Bj��W�C��N�$�2�����ڎ���X�+㗤J�!��ۓ��t�։�j�7nT����`� hvQ?{?9}	�Y\�v3���sP S.q���L�@N�^�f��J�ʯ�\Vӓ_'�0+_�qD[��w��e�SOK�����A�Q�[�ݺ����7���g������k�m#6�W�п�v�C_/�;�&]�. ��i �J$��|,��A��]쪽KY���.M��|�>�y%�W��6�}1}���N��9\{���Ҁ U�P�-Wt �4��)���t����U$��:�a�����e*�K i���E���Gtf,��+k(߆�Ve]Z�i���6�3:8?4��B�<��,�G�)��Mlr"���M���;��(n睢�v���Ct��>~�u������k��	�;���^��b!w�]�D
���B�����F}�(+20��2"D����*ƶR�E��;��w��%���$e���O6��,��1�m}'�|��z����FL����*m�ipL�H��h�FJ6�<�6e���q
sQX�����EֻVLNaH9`;(G��4�#X��;�5��}����o�s<Z�&Se�@�ۉ��XgY~���̀-#�����6<Y �r&������R�]��9%Z�'��,�O}m�����M^���q��.T�(�� <f��q�b<H��_� �2�0�m��7ȉ����7O���1�l�f٘DD}��_���L����7(�+�ҺF�2�,��w�J��$!�٧�pr`eO��A	x�Ո$ �zۇ����x���	PM,P��Fq(֯�S��v�,��K�B#�0m�����j���go�&t�y;2̕re�����$���rA�����i��i��g|�����Pz�v|��)�FWd@5Y�t6�O��kz�Y���OY�+��U~��|��.�bc�+<� �9�|�@.��Ė�`��D"�瞅u����q8�58��u"�-׸&��c�(��5K��
&��3�E oO���s���{0GV7l��Ψ3���ktV���ji�a�"ďa՛��nЊ��*�PB��=��T��1�(����Ł�H���Z��\��:$VvK�Ƒ�1R�S�����b��h�����gjY_m��2��͎�ݸ�ݿ��m���0���T��7�c-�����r�KB^w�JRV\Z�1�s7v�����v��൰Oy�ӛ�XO���67���D�H�6�;����5O�����0�i�����\���bȉ�*oisK�C�B7��m�^b�)oKd>B�R�wR?�`3�|�FLڈ%Zf�2]�-�@�Cmi���B�P�c�f+���bs7����W�Y�7XYƯ'�+�����5��k���55M�c���:�\�1�!:��2��;O�ح*��6L�ڀ�j����Q�[AE8��zD�YP/uޫlN�9�AW ����O�ǚ��#=�ఄ~�_�+���4C!���<q��m+���6�.RM�ѓH)�lH�2�*��0ޔ��=����yo�7�`�_[S��3�l��sd�H݄3��a��>5^�i�ڟU��^��p	�6iӰ_�{je'�����k7�B8�U޵��&���%F���/u ��K�B�..��2�(���*
%'jf8��F	�L��wks=u[4�a);$P�UiwHP7!u�M��3��aS�iã��	�D�Rя�o��m,Y/_=�L�����[Fc0Ө�{����D��K�>��§���|(\����@҃D�`�l$�J�lE�M�)�{˺���H�?�}T�₤��8��X�%l�ܝ���}N��*1 �xH�zU5g`f5 �Z�`MK��s��]a��՞�l��Ve�?�"�����Pl,U�Ŋo+���Fq"���p��ۊ�Z����֛���H�0ù�x��e�3�b5��A[e���%0�����Z��[vV��	$GZ�g�P���|����׫���)�m���a���
��T�����nI��Fw��C��?(hf�oH��=#��O�#���S�_�ѿ)�KSA5-5��-t@[�����$�Z��rW�BW�c�͏<s�;Z.�M�gu�څfn��#є�A:����B$�y8�[/'^�D6y⑗�G��p�
�[O@3#�Ж��^�����^���&�x��	X�EK�+zؿ�x�3�]<	L?�WԼf�z�l�vw�V�~�����У���l4	��oF^z	�t2����f�C���C��N܅!��#�`��hȯ6�����m oOs,Q��*��>�U�w�ՏV����^��;�^�3u�ߐ�����^Ms#��+��ع��<�˷��5=�9Ө�%�O�e������G�I\�2?��Ga�W��x03����D�}J��?`6?s��h	�?��ӣ<���e��j�')_���4�SF��,O~U�e�/a�y�Z�N��jQ�4ʨ�_��tJ�F�=2i��:��� W�% ���%��j4*Ǡ/>]ǌ�*9.A���H�b=v���<iO�	WPn���PF R�@��?NioHPZ4GSs vJ��`^� ��+���XN�O)N��ǲ+/�X��Xn4��Zm,��1�Cv�$�d恘c>�Q|p��U��U�V��U�˴���.�7�n��8vR:��s�4'��Y��6eza�\��rCɥ��u,�.M�0�C�Uf�Kd���Z��0�~��1KoӲ��&�*���݋���\.,R��nbPx�x~�/�a_���Vzz��Z3�Q���ÍHTB㼔����� ���f�h�����%ZҞ�hcq�cM�ԩ|5�e� q�"�A��B$���,Og*�[ O��њX+]�\��a�~wx�<� Q�p}�9ה��"ƃAL�>h� �W`r��B�Ы�f���)(����Ѻb!�I�IV�b�P�Q�0]H}3�|�VU <�̿Tc~�1^OxGSȕ�#�.o�)���& �ƸQ ��Wץ����BeZ��_K��k����{��dl�T��D�X�������p�c��P�A�]JU���Ӧi��Ch/��pKToP�ER's3���º��k�K��2�ah9�Z��gM��"�����+�,~em�&%
�	ܮ�;��I6$ٮm����n��0'p�XUD�����Hk[�_mN�O��Ȣ��ͫy���Gg���!ҙ�C���1�&:�c�A�,�k&ۊd��6�h�S#�����v}��i��Go᧨zi�u��po��ः]�r�jj�{��D��j����z�9��k2��PK���
VJJ���M�A�9�S�pu≮ʍ�>����UB���#p����(�at��0�ʵ>撸��j,�e�}��+�r�6=9Q�z=��k>C~�����k1?t}"?�e8�;O�I��a�~_��s��WK=[�K��[Os��.��,�H�)��O�sJ��-���/�GF��'�.R�z�qJϳIN��L���y�J�_b�+2E�[�?	�)U٥I6�� �睢�J�+�#���[����4��/M���K�p7d����7�S�QϓHǨ������[×����I�2��1h��z�x�q�T3�ǣN�gIt�irjPzj:����;y�'NΔ7~�Ӊ�t�Ϝ##ݑ�X����V�x������_?�kB��"�5vps��B�N�*�*��Bs�ċ�a8�UO1��r����i�`�v��0�l��S�Ј/%�'�_r&���6lPљ��n��\O��+Nk����E:�|Eu��<��$��Y�tp��� �(}�}����߉}�AgV%���C��>�9�y�F�/�}�E�s�K+@�<{�7��t$�:�6�>ã��fX�l��<���u ��ޣ���F��~����F���V�*B���
e�V�H��JQy�oL7��£O2rw���s�æP�49
4��9
�J稥�R����[/2̱��%t)�)[��ŀ0��m5�nr�+:/�9�ճW$/Ǩ�rX������ǨɊ���	��"��՟�^�/7hVÎݶJ���-ǲ+�q�O��t�`	����I�W��{����o{/�y[K�7�@_�te3�/#~SP] �^��'��@e�Z�ɬ�,е�|V
����_�n[R��LgW�YE��@,$Lۖ�u��N�U���9ԼH����vX����z�~�~# �xӞU�:�VQ1)�4��ɭ�~{)`�r�I��(K�F��Hs���I�7$}~%������>�x�P�?���5B�-[^�A��0rl=kzl~X�>��>�ه��A�t���wX"�7����
JO�x�*�������{+��p�N��D��=��1|(��`ܘ�2�Z��H+i��:���K,u����Y�	�����0���TN�����@��d��*��%T��X��ާ�V�A63��ԇ��e�+��osѪS`��W�m��Z�\oue�V�w����OY+� X;���n
{��$��V����_���?վޫ�<�̹�Þe�^&=B��m��tn���n^;aZ�{�y�-������{��=�����>�| 6p٪�B��Wl���NB�S0�.��my{�(��3���E�]���6q
P�aåˮ;EU�eМӀ<���->�:,���W�/E�>�����M���k�V���J��i܏��\_�?��tJ��#?��E�)V��$/�3l-?^$�~��{�7N���S8�)�l�[ī���mᛪ�EՑ	)]���^�،x�C�֝R�ɾ*���й��u��4�^7!+�7h��m�H�q1�����T�Hr�����b�%��)�j���ԧ
?�%Z�{��23q�:� I�+�TSP m=�4[����I���4���|�#@WQ�d��rh(�ݫ��c�@�?�0]�j�5 6��b�<�q��Y-˦���KSn�e�"Ow���A��K�❽ñ�j�c�2��Kuxluu�S.�}��i�8s4���Kyi5
QWO,$}\�>�����use�T�/�K�޺t�֥
��h�҈�pq�.]Ĩ������+;O�WW���+7k]�N])��Oەu>\/�n�Oۍɓ���hPH����JUO��k����M� �'�㿊��>3��>��'�-9n�I�����x��ҷɷ=���3`Fs�r�:�Y!+CI�̥X���~�O��SS;�iI�n��������UPA_���2�/W=����ʫ�x�}�m%�P�	���*7S���Y�-2�=ހ�v)}uS��m��r�*��{��Zڞ�@���/B��1'�Tآ��S:�z�g1;ҷ}��Fu�_W-��=I� J��
��y�U�Tǃ����؟��=���*�EU1-����v�6\��	w�z�M�.�ry����a5��l�e{�ʪ�"%�U~6���H]P~4����\�1�^ٰ����݋a:[án������8��7��=�d�cNuJt�X��uu��U���]���ۮY
���V�d��F� ;�h29��W���j�+�G�߭�[Q|
r���[��8�D�`�`?!�R�D�����<�b�����^H����}���f�.����C͝�T���n�I�\d�3P��c7:�v���P:�������gF�SD�sX��Yd�`����Q�r�B�j.r�p��Uᓫ�z�7��x����!|�㳈�	~�Rn��(�Z�n6����p�'"�ȸ���n��@DoC�%�~�@M��ɑеiW��'�ޠ�(���t�A�ާN�]�}�T�[����q��X=�l�(Z��?�+@�+�>`��x~m��7T�tF���O������k/�D��(N���Ll�(T����;@B�)��ԯ��&�ȍ��@+�ˀ(	���)��ֺhiN8�l������n/�c��&�UZ5�Y$#�����I������p�13�աS�����g�3�<�P�=lx^�2�t����a!�rC���Cz�H�J��y���;��Lϲ(?�G����	���LC>$�)r�*��M6;�`��p��c2^#� cAFl{%z�a��1XkO���	�Q����,�{U&@͎Θ�8���ep@��s
�d�Ej���hu!�ڃg3޻Φ��Fw��T�@ʃN��=ï�D�L�E)��z�|�y!Dr�s?~����h���U����7��f�C��̭�j�Tx!2SR��hG�8b�G��Fbe���I�Š��qhNl((�v4]�����Mè��+�%�U���ln�Jwni�Nx�gp(G�O���0O�S-ou���	�x�!�h �z��P�N��w����Ɨm820\�_���wQu�?Fz���#*��+{v�쉯؂��b˅���Ģ����FtR+؂�<0H�8P����.���%�{�84-pG�-o[4 �mY&�n��|��:r��؂���v�&h�g��a���s��� ˣ�h��zR�����	3���|�Rξ,��;ب�.VY�*ܿ8������N���U�h��1�K�����*�MZ&��}h¯"�}�!�?x�]��Ӆf��ȅe�z�Ĩ�|/2ɬ�x�T�-:��2<jܓ��<�4ڠE�`ؖ_��;�$W���Q6��,7.�ƫ��K�����?Q��&��vt��gi�s�}��R�1[��j���E���r�LuKc}(�%@�˴ׅ�E��	�b3<�>�յ�4/��o#�v����A�#}��$�5+���Ѿ�44-ߋ��q�\����-�O�u��=��`k*p��e�1�)O��c)!��b	à 8�������!�ô9�Ɔi��y��u�bT[a͇,#��`oVM+R�֘�J[r�!�M�c�[�C����r%h(�l�������74�����=� �`1�F+�4�/��&�I1�]��xDi�R�G���+gY6��)���e ׫η���Q��0���سgY�5��<�R�!4���:�\�����t%m�Q��7^��+��Z��4���ڗ�X���`s��+h/�2�v[�u}A�;�ьu�`�B%��iy}��,ˋ-𬼤թ4}�s��a{�4�qg��Q�د�m� .eT�v%g
��������t4y�7�C߃O�v/��C��_��l���]D�*�]-�ka��F��<�@������AK�)��S�I��,
R�(�ɟ��1H��P�$�G��Gm��)t`"ߎ�k(b*��Pp��|�D��C����13���Rv�6���!�R
 �'�e�Km,Pc��8�";S�u�bc^��S�ш�)?���(���泊Or��������U�����!�R��KΩm��iY�`�Eq�U:�9�8Ms��x��ƃ[�i�X�a7��/���� V�D!y�2��̸���s�����HU6���y�&��j��CZh�*�'U��l䯰�f��/zZ��0�z�&�=!W��h�y���C��� ��Ó��|�"[�QwE�����n��!�Ċ?�g�3�{�;�,�5}�WyO���\��F/o-}�?h�WZ�����E�zճ��ǚn��� �yN�K�W�����D���Np�C�{��1L򣏞��]5U����N�S�{4��-E�R�5$;��Q�Ev�S���޼��K��=�$n�O?����[QB6D+a�;�^ n:LM��ߣ�W������x��mu0���{�� ��A��e��L�Ce��v)-���lxi�,��L*����VY�`�Ŗ���O$g	^���R!�4Kh��(�=����dHNh5ۣn�z�*S���%�>�F�z	�Aځ�����8�M�����"R�����币2��?�2�0��0�0c6f�2�?	�=>ax��Ga �D?����nd�q��K
�Y��C���3�d�D[9��������?3*v&�����뛤����O?�E|e\_�pKN���ii�ǣ���e��/J^^���-��������9����V/�__^��(�]hX^ׇ�&�'��2S�/�vA�������%{��;�-��6�|n��p��b}�M�řE.)K��U
٥)6�7��D���'�����l��g�ow�v�&-Lsl�)�e�fxsW��Fn��i�;�|j���B>���Ě�n�;=v��I Q��<��h�c�	�Uk{
��a�1'~m��~��$��F96���'��:�į�>�1�	��y�K9�Vσv����,��Y��c��[qD�͢0��ȱ��ه���m���ه�ֿ�����#��c�f��w�N����-oo�W�G���O��?[���k�1�~Jcd��h��-�[���ǎ�O0�μ��u�3���^�������w%W���j �7������Yj��j��t�,*��G��m6�~�	8Cΐ�3�gW�=7��s��G�2�"�NZ�����?�:��\߅:���	Su����S��UkJ���gyj������	��2�ޘj�j�?�'���?^�3���3����v�����6d�1�>'�c�1f���gG�������[�1F�c����3��?�Qs���������g����=�) �q�؁=���-M(*��6���� ���D�J���$����R�t�8M��%��s�f$[�a��J ��,ǁ|�����!yUh�h��|&���c_����htB{w���wm�����n`@'p�KDƝ
�&:�V "G*N���T�F|9�*ymR�.	Fy���4~�����y.*B-�'�Q1R�]����)Nr"�Έ�.�[�A��[�� �S���	������{���`�*h�(����Nx��k��B=&�����IS���;0��6'�� �@׋�ku�-�"ǥES-��w�d�C��n���:i�ճ����[ZR��FJKJ<;���-�����K����T)H����5�.58���ؐ��ٺ�O�Y��=�얷���Ǿ���t�s\����}�tf���N���N�qyM>�.)�{�C��N �^���>O��>yU���t��)��D������{:嵗���O=_�I'~���<_�%7�������'��=�e����u�ǳ�zbC�4��n�]��Ny� �����9)C���8����'�U����e�1�8�
���;���������	�i)��ǳ`�AO�M}>���H>`�s�od��+9'�F�J��s�ol���8'�&�J��s��d��=ǈ~vg�����л�z�z�xbԻ;�?������W�ݗ�8�����лp�t���=;�Q�g���h.�	t�_�n1ϗD���w@��Es�W�k�^��W�^{5��^��W�^{���^��ҫ�ExU�K�6��W/}�X�d���"��륇����N�9W'�9W'ך;)�j͋A�!�`�n,B�-x89�����[�����[y��a�m,B;,��!'��K�vB;��Vo�����"t���|zH��Vj���h$�J�����"t̂%sb���m��}h���j�;����"t��^r�5��v�a`�X�YX�6��0���0���0Z�s��0v��0���0���0>:�a<�a>�a9�a=�a(�9��È�.�N��?n����K��-aj�v	w�%L�.����A�%�^����AZ9CF��:�E|z��r�NR}��:�:W'���d��:Yx�N��������su��\�}�N�����3������FR{�����4
T���W<h��A;h(:��s�Z�8�&��b�s֌ٵ�bk:z���1�Zӡ�u�E�x1"8��)�D�z#�(�A9�9Ѻ;~�X�	��`�"U�5�S��tz���̂"6jc�剄�W]Gm@�r�s�u_��S;,M����Cm@�r����~�qR'� �#7�PШ���nݕ?D\���k�����k��MA�}.�6���������bjS�k�GR������ڔ�����ft�}.�6���y,��[�G�zk�|��h�Wv T� �5W�N��G���Q�QB�������j`H�W'����GO�<j�e� ���X��������%j���g2��� F��
�.R��b�!Ã��K�����X(��40/�.�ע~D��y�!=���.��8)�o�4���>Ƒ%����WJ�Ҁ�sr�^W�:���_�4���>�Q%HQ�Ӯ��NՀ�pR���(�)7��N׀��F�b�n��w��#u��E�h@�z#D�N7/������u�M��A(�!Ju�M���4�Žb�N���w�T�!*t�͡�ab��h1A'�\��X��sMo�֩���wz��]:���`�4P<�F�N��ڔ �#Roԙ�3L�+�k�A��:I��3��L����xt�9�4G#,'<�I@�3P
uS�(ұ<PV����5W'r��L�z����x(�C#\P��J�cm�+��(�J(�C��<��8�u	D$@DPο�Eph�����q�c}��j�&(���@�M��D��8^I��x^4]l��g�Æ�-�E�z㤬��'�l=�j��05������󠯶���?lI`z�<��	 �4���&0�<Zk��0Y�CKӞ� �&��:x/�i�yQ|ô�Lhxؙ���yQ��i����'���yQ|-ô�Lhx؟�t��(��az�Lhx�(���yQ|=ô�Lhx8��t��(�
������p8�I9/�o`�6�	G�:΋�3L[̄���	L���9ʹ�i��0Y�%���@k�a��4ac�����#���@e�a��4Ic�����3���@_�a��4c��#��+�����ô�i��0)G�Cw�0z��N�c����Г��V��h�����LJx�h8��M�3ͤ�k�Jz��G�a3)�����:M2G̤�{��4=�p5��	���C1�\	���Q���LJxp'p���
��i&%<$p���G����P��1�4�d8�ͤ�����sд��Ч��qk8z#f7�4����*�0`��x�P{!߿i�b>���oL\�h"e��*+e�����q������U��يŷ��TlZ"�������	9xW�NLd@�.�
�\�:���ܵ�W�W�jRu��1�	۟+o��$��6�,���x����3W@j�k���0�k�%f}���B�,��Ȝ���2U����fT�N>��t-���Vv�Q�C�=��}�_!�ݱ�E��VF.������U��i�#��5=�bZ��\@�����C������D�e�{ؗȏ<-��r�U�Q�}'f>R���tljI��Ux���d��Y'�n�����l"Cv,d�a��Y1'8��,Dn��l���أ-N����$��"�G{>(�����րt���*��5�j/��tΖ&YE�Xe�r��,�SaMQ$-G�8�A����I��=K=�&�-�7B�  -'��6 �����E�~�bv�B��+�1���*!WFP���ar�J�٤�.V[�sl�м+�Go��+������<9�gu�%3�y5	���&h� ��jE�Gx-I8�މ?|��)�w�
H��M4hq��pN�^����ȭ��p!Cd�R��&�ʳ��|k�*^ϑ�6q�U�?)���*.������7� #}�Io"ָ�R`���VW�!-�6���0-Υ�#~��% �<���@o�~L�~�<�i��k_��0�|��O�/�(�QY��)̛b�aN>��
�D���Xz��� �q�/�VcraL���`L�-U����"eu.J^��hs�ň- 7:��mG�f�E�-�R��U&?�R�þ�����L22g�a��ݰ*j.��YT'���-ʆ�NN�������O�F�-�R��e���iI˴\J����z����^�ĳ\��P���_���U|y��P=р���UZ*�ֈ�9>*��O��o5ƁY o�
!��D�3�*0r�ĖYs�G�(����������
�hKz�^�vx-��D;V�)�`��Q��X��O+Ø���{��ȑP�'���;na�W#�z�1!# �G���[a��B����Sr�*8<�P�l�7��B��`ý�f��:o7�����	�:�R���:���gՕߊ%�[YI�sI�r��-Vs֕@��`��Jĭ ��e�brĚ��s��g�H �x��ߜ&9e��E_�n��si�r1��)X��� �G�b
��K���~ ��_W��SUuG�tM��SkØM�ψ�EG[t���R7B���O��@:5< Z��*/`b�l ���q\:�ٸ=j��e������H#g�8`���n����'�������ۿ��e�S<��ˌY�c��5���B�H%b�4w�8-���&����tx0�R5�2�瞃}yB�W���\���C�0^<K���������t��	�:=V�kNI��T^K��4��\����.>��i��lE��*%�4�NDۆ!����7����A�-�����JgHPJI�IJE�Q����4ъ�)Ć.P����r����hR��,��Ѵ�쎦w1��-}�v�!/�D����O��9Yڧl:�.��3��N}��1���9�iη��v!�J'���HN�;Vqj^��u������T�'�[O��TQ Nț���
�Χ�`� � �h��g��	�+�S7x`ѺF��b�C��J���K�ܙ���ͮ���	B=�'��������:�;ڭ�B��ex���nJz�;��B�����귅�>y)_�F'u��^4�^��&Pû��S�D�T�"ޕ]LO��X�� �SA_��jz:O�+�Q��Wv�h�M� =eB����l��+�g[�B��ɗ���D+���}�W9��9L�hia��;�é3Ǖ�q��,׀b5GQbD�\C~�΋���u���
ңV5������#�F���F)
J35��l
d]F��/����!Z
t�)$�>'Mt��]&�iO}^Q^CYU��_�̀<׌�|�[���g��:�9y�
���?��O�e<(݄�RT~F|�qJغROغ�r�~l����M�yo[����Lv�U銚����h��'2��r�,���5�K�:B�X�i�W�	�}֮��&mBͧ��[#' ��H�Iu�MD	gE�)��U,A<6�}w�]��f�~#/v�gգ�o�S*[ln���Yb���^�fh�����"�۳��(��1g+MbS�m2`U��
�y`�1��i���¸V'��&�磟)T�ǫ������P}�F�l���M�Y�_O�� �=L�MB5?C���?I$�G�����؄!7�D�ʋ�E!�ݺ+�۵��y��kmh��[8l�w�L�G��(�NQg�A�m�밋S�����7��I�{��� Zw`!0�e�.�M}����O��TM}+��Է;��4XƧMꖛW%z��v�2�h%��Dtf��X��l1�Ԝ�	��w3�:�T�����N��q��k��_��d�U��m���L��s*�p�ڎ
VM~iE|������,��>Mf8y��`��vf�|M|��t�bl�ĥp��}y����6�0���v
k�S����nV?�<�p!�]`�� ܢ�0��om-�휓���wVїͤ_ڥ�����G����#�K�a~L�»���Q�ԃ��f��V?�6:���x���)��߫����Pq�O������%
/����;���
age���Kz����s�?������W��:X08�7(�2����a!�]�4��4ʊ�#��H$�C�}-���A��+N�)�#�{�5��U��E��D�Cc�:L��Ȧ��:Mm/4 8L>6 '�vƈ�+Pq0F��, ���C]�m`r�I�W����MXzf��W|���?�u�X_�'�D�W߉k=|ۀMx���-Y<$0?��0�Om�$"��r�����s*v�y�k)�Lk��=���
Η���B�u�}d;â�A*a��^�6���5V�hZN,��ٖ�b���$��@|�8�G�ՙyS斔�k�
�1܅D�R�%���+���5N9�ƕR~Ҽ��X�� b&���~>�����.��C� ����!��#�&G������ �ܰ��
t������\/_�舝�u�%�Wc����8/7)?�%�n�x_�_�?�*ۂiu�n���?�ĜydE����kmf�7z�+Wvz��]�:�p-��t#�x����C�[6�	,����F5ҩ|�U����~�e��1�c��\�����Y���N�7��oٔ�����B���*����^&�Ш�N��W"�z+�3�s��ƺ��PXG�m��G����������y�����r��˜�I���"//����#�d/����>LJ�c��;F�Q�UW����܈��m�)�GFV�<L���GD��U��+U�*�>���A�_QbE@��񛋇�)wl"�/+���N�}��؛�����b��/^�_��vF���%C�/ʕ��i��|��U�]�Q�1|w(K�Tfȕ�������R��#u��\q�)5�����sEeO��杲����7M/�o�9_�׳�FFh�Z����E��u�����Ԉ���u�?�b��jhT�z6aTV��X�K�eg�oX�>��6���EL'��l�-��a덏�ZVmg��� �� z%�0 ~ ]݉��s���~i4>G]B��9U�j��ې�X>p't +����r�P�g+ם~��O
	�hk�6݀�W�>�&���]p�>R����J��6�B&�*�u"}��v3	�:ĉ��k(�V6��������@�| *��h�9��fW�g���֯�t��u	|�tZ����b�
��Q�p�A�r�X���Sj�:ϐ7g�Vs.,����K��wN�d��+�,��O����Q)[zҰ�u����~�����#�����
qK\QLEכ�(�;�H�O�P�&ծ��8�It�#���\&�ʐ�,I8��7�MS"[��1�kY��cgҌF�~G�u�א���4�@��j���%�r��h8<%V��4K�)iY�9
�F�t�����X	ǰR�J�E2�G�<�a���2%�j\u��^�f�eMr��h�o��e��^r�}���e�E�3�E���sIhR��b��%�jnazB-Oz�,S�wLbO�hB��d��6�*֤̇^��q����H���C��z3WǛ��p��jr2T�t��cC�:ɭU�f�Y�5�rc1fi�sя~����p �[��p���b�{kck�چ�s{Z��ہ<�D{�Tѝ��ǩJ����K΀R<��u���a��Ft� ύYi�U"���r(?rw�OmS��9/a|t�]y��J�������+0�Ar]�c�D��ީ���Tux���h\����@���{e���t�ix����x�A��I�Xve?DK^�;��`x��� f�x� 5ڣ��a=��fGٴ�se2� ��Te����V[�kۂr�k��k+��#��-d�1ok���]/A���`���:�.u��Q�T�5�(�"n����)߱`&�+�*7������DBo�J�u���څP�4�Y':%<�H�fIq>���F��Pqu�Rlˠ�\�JT?��v(�{zSg'<�W?���\'tJ5�t�SC��k��b�����Ul}��?�$�X&6P��"��Xl)6������R��x���z�f.���6-^r�'yX��X�q��C���H���cn♄�"���ȕ��Lg�-�o�.A�'�^�)|Q�[T+����w�Jo�(���>A�'��!���]E����L(��Q�!�:��c�(
��˄b��b2�88�����vh(���τ­��O(�:���ゎ�xJ�g�P�O������(
b��@1rJp������b%�����4��_�����n~Z+�@P��.�ߠ��7������k�_��^i.9�ӊ�@�rA� S�� Ŧ�����`D���T��h��)Km�#�8�L(���
�Kō	��B�FWj(��(�ruE�B��P�P\�Q�&���\(BQ��8\��x0�b�P,~Q�P<�Q�H�(9�BBq����Q(9:���BѲ Q�P\�Q��C�fb�2'����	�X���r���2�lOp����CY3F|Ȋ�8�6º����(�����9�G|�hBe�p��q��E� �;�$o���8/�g8�:��#��Ŝ�Kb�PP�^` ^�|�C��:���m �<�!���8�X�դ��S�d[���B�r�� �n���\�_��۝�f��-a��B42�]�v��0��[W��Vo=">R�ݖhm��[��^���k \J{ҁ,c��
c9ݫҔ���{VӮp�J[ŤH���a�twɅt�)'l���Z��M��NU���/W��X�4�Em��/ܕ�Pb�I��Z�X[ ���Eʜl��˞dq�y2aq�/Ncq�FsN'�6�K��N�x�éݗ�]7�`�b�	q �!���R��%�w.�Ny�s�0�;�O8�l�-�Ј��Jg������D�ue��"9�xr?�|��X�U: �W:٢�vxN�u*�N�C���D�NSW�G�P��4��,k�9�n�6$
�W?MJ�Xio�^��l3�7��>��u!�B�ET!�$���y]+�u���'rM{��L�p;�oeh���O�&����Ѷy�`�7t+�jsݼ �A�{@���&4�_��ƃR�k5N��O�(A�sѩn�U���D84�����O���5Zd"���i.���E�ngs��y���0��m�Ѽ�R}�V���Sr?��L^p�V��x�x9hy���j�����8VT�v���,[�,[�`���Яɩ��s
�t�=���P��b)޸����)6t���У�(�}���3����}�a���{�=K�H7���vv V����#צ��Kp�����n~M����ux��4GG�2~��]q�������g�����{A�U#�j�Cy�	r�"��d�t_1&��3��~��n��L����R�t}��\���O_)�v��v�{ ,�0��=�
ͷ���̅\���%hvb�!�����%��%$��.A	^J�-�u���f�B��L@K��y1E�&rU��U<}�k
��L���\B� &��:�p���-F���>��$Ϸ=�=��n#;����+ M	薀�.QU�Ύ�JJ���w]�Y/�v��薋����Ric��:�*�&G���v+p\GG4�R��BǓ-��t`e�X}F8�J���p5R-E2����s��CK.��N�� +*�F �p�7��Ym5@�x;��%�G�|P3�xP7.4L�r���.�:�Y����|�nkc�v,��\��,��m'2��oM� ߫�� �0V�4Y���!x)y�a��@�+G�n.���n0P��ƞ�V��d^�\��?@��q劁h܇��Ѧc���#�/���C���a���:��&����AX���~V��w:$A�ʣ��u�ԣ�}\$<;��x?�+�)�<���8��W�z�Ҟ����g!��P5�	B6��龀\[�C����a&�n䷹�>��
Y�K�Sh�Jut�3/ĉ�����M)l�˪�K"R��T!8w)�UP]��T�dЪh���w�C�aQ������O��TD$a�o�r:p�J�2M�ߓ�c��O�������x�A���6�n���������#$�)�g���Z2�m��2�ݡ���g�A�V��\��ZXw^��<&�uĺGx�~�Q�n��U��>��a X����N���4�NE��~�B��5���\.�&fM�mɫ��5.|5�]�%J�MR���%8.��I.��@�eص���Be�g�" ��'z=MtK�6�:ڧ�#��J� &R���������Ώ]�'��Ua@݌�����7�sϮ�"��$io}��2_���o���(�4�F�Ε�
)��؂V���^{P-߷��پe�̸o��q�XH����p����YR+���J���8<E/̓ZA��xx�Љo�`�ug�ک1�����,�*��&�63S���/0ei#4g�G�1�t"S���)	�o�U}9SV�p�4W��E[�t�?Y��}V����x�kd����A�yF��G�y>��l��V�/V������&x�!wD����;�}�YB�e���������Э���	�N���4Z~'5�r�Cۚ�h��a�qd�� �</�@;��D'����>'��Ȁ�nY��!L�Fw��ʅ$�R�E����$#`���G�l4��5o�E��W��՛l�����@�f�Wsjg��N�!	�Goe��S�wp�vh4NW����<�|F�����U�1�_��f�F~fb �b�\���/�7ƺ\�LG2xk_�Ct�K`�X�gm��I㬛Q�<j�-햒Gi#,�b}oL��69��������+}͜u��iw���N_"�ԁ蜎��&�T�+�j���a�}���*��q0]h{ۧR�&��[��y���0GQ��K�(���T�)i�r �O�(Uo2H����qe�x��j�!�Ta�9�`)�-�zɛ�'[N&�E�$3�ͫtq����P�Z���r<oN������}HH^ {�Dsqy�5����ţ�M΁Q1��={��x)�9@<������ �`ڇ��-\@�z�a�^{��.���^�؋3�����gG����T>3V�D��������l�� �'�����<��v՝��L=��7��_;;��D��_�^���eăoL�x�0�A��r�4����t<������m��iO�1��RS\ݏs\�/���q7��؎���L�m�i�k�a�̫,[��p���P����7��hC7���0���'��hE�R�nϙ=��?�4�!��/�mf]���_X��q�����ǰ�����,�������a�YvQj ��ُ�\��gĩ=��Y|���nK����/���p��ߏ6�\閐 ��?Z���y�*D�7&M�J�Z�=TvD�Ӏ�.=j��P��me�Kz���r#��Tn�Qw:T��9$?T��d G0�˻-��=�]�E��N�W��˾`���24W��nz)[�t Z��q���k���g9�_�ވ;lb	�v!��ۗ��P����\�E������e�HR�>C�laْ��~,��������� t�����4˲rR��F�''?�K���b�b���yZ�x�$�4��':��B�ЭbM7�ax�g������$)��R�k[B��t0�t0��!;@��B�t��g��GY9�&�!��+Zq��C�a����;M�V�c�DSGC�p>2��ή�#��2K��m3v��޲c��=t���N��^���)���Z�
c��=�P�?�N�)��&,�ˠoI@���0��0��l|��P�ъ���8A_�A�9k6{Oƭ�k�~c}8�Q��y��k ����b}���b����f��y�}�T��V�гhF]�fKd�췗O�Y�.:p,�W�8yn�-]�z,�>�1���m�{�B��y��MV�	Ǜ^�Zi+�f���>~>�ڶ0ɞ��X'��g�?�����&� �ґAi�����d�Q2��s4#̑�0G2��m� �3�:����8O�Ȍc:�]���g�|�\���? O�Q��QӀ���_�~=U��A�Z�Ub@�E8S��ou�_�"r8ݯ�۳*yR䪰Wn��O}npːV���=V��o1�w}��:6g|�T�'͏�p��l�`�;�l@��ՠ�X}�B����H@/:d�R1����Rk�����@ʖ����-oJq�7�O'����x�����"�eNz�f��ɷͩ#̏a����T�%^沗�o���!|E��~ d��h/s��'e.��6��]���[��~�çaI�KwPg0��㛳��t�%@���I���e;��oC�{P�[��^��ID��!���8�t��{�{�	��;Hf��/#�`�R�h��v�h��:� g&��U{)���d�����0�Xr���%O�,~Z�xUL��-u�@�:<���SURe���|�{���nF�k���{�/�$�ub�6�W���������:6/��V���?\�O	����)�ם����[jA�9�x4n��K٣N�^b��U��S a�6V���eǭ�7WF�N���`������w/?��p���c�z��թ\|/v<-ڀ��:��+|x蟦o>�ф9^��߿�Le2�K�Ǹ^���u�W�/t�6�}�A�"�G�BdX:_�[��{�Y�br���Q%��]A�o"^h�&,-0���nF�~9L�M���|�
n�=C�Se�Ҥ0fj�1^8i�֡�P�[ZX���~M�)L�����'ϪH��)�h4/�y9�,��њ�#�V��>7
MO'���ɉ�Y�&g��M�(M�0�ir}rL�\_]:>9���1�:�7���������6͠1Oc0����@ϱ���F�uD�6�	����C�����hk�X�Ή��q��X�i���]�r���\T.��ͨчK��	K����j��.��Ӡ�۳1��4��,��g[�yΨ��h�����>�|Q�a�]xFm�:^}��P��'�Z�����i��?�0՝ႲG�_P�U�H0l��tY����8~�/I�H|�� _p~ѻ}���������Y��uR�N�ź�
�E�z��v9���K/�Z��(T
3�cLב}���òd1�&A��1��r���uN�����~gx�����nqV'bq�����Ϙw��:s~@�9�q�nolE�wJ�1Y��p��0�.�P�x	G��si��y%�
k=au�X'�fcl�C�?S^V;/|Ay[���GS�T»�)^��ҡ����P��qJ�d�t�z��S��T�]R��$�|������W������i��#*������iB������Ҵ�軶)�3��I4M��KA�W*�c<,G��k�F�BG���O��U˵wA�o�
KN����	��S�,�"z�����n�
rX�K���$'��bb�ɓYT *�lT������Љ��p@�Ⱥ��%m�iF6�'��<�6��~u�?8'�ʂ;;�c'�5���sH:��I��z[Ym���#6t����m��3�_�&�o�~!����.X5��v;�0K���s�U��z��@�j��?3��9�:�$�]m�0@J�!7.ƨ+yR���_�U��{r��q�M�	���ӈ)I}Й�7�2�Tf�����"�}���z"rlޥ���ei�[���Z�S(�x�D<��]�G�}%i�dD,k�IǙ�'iC�&�nq4S�^1%���*UT1�Ѫ�k��-d	�A�g�:��0��}�:_hf��u��\z��ٙ̉d[A������]l�n}729pA_h��`W���m�"vaAgXH��q(�N5'W�O���������R�&'D���;�@q�>��#=b��;�o�&v��(��4v��}���ǉ͡
���HY�I�JR�0
Z�<"U:�ʣR�+�}J�t�C6��C�,Ж� (�4=k^{�5�n�4���цc|	_��ʹ;�n�#�O�$?�Ck G_ԩ���X�Q�ޣ!�Eg����k`6O55R�\��25'[K��6d(��������"V����:S��N���d��*��"u1�/�'gO�6"=<���^��b��V����җ���i��@w��B~i�[4��I}�6���\>��9�wՠ�h���r�	�O1;n�?�W����;���䟍�J~��Q����un�'��q���\�?��O��+�蟒����+1����RA,ʢ�UU�����ըZ����-�`>Oϣ�$>��]K�����������N�\-VMk+��	b�\�6(��k�׉�S��j�v�X;G�ch��������!9[�~���+�˓zP"x���(�R�G|�jb�@���Z/���S����*g�k�r�|)�s`0�����}ʯ����N��)���^ٓM��~��-^m��5=��O^�4Q�?��3�P��>y�be*=�F(#<���Ge,����G�Hje{F�*-�,�U���mF&
����)h����y��_ҝ��p�x�L�oM~��g�}�.�RX�`iNʆ'J��������XV�/O�8���;��6�{g���r�;z����ޛ�7Ue��/m(A�bՂA��K�EiI)40,�Ҕ�t#M
(E0��|DQAQQQQ�aTFY� D@d�Q�a��	�(X���{�}K�6�q~��?���M����g�瞓	߸��G �7��9�+'Ų��o�yR��;Z���l�|�zf�+jh�S�&������G�<�IbU#ZJ�Ƴ��~#����|Gpm'����ㄱ�j������Sh�/4��q���bp�Xa*�U��0��8J#�q}�H ����u�[�%�9Vƴ�DgB��/^
��߭�/P���vg��L�}����?������»����E��ĳ���k�<�WN�q�s��6�л�UZs�Y��;�������! ��z/����\�]���+��h����yɜ=�;�b8ܳ�������8�q��������[��tD3]-�I���D �Ѓ8��_ĝV�|���Sѱ��c��K���� �!=�Z�?��H�G2)x=WD���Ny{��M#���d�%4 ��1BI��xH�p:��>���#A������7D�6��Hl$�����9+C�I?(tt;yC���d��O	Cׅ����ĆG(a����� ¾�5��s�id_ׂ�9��gB�x��
����e�̐�����3t��nw������sx�<�r&����Ʀ�;�P�謃�`��@�xe���Q����H%�Y�o���JT�v��SPгXz�y�1�4NT��r���qc�HaL�ŉ�7��q�7���Xʅ"6���V���x�E���V`��^���f�lR������2�U,�Ox|1=˼X$���2�$�,|!��<�&�K+(f�l.�/�����p�ו'����_}C ӕ��ɗ_u$? G����:��=�@���QfI͙�
>;�?��8q�\��~l�A4�h�<��#'��t���6(}Q/E򌶕��<�4g���02z'W	{�z�=^$
��ć<C>^$*����z29b�3�4;��l�'@΃����lyb�����&wE�Aj���~I���M�^f-?�$��d �e��6���' ��ͳ�#L�3!<���ڸG���Ӄ�h���˞��+�[QI�QR��h�e��8-}K$��Qq�$/�5s\S���M<>8e�*z�� ��5�dvn���)Z	 ۲���'�F�MP^f@|R���Wp���#�kdLH�����}��W�*���.�g)�g�L|�dh�ڤ�=�o'�� �kۇ����
ON&hqT䘗S�w��pB����.\�D�xMrW[wϲD��a��z���	OO���A��.�ر4�z(*O��5�Y�pp�T�����~?>,hU�nP��������"�ˣ���An0��<��N�#��Dw�5���5Z���4���#	b�_���t��:���u#�'�A).�b�F�~(��o͑��8 ���e	��=#"<	F�ݳB}�z�S�2;�v����҆ͻ�3~K0�Nc�sq��¡��6�B��f>T�xUN؁�B�r|j]�#�ƍ��M�PH�d,�2Set\����D}A�G7��/�`�v�ȅ��� ��\��Sa�V5�i,�|
��f��ǹ�ҵ��7��͙q�O��c_x�wwI7d�{�pB(��O��J��FQ�s�Q��]��ҙ�-�0�˨�}Q�� �w@�
�؛�����59X��
_<�Ta^��O�yi~&1Y��f�4���#�&F;�#�|�����D�p
>�ga�z�,�V�,\�i���,����}`�ʥ;΃�=�ic~Ԟ����^.eڦc��*�N߃'3�o��$d
���+�К��c$ya�44hGj������O!���I�����Qw��ycR����@�*����F� ��y�u����r-?J�+wqt�~6;��`�W|����v;�;�%n�Y���2��B�9�Ayd�1B�'1/O�
k�������	�'{]{��)�t��]L��7�A7�%�H3���9B`�i�r-DZ ܍;�]��M�#,vb�T��O��}wD6���Y� �i�v���].��Õ�'��{�t߽.��'��Q�MtD�fA�H
�? ��
��ǰ��� @Ag{@���G�[B��s�[q��C��7[]���a��k����@��aos~�
�+�g�t��wP�Ít�����ZW�:���5��Ϲ=�؁��pQ���+0��e��ĥ���c�,i$z9�"4Yyz7��oӻq6
c����K'�~�p��<M�����eA�N�	iO��ȇR	���ёW�M��e7I\�$����5��X���טPq�P.X��n�#qd�;"��t����2&��s�c�XU�5�_?�1�dY�w��}$���
�!T[�ʮ��C���(� ���X��y�a���ֲ5���qy�4'�Y����S?A/�ͱ�<��␘C�#�Ĵ�֯܄�o��O��,�t��8?�������x%�sJ�Đ}�xi�&a?	0ml��x;����ia���E �!�R�rV��n|Du]��4�DL��b��:g�ȑ��(IqXO!��HU��� �Q�e�Dԏ���.����Pf;�π�l��P�����O�w���T	t���}�@J"|��}N����w�o�1���x�3��'���溆�kd?�y]C�<(�~]OV z�QxiN�1:�}��<�U�us�k��5�4f��5�M����
}�O.�B-��	�����33�:�t����qq�s����4��R���U���p�c�\x�u4�}x _�g��Ċ�IśŊ-7H����b^T�r����3Ѵ *j��n�T�ᇎ����˹�䷿��+8�G i�^�E�����>D�׆�dp�Y��dED�i���aZ��d*�x&S�m�U���c쌏Q/]��I\���0uɮ<~�n�w�|�l��>qn������ԑk*D��o) ��X}�#��x�iQ��I I�*9BU&U����Y�B��O���.qM�L��\�Tr@e���9�"U�)T�P���bU����bU�C�PO�2NS]
�G���5���4B��RS�X��7x�����|��=��!Ol ��e�o���*���ˁ�}s��>���n���P�ib �m%p��F�D��A��z���cI�8��0{�\Զq�4E�����$N�sБ���p��;�����菄s��MAfĴ�gF"NA�"���(�뚬b?	敛�&�'n/<�q-7PM"^����Dއ!�����R)� �]�=d7��+���kz~ l"i@��������C�d��q1����p�183Z�;;�p8��7�B�I��f*y%�D�m���amk�^�էklZ2r��x�����|��Ҹ����)�# ��u���	u��q[c��H]^����B��-�B�ky��&�Z�ո� ؎#�d�PWoNKB�vP�TyD4��\4��ё��]޷4u�Ǻ��T���A�Ң�͌�)́�+������X��[��>��-�t����������g��z`?0&�,�t���QW>�(p��(��sO�Q�X��3,�Q�a��)r
 3�ZC��������~4V]/m�����A٧��M����=*ė���u�+ʅ[;뒷�BZ�b���wYg�~-�)l��U^���O��J14�K��!����l$h�;���'�9��#U���{̐a�iZ��C��Ѯ_6�@��w��i��J�=Ʒ���e�C��vD��$�K|f��Ƈ�gC���6��;[���3�9�<��(���2��@S\��x 
f�pgZ>'FIr��H�>�g�~UԒ�%N�&�8paIVR�c��'��)^����,���$Z�8Wd�
ᄾ:�j̗F�Y�b�B�c|��.K*��l�o���F|�����?�7'�\G���u�~�����S�-������Ͷ.��i����w#iw���ϯD�W{��[B�2.J��G���yA<��p��f��)#���uB��oi�[�K��ӣ�)PΜ}a���1	� i?����6i[�~E⚦��?r�@D/�r���@�&T�
��`^1�؊Z����&}��sѸH��S[a1B��~!H�B�Ā�l�^rrQ��H0>�!��|wFp/�6���U_��c�;���/<�7��@ps햇]�`p)i���-`'��ȴ'��i ��HV� w���~�̔O:���vr�M{�3�wԇ���O��09
(�h���"}��nxsd�����H� �j_�q�8�z�&�A	�'b6����"���C�W7G�L:aiN ҄_���NF�%���o1�8Q�F������:I����y�� ���~�:;.q�.zd&����r�]�/�G��:��&n�W	�L`Jm���myL���.�n-�qE�{��MP4����s~�߱_�� ���m���&�"1�b%�8Ҷ��|�_�jq%љ�e`���I��Q�s��g ��}=(V�qui������?�㍀`��Ft3�굳{���5q����#�@g�h�����4WA9��r~�����u���#�o��0F��������#ș��Y�W�<<ʖ�e���;�  ������[cĞ��sD�]���:��9m�m���(�z�W�D���$��8� -g	��N� ����
Wx?,��)���#�î�ő�hp�S�jm#�k �e�.���Ku��|�3GJr�#�s(z�d��T� �9aB�U��c`�xX�T�oS�W�<�i�~��{��Q�I�����S@�v�u���Y�.���1�l�l��p�1o���7r��G��G"{�TG��Dۣл�g<�+��X��;��~c���}o�o��#��w����:���9�]�&\qra�K�x·u;`SvæX>��	>&i�/1A���0���ˋ�*�T��fJ�J*���A��2��v���b�X�
^w��~	A{xw��~�p佝�d�xlG��٠`_�`B�������\����y����BT� �Ad D����(� k'�	;c#/(D���"�9��P1�/��t�5/D�&��R���"�6��j���������z��;;��ȱt5;ƩG�^BDht㮤�h%�=����a����,��9b|�
2��Ȗ����!:x11�|�	^���� ��MX!�[2���,i$֬�W1��Jj��ʐ7@���p�O'�g�t�O*mqv���%�ۑ�\���fM�[m ��o��`��5��DL#N�-��Ε7gq��et&[J�J�l�+�Wvᘨ��~�tu}Z@����,�ˊ���K�q�L7��F1\L����7Fp��3d�[�B������݃'D;Z;���.�����s'�Ļ�h��t#���%�h�Ym���^G��<om��4MlxJ�8��<�@dɳ�'�J%]�N����L��S�9�S5SNp@�?�H����Z>42P���4'pU�qge�g�l��^��v��� [l����}Po�iB ������[��t�2/��ǧtu鄆uR�(���|�3S��,1��a&(�/s#���@
���$����C���S�b��ҥ+�f﶐�Bڋi�~�&=%4��t;��\v�LLma.�\�g:��ܛJ�S��G�驼�I�~�9]�W���?ъ�Y�:@�R�J�A�HBex�&=y~���޺�lR�No;=�� p�g,B���S�!�n恤��a".�D�)��˿��Iנ6$t�y��7����~��}}v��F�z�4@�lY����AH�R�9p��[��5�@�B	�u�p��s0������}q��X��ġeO��!�0�&w�{��򮰀�5GNu��v��L6s�@ J�\&�s?��m�m,_� n
$����B1?2�4�4Ip:N��aCt<W7�:��G��;���E̒��s@��3*����!���ZsM(_�ڑY#t��17��b�%����ѻ�,�8h���gڦ-[���p�_�,^��%2� ����sf����ѳu�l=���~��!��G�M�߰y{��j��dޅ��{ͻ*��j޵C���܏ï��D�C`a�K� ��U*7����Th�-�i>@2	']/���o�������,��KC~j≮$�3�Mz⣂Z�LN~���
J�	��L����hy���+N}�'�XOR���n��G���/"�Ε7�����J���u�4��P��@�u��8�7���x�+\'g;��%�����#׏�b�C�A4�r�,���5��y#�� ���@Z��y2��7^�lQ���b������(_�`ב ��<+�s�?�v���ځˡ��}��?��wa���G�M�{���&ˍc��[0R$�> *�Γx�}���6k�����UA6T�����P�6��x&�	J�r&�f`^Bw���3��dR����e|���۳�;<���%�Bc�O3B%����#���&��[�nS�ʘ����>�~�s%��Pb���׵~(��
\M��K�}:+|c"�c��M�
��&�`YCS�������ᯜΖ�-�4+����MϷkH�B(�A�70� �Ӟ�]�����bV�VGT,�愓�O>��7D��>���?���oƲX}/!RH'���|_{Gt�;���	�l���Nn��Y"&~���[>y��[,�Tv����hO�K�ۯ�Q��݌� �w��='4>B�E���h*L��8�(� �M��6����)�y/�%l�F���#�]��(��o.�Fi�N��a���2�on-�c˛�q�f�8�h���(����V�M�hl(� �P��n���`�ozC�}3os��J�F�\Y����U�FIg��Ӓ��t�|�
�ts=֕��zs,�@f �`���<��W0�DV���y��ⶠ �W���s����5s]`(l:Eg���/cPr%����\�AX`�����wƛ�C^V����C��~�p�&�<��m���l�.������þ��$ަ�����˞�^����B�� ��bᾡ��{��$�e�]�wb:r�1͡BO�/Á9IT9�~~�3Q�-/�|�ƈ7�n���H'�P�h��7�8L嬏�q�=�u��tV��^j�ř
7��s��i�{�O��浞LY���__�21�LI�~}�w,a��x��׹%�c]+���m�꾄Q�I�W�J��� �Ⱥǋ�sh����t�7�CC�q"I��Y�u��>@N84�Mt��k 妰C&��͏���4*�t�8��ؽ )��۾�[:��Q=����6�j�B���42%E��et�D����9)��Dĸ~l �����a�/.��t��׸���1�xK�rei*pr^8͙���R��1B�s�N��B��" VE6���|\Ƭ.#�D�?���It�&�!�^��37�9�霭1e�A�p���>T�2��	��@8�c�W�g�g�3���뇢� �*I0g{PUw�~}EFZBl6C#\K���1 Ҳ�_&���m1OT֊�����~�$'*ĕ@���͓ݮ$�]}k�I%���Eb-w���09�}	��R���dndA�ւ���+<Yэ�Q�J�t�N+� )��M�h�lE�4Z��F����s_� ��9���P���F�d�T��C�< ��zv:*&G9� .�o�o6��M�ϑ��935�z�׋���[J���Rv!٧6>�e�Ñ c��@�
��I4O<���IRE�H�\�-ڊ��g��^������ TP�� �4�nF�LP�J�C�Y*f����_Ǿ���KU!���]���9ԋ9Ť!gr��\!�-�u�ӫ(Em��P��Ǥ�%^���r�E��k�B2�B�^�F���U�r#���ɠ]�EPȟ���e4w>G�Q�!nv%2
q�%�0#O��Y�|z��뽶iF�b�H	9��)�$׋(1��HȰ�ENb8�JQb�h�o���~'����K�������G�?I����>I�?"��)��L<j��'m����ͨ��M�H��|h�e����l�v������ءɄ%GQ5+%�!8�"A5�<����t�Q"�D��W<ҟ�K{u2�L@P"5WfRJ˕�%t+���Z����j�ȭX�q�9my�iw%S��f~��H	e��.��u&<ܔ���uɂ�%��*�P��9��A)0V�Xr�6����w�Ć�x�J{O:Rٰk�TH��?7��N�H�!�O�"{�BgJi����j�^���2:z��)����O�~!~Yc�s�	�^�k���;���)a�0��\�u�7	�dp���ٌ��G�Ϛ*���)aw�n"s��r��^	���q�t�ڀ[�E����5�+� ��d��)����:�F�ѹL�k��61��UzO	��E|�D���@3�C�8Z"�2	�@��`�"�I1��g����m=o#A�оV�p2����
�?�I��Yx�o�җc�J��X�pA�����lQ��Zs���gҭm���Y�t��m�ϸ ���|��"��O�(�)_=iga~�q��Y'�^@OcWA*�+��)��CU��j�
	'Ka�&g����S0��䎐���S��6z|=>C{&º���]O=�(��y�oC+�eC�AZ��g�zFI����X��$T=�g�ٿ\Opn�x)��G�g+���J�+\Y�w��)TX.�N�y�g�@AWV.aW�L������fu���� !!%���K1:}����Bz���=��=����:�UR�j�� 7�ɰ��d`��}!�VH?g0�tw���jZ����O���K(����#��!�]K�U����� �������UO	����Q�]8=~SOp!����TE��V�Zߜ-���X�ːFw��������~B
�ی�����卵pȳ�i(G��/'7ɸ�clӕX&y3Dǣyh�UzJ�G�d�@�E&�.Ǆ�^�մv�ú�{���ڙ)1f&��Q�L8{�3g��J"<��tV6Qո���zi*�t�4�^:�g��\#*mT�Φ{P�il����:�cVG+e���� �9/3'��r�ĺ~����������!��/V�T�t��ăoTK�-CTIL�[��b���pp����B�	!���f�F�0������"��HϦM��� �������ӡ�2ދaW�4�*(eũډFm��Y��m7�
J��%�ն6��YJ�giF����d���C�ly��V��R:[Ig'��m��B�������+Q3ȕ��rL� ���4as'pvJD[L.��s�Sܡ��|�����M�:�+����"3��4XE.ċy�ܷ�<K��g�|��Q~����a�rkW���5�}B����K8��H^�C2�;KWl� �f��B����)1���t�O�@SL!Yu��'x����#vP�si���V��m"��2�������D��ήr���8I��F��}��%�N�2H�kx�7�Q2� 5e5/��"�i>,���y�2�6%5�o�q������@n�)�{&�W���'	� �șI�pA`��waƋ��K�W�>l9L�q�6�Q��
�7�����li�D�ɲ�B؏"`���+Z=P2��Ġ��
$��ǅ�5��`s�/��$�J�e�\ߌ��G���tg�F��>���#`
d��q~�{L�B�^̊0L�q�텐�X5'�E8����TR��nN(}O���8���`\tA)��"r�ο�ѩߚ Y'���&z��'�U�%x�t�(�l�BJI�s�
x.Ø�֟��qԷm���&��H\����v��_8��p�����(�2��� ���+A��ݴ���9�"�J�:|�G���]�D�A���}h|���ԟ�1R�r��U�e;�t�Q��P�c����/�٤���g%����궏9�ܫԞ�v�S�話t�!=-ȫRZH����\+��ֆ[��/�f���0��pO�/䡷���a���ko=��(�.�M+9-s{Lm�Fq����㼠�g�����4C�̑��R�w�^� ZC&�M�.��\$��U�\	A�w@OC�3��t�6�����<�����%A�=�@�<�(>���-��sd[����0������ȱ=�� ��h���vx�-��"U����7�v�<#����_���&����Q�v��ZK�3�;�,��Ԃ!J`�"��7��pb��j5��f�د�g�e��Ӷx��̍)h�zdm��!�Ո�s?�t�F�p�V�K&%�[c~	����㎕i�|�M��\1�_��}�����hd��of6����\�'��E�(�m�X�am��f
s �C�%� ��deM�a5�P�4ͨ3d�V*͗�dgй2&-�Βa`�@��39+�Nmh��P��tm����ZT!?�x�`�빙���o&;w��s;5�P�cnN@��jţ�d��³�8Qi<��^��'�4�4�w��*!���>����^&7�\�f��&�WVo���7��~��T�J���%�k}p܂����$:)N�YA:IN[��AA�q�!\���rH�hY0C2:��c�,e�/�H.���F���l���ޛ8a�2e��,t��O����Ԙ�95r,�A0iDS��,U����LF�l:�� �9&C��w�{����Gx�I\��F�;V�`�Rđ~�#=�'�w>"�<�S��8z��M�
�.ܮ���DG�4�۵D�S"��{�|��톇���	��(���`�H���H|˅D��6(r�Q�j-V��1La���J<n(Oa��l�w1ea�����<���{,'�8��k���0{�An=�(к���H���S�$�秬���S�	.ް��;�,VR>'3Na͔����XHk��+�g������嶕x&D�m�[#曟�1����&�7<���wI�3����Lo���R&�o�-�,�j��)���v7�4�W�<�ןx�3r�F��`4;��W;��v;.PR����� �M��k���Ol8�Ho���Lb�>=����FwQD����Ӌ�ׄN��3hO��ɰ"�s�E$$���G���dI�AAy��������7���Ϧ���8���� �a�t\S	qqS���D#�&*�A�&�ж�+A̾ ơf����ڦ�^&z���6���Tb��(s��Kg����̧��Rbu��K�m�A%��q%֥q�~��_�G�s��^7�|�Ol��`�Q��|��ʡG�ݺ���C�ћ��,���i3���������0k%��Ī�*.b^�bW����8U
�[�&���<|J.��Þ��Kr�"�K���9��x���Lm�2ߍ�hd}�&R�߁�d*꬟GR�A`���S�y�L,yJ�J�)O�__�a\
䉪:^�R7��ܤ�e�SZBH�Y��L�.�!U�~Yƃ����LH�T' ��"��q�c��v.�({f)�e�S�I�����}|�� �j<(�|�wL�Z�I���&���/�14rG)�P��q�����6��ô5G"��?�r�q`����Ck;��@|RwAndBx�L�g���u��$�O�̨3~9��j���\t�v��w3�w1���0�&<[���C�X|i��'G�"˷��`E$Es�EEO%���t3T��%�˗����R���P�:]{��av��rә��#��N2am{p����3ybc?�9�o4K����wk[A�*p��B4�J��.(�'�x������� hb#����j����Ab2���AK̵2ΥQAAy
�cvD�Y�`8sk s[j ssj����������P�q�#����7��J՞�@Qu	�	��Q!S�9��r���ǥW���*Jl��,�[i�6fFR��]L<�1q�\+�Y����������_]^%�� ��� r�.�BA��| �(�L&r>�`�$?�i	/�^���d�%�'�g�b�̤QW�Ii���z�5��w��TLrHF'ث޸�rHr	z�K�a^�iz��BRרM��:S*���?�wqn�J�爫�U��s�C�-�����ߋ����<АG�Dp�s������'������J�$�{�΀c󼊈��O�M3ءu]����#���G���b~��;O�I��im�r�;�&^���T��6jRh~���:B�=`���8گ�[�]\�:*���,싿wD_/��sqp������#�o�sc� �o��/U�!`%��,��7RBAE=P��/v�kA���b!N�3�����}n��9�2�?�AVs=�Jx��i9A��Ż#\4��� d��5	���K��ؤ˾�$�)�����q�ʢA��֦�`�9�����!?���[����1n���Y���C5�Æy����s��?o��g��0\ 7�m�;8Ѕ]�%9����<v��h�J	�{�[G<e�Wv����Ć�"�]ENW:�{HKe��Ku\�CI�d{�f�,�%f��~U��oj�׽~�ck^�^��WK��wq���( ���H&VC� �v�0� �V�Dv-�<v�8I���c�[���a�`�P���Jv�-���7��
�������F`ъH�^�)��K�	~�/7R���{��I����ɾ��TV��>CS�� �;UeG����o|佶�{%l�PJy
��{?��w�o�����L'Ĵ�#]TJ��x-	'Z&G�K��f�*91�u(�'6F�\�%����*�^\>�l��W�����H�x�2P���JK�1$D����='I��K|�ݔ�����O$>��M/�4ZX���+��j�U.�a�&�>iI`���e��Y�OY������0I]�ND�N/Jc#\f+	�wP�3�!\Y�(o�Z���J����$90ͷ3ea����/.��_���fK�#�W��@��:����͘p|{K-p�':�����N�=�!�Ԇ
���L�z^&Ao��U~�La	:r�n���HT���
ؼ���p]J +Y
O�yj/��/KvB���@��8&+ź�{�$7y�^h��J�=�r�����/M��>��ժ��ZF��`I��BD��.Q�hD��Q���=m��t��&��t�-�\��"�|T©�>w����moD���K���y84��YQQE�F���Mz[s�̩�?"X8��|�d��Άk�hC�Փ8)�-�S�eh!�&��l������d�X�������}P� ox���K˘{�t���WFg˰�`��՘�� lY��"�#�[���>E����I-ɼg��Y.S�����oj�6�x�����}�.�_b	��@���]��Q�|q����YXn����/�����w����/��6<3����r��#fV<ag���mf.�
��
f���6����W`���*q)�+�,���%�����%˕�˅�߳��Vآdq�~c*Io���糷��l}�u���:�~Y�>��Z��{�DsH\��k�q�1[1B�1<8��V,�~S��k�D�F;E�d��=�3��-�WY<؛�؂.w�b�Y#�TX@�q�.��U@�_�u.1m���й݈����3>��56�w�J�н_H�CJ[c��S�q���uP�	� ���~��K����r�Gt����PB]�Bo3{aރ�2�Ƈ�߁��ćP�ǎ���8�4H8�<�D`���p������|�4���]%��8����7L�'�{�36F��e >iXŵ)�P�<_8�Z7��]��1��cN<-
���c��t�;N��,�O�4�ڦ�QxY���'	�$���
 +ު���N����-��-$B%�_�~�NJ� $�>
>�������wOt=G"�㧱)��Ɉ�����k����H��$=���m�d�ے��H'�L���{o��L�tnz���3AjSPԈ?t>3̎���Y͌�g�g�P��g�
�(�@����9q�2�w6����36��x&����gҢ8��l�>�g3�Y���g��B_�l[�8�<q�9jUD�wK�(�����B�m�>�t�Ѣ8��(��<xi?����Cj�t�{ڱ���R.�p�%�Hg�Q_B��ېVB�:H���C�^��+!-��T)��h�?�� �\G]�t�aH�!�
i�%�J!M�t7$�r��+��eH퐆��A��lH� ���<���@:i�I���[HG ��6����T�R+��@h+�
R��Y�<|�yr�})�a�͐�n�d�t���y���ėy�o$9��|��R�Ha������	���;��l�,�t��øN���!�i-$/��!}����A�|���s��N�g�,H���A*���0�W!m�t �0H��)	�pHc!]�v~�$�6� �H2H�0��ڡ��A����Ӆ\�6�=�Cʅ�^x�0��<����P饞��T��T�x*��xkK�j��H&�x���z=E��%5D���x�ˊ�[�q�s�|�qU���|eEe��WԸ��q�	Z���
��K\��t/|�[T���+���2���ZOvQUq����d��7��֗��V{)�q*��yr�>�"7E���)����&T�T{+�HԛX*���z�|\_�I��Tx|�ڻ7�ST��1�%�Y��x�=��{�Y�C&ƻ��s=��`B��rM���D�A�AUK�Ee��jo~Yռ
Ϥ�ʡ^*���Ĳ��E��԰8(�E�{�E]��X]T̿�6�͜��9Q��W�`���������a�%���<���ʣ���WV�C�(�������ہN�V{�T����)q��Z_��̗�*��n%O�_PC)?;\SXfj~�d��G��j��x˪|%����֖ͭ�z�*,���U�Uy��RJI�\Ϣ2E�')$_ʩ�isk|Ye�e겤�����*��>.����*,�[Y\Q#),����DRXTY;���:	-�z|�Z�K��P��+.���
K��� >!OMa������bJ��w	��WCaQMM�oq<��}������긲UTem�\����rb`�>OZ��qӦ����Y]��VW��,�_诂-4�
BP���t��B�4W�?YB�g�Cc�<�վ��� �dgN@"������ݐ��xG�7垐�?eק�=%j� 
<��:�9��y���G�n9���)���H����v��#����z��L
��C��: ɢ�
E} �\3�{2����`BI�"j3���>�u%�#�dBe`�j���2�y5���nBՂq~_)�
��vg���*��'�#��(�'��T�Zς��c�+}�7�qS�Es=��><5��y�3�%F���Wx<5Ԟȷ�Օ5E^����!�5���5�|�)��U�au p0������5���_���q ��d�]/Y~X��j?�I�c�S���'�.vØ���I�,TN)�􌫅�<��2I���#7���15A�c�������;q�F�Z��sȃj�+��{=�|+�K+=�sk ο�o��(��dR�gjU�HJ��<�$-Tu�����P!PO~!ҥ>�\�	Us��J7{#�gx��g�a�'�'{j�_�n��W��j�3��Ǌ-��u��M�N�����*�ʉ���l�t����������FR ���(�?wm��M�-�)��Ս�w/�0���?fpSǄ��|>o�}@�k���ImYe�Z��R�'��E��'��WT��O;���5�Cxԣ�onX^�Ō2  _5�z�y
��6�@����Ub��Ɠ��{1Lu����(�K��k�H�Y���G ��`���
��5N�^��SK�Qk�n`H�@uȞ�zx�M�����TFYmM�oni'D'ǹ<����{���΋$�c�ZʭXg���:Q!���M���yB��a=���"ޗ��W]�-�"�
9+�[g��`�%>JMeV��G<I�C�|�dBm�����U݇s���Q������+4�� pԜ^@��sK�T~�/@�2�E���a�u�k����䋚A�
� ?U`רV��ky���ވ'"M5J��R-B�/��ؘ��� I�q9_#��>��]F��n��L�8WE���2���?qS��]j!�����8�2O-�*B$�q�7"����Qs�-	�1�N���ZC$����ZO�o^����_	;�J��q����cdU8��ŝ��
`n8����?�'����P�/�2j�"�H��4�$2�|��5��e�`J��m��qO�����-��$%���?���G^�*2<x�{ӿ2�е��_����O^��_�ݱH�?W��߄�1iN%]��C����>�Ӽ;�<��Ow^}����7�����s��Ak;޹�����k����N��鱼���}��U~��s�$��2��}��l�Ti�S��d$$������$�t6@I6@�)ҹ��,�H*H�S���\�ږQ��¼���:%I�$��n�w�6AZ	i&�4H)�d��5J��
H3!|��_�7��sx��>�?Bu��������$T��5�4�L��iȀuɉ�Q���=<��y@,;b�����)��z-.���㨆���7�Q���O�PS�	�͹��"x,"���cU�R<Us�Q:��:%k�iXJ���"~��{j�9���3&���l^�/e�ܑ)9es�յ�%>x����1c07pE���*�@sU��a~o�xOeQ�J���-E��c���R@<*+�� �o�UM(��̷��u)�O�~,d����N�����ƹ>�`���|�* ��ab��r�N�X^��@��;9Å�/�z���eUZ<��U쩝�-#�2� ��2����Sr�A�����	}^-ї�����i�N�j=s��/��g^�?L����-�vf��6�ut��EPvc"H�ѹ�_>�+��PUW=���=��l�\�a�����ZO�wE�쮞�f�+b(���!�������!^�|��fR���j��'��,���vI���nK��fyo>�|=R��+R�{�ȧ| ��QU��f�g做�����&yT���|���S���t�S	���/���/�;jBi����Tm���^ȍ��I|����P�.��H��l���E��3(����K�V�]��:�_uGD]��P[gj,�,|��?|SS&�]���R�0��P�J�`<cő����_�F��T����򑶪`d3��Y�1"±�"��Gr�����h�A��^���;�o,�5U�gg-���$���CN��rh����0_U=�{,<[D��S�Cy�Y1�>�~c��B]i��,���d��ǁ������<V������uE����/�P�h��)*�p�SHO��ފ(Ȥ��l��'�t�i���!$5
�#�/>ܰ�C��/�<����o?�3qA�:�v��~˺�3��K�?���d����6���餜��Q��H��b<O��ᚎ�w�]��6�NM���F���L:�n��A�B�R7E?M?S?G�I�]�p�p�p�p�p�p�p��...���(5ʌr�¨4�6�5n5n3n7�0�6�L:��d3��2L٦�&�i�i�)�<�<ڬ2��&�͜f�0g�'�]�)�i��9�bs���\c��������+�+̫ͫ�k͗�m�v3e�Zd�EaQZ�,ɖK�e�e�Ee�Y�,�l�D��2�2�2Ӳ��`YaYiYeYmYk�`�h�o9h9b9n9i9e9k9g9o�[V�5ɚlM��ZGXG[v�=ɞl�f�n�a�io������������R;a�6�6�6���l�4u�:[�ROQOS�T�Q�K���O�H�D�Lݠ^�^�^�^�^�ޠިޤެުަޮ���l�D��0�0�0�0�Pl(5Tj>�"��2C�a�a�a�a�a�a�a�a�a�a�a�a�a�a��ɰ��u���%ɘlL1�GGUF��d�ӌ��x�y�y�y���oζ�b�1�s,Ŗ%1�}�e���<��:��j��Y3��։V�u�u�u�u�u�}�}�}�}�}�}�}�}k�Z(I�dG�#�1�1ڡr�&�͑��pd;&:\�)�i���9�b�f�V�6�v��NG�c��~E-�����dK���Rm#l�m*��f��li��5?g?og����m�v;�:d�C��7K�����U�Վ��v���m��ɶ�v�v�v�v�v�v�v�v��ڎۓ�)�T��h�ʩs��6g��������u^p"���V�V�֚6�6�6�6�������v�v��L�MMGL�M'M�LgM�L�M���鲩��n��R��,7+�Js�+�(n�Sդگ:�:�:�:�:�:�:�:�bUTU�Um�v���ej�Z�V�����u������]�]�]ֵ��u�^����z�^�O�'�S�����z���������_�_�_�+I�dC�!�0�0ڠ2�&C�;G�yr��ɺ�z�z�z�z�z�z�z�z��Z/X/Z/[۬�V�&��l�m[m�l�m;l;m��"8�>���:#ԣ�*�NmRc"�3��6�6�6�6����v�v��T�����}�E�X;5z�F�:�e��A����� �[�m��Ҷȶ���m�}��N$6H(UoU�ʮZ�zD�V�<`�c�oT�ջ��wj��LM�f�柚�F��ioԚ��x�T�m�v�v����E��v��=�>ݧ����eB�������0�HX�2��k����2:�0�3>j|Ѹ���1�4�4v�Ǧ�����8X���)���-��G-�è�Y^��f�n���/�����0B��8d��x�c�Z������j���#�e��&[�m���6��-����b�b�l��	�~��ϧ�ﴫ�&{��^{��o�z���>0I��ܱ�q�ǜ�t�vt�v���2�Mu>�Wݢ*V}�����ՙ��Tu`�e��_QoQ�I���>�a���S��ߪ����nWK5rM�f�f�f�Ơqj��L�����Ti���4�i�k^ռ�٭�A�����Z�v��A���5m������Q]_� �;������2�����bXi|�����)S/S�i��Դ����)�L?�¦bK����N��g�o���[��Z��>��0{��C��`/9^w|�⠎ST;��LU��î�����P�R߫�8~F��������j�&Ms�f�f���s�M�o5�i^Z���5� �{uGu)���}���?���o�_gH�]�68��1�L�M��V����ۀ�k>`�̜b�ݢ�ŲͲ۲�r���)jk�J[���ٺ�z���Un`��v��`�A@�o�{�u���Q���̀�e�~�!���9>rv�8�sH�7~��,v·5or~����:ǭ�\5@5\5Y�UoWIԉ�ǵ��s�u9��Eu+�m�F?^�h6h^�lӼ����k��%ڏ�'���ct�x]�n��Q7D�~�A�� v{@�f���+���
�:טol��4�4�TdZd�71�U��5��{�z�M@��Y&>oi�\��[r`W̳��~�������M���_��\{���^e��G�G�À�}7:n�ew�Tt�c��5u�K�ɪ�T���T��G��q�]��nVQ	}A=C3�V��y�v�fp�N���Z�v	`�ǵ��/�n��G{I{Uۤ�Hw(Bo��7�'�s���2�����/����O�O��O�s���� ����ƀq�q�q����q��c�u�j�3��D�p�/��g ��a����Ɲֻ��`z���~�m��k[h[	���a�ʮ���m�g��/~����4G�c��>��N:N;:op��|������NN��̽Ur�NeVMRMQ�Wը�.~��J5L}`�ݰ�O����СVjn�� &&i�h4��i��9��4Y�{aoφ�Y�}U�O7Pw�������t?��6�8���:�%�af��;�r�zË�� >��9�)�A�!�Eqn�2?��1����w�v�e�ephU����=j9�s� |��:ڦ��,����s�����h���������8�?:�λ�.�Tg������RH(�[�R�Uw��*�s��du!p�����g�ߨ�S?�Y�Y�y_�d��ډ0�e�F�Sڡ��z�~��{�����>oxٰ8��g��C�kc|�����C�V>7�1�7�����Yby	8˷,;-{-G-/Y_�nj��A�$��6��~ۣ�=@�?��am7���i������K��M��{�x��Yc��p~x�+�/�����_5H���A���ս@�g��C��U;4��f�vPF�n��V�X�Wuo%���]�~��.�N?v���_�����vÝ��]\hXgx��aP��c��g|��$HT/[��������F�DUb� <�����i���Ls�e�����Zf��n��i}�:�6h�:�����I��9���B���]�d������u���X�]�g�8�w\v����8�NJ%!N�����X4�4� �[4�h.i�t�ɧ�̸_���b��8��dn�x�ˬ�X����`}��!�p��>Ǿ̾����U������f���J�P׌�=������d�]�C�[^J�hl:pNSA�z_}N-ꙡ�Ӽ��H�/�\;X����_����jC�6�F��!�	���B�Q� �VM����z�k���O�'���V�6��r��>C5�]O�h|��g���
r�w9HPF�?O�6n2�i|��n�odrD�i���Dê��L�&��:؋i�>�͵��/���l��2�^m�S#,c,� ?Z�->��x~��H����y���p���j)�k�u�u����i�q������ ��a�a�^������H^���-H,W�#A&*uT��U�	tn��.g�s�s��9�a�ί����I�$T1�A����ל��R�j�:ի��.w����Φ�JP���jV�<L�����5;44횑Z3p��y�#���_�}^�U;v�R��'u/�^��Y�[wP�W���������f}�>_?G_�_�g�k�������%}o� ��Wp�p��5�8��q��V�m�t�����2n���i��x�����i ��i<���=ƚM�͓���s�U q5�~�U�ͻ�-�V��
�� �Zam�[J,~�C��-/[�,�u��-�.>��������,���mZ��Vf��l� �n�} �i۷��lq�i�f7���Q��L?�@ۭ����2	���R�W}
�T�z8�3������i�Z!����ު}�;S�Ч�]�)�_��U�%��Ɇ� �� ��b����q��7�� �L��:���TmZ�#�|��
�9�����4��m����濙;�ɖ��C���z�I]o�Y[i��{����F��_�ƙnw�or���=��u<��� m�8�8G�)���y���&y�ੂ ��E��JBe��UiU�TY�U7���i��	�Q��@�F���I����igp�kԬ��O�w����I;(J�֧]�]�ݦ}8���j�n�!����OxC�z�JP���"}5H(�`��Կ�7���Y@I�K ��70]oJ���ۯ��hzd�M�����<�u�?��7z��O��7Z�L���~.�;��$0{���� �}	�搵Ú
p�d���'lo����#�� ����k��~�HW�7;������B킹��q�!V�$�΍�����6�Ǎ)j�J�r��A��Ũ�	�U5���a���( g���j�5e��=��V�͓�Ӛ�5�A�H&�[;S[�*�m_j��e����u�tf]��J�D�E�'��߁�8ըG��~�������~�
;9�'��1�o8f8i��p�� � u�	��V��e���*�d��x��w�g�3�`J6���~����`Md�oh�������bI��E@EE)ª�{AT��]u�u�ݵ+v�]��b]{Ś�~�L �������}6>x��̙�3�|���		��S8.u���ԩ�;r��1�_qz��d����n&���=��O��9K��b0"30o��U\k��wm�����o ����(ՓZJI;J��٬tDzQ�@�D�/�*m�&A���,Ŵ�&�7���B_ag���7�b��V��M�fp�]���̵��w��"�B�����H$�D�"�)Z���-z%�.vG3M4]�V|T|���X_b&	Dߍ��#���K�!Y������ն��v'��)�W��m���������ۍ����	����]M{W�1�>=�����n0^P�0-k���Q�8�q��z0��cz�kGS�Zh�p�h��N��.9e;=rʃ�6��Jv�p^�XPm��e�)�!�#�+ֹ�r����U_�E*�/�K+�Y�Y������p����M��#F�CSY
������I�m�]�c·B}3���c��{ی��\�V�hs���V��'�AP��D��귺��kD��.�<sB|I�A\Y�"i'��[(Y'�%pVrK�B��X}��Vf�ئ�N��g���M�{`�[�zvVp�G�N@������������D�A�րGN�������˱�cg���1�r|��X	3���/c�,�ߠV�;�t��8�_ut�Ek�9ov>��.������e,�j9�nsWK��a6�K[HE�qP���;��n��~u[���[��C7�y����	�C��{0O2L�.��^��I�e����E-Eb�/h@�d<�V���'����l�ǋǊ��37���_�߉�$���l�t����O�=IG�e��l����cW�Nh`�ɮ�]_�AC{#�����0ʧ������a��^���,��$�����8&�q�
�r���}�'N�0��Ne���k`6z�l�R����]�t�6um��
g��u9z�M�����]�c<7�zH[K�H�iP=�נni>"����h��j�9�1m ���Q�[8�g�p�p�����p��4���Ob>zkc"25Y�:�BE��������P���~⩘��b$_�,d.��#/Y � �")o[Ƕ��
t�];1<@{� �1�3���b�zFj�.`��L���+�a���N��.^�c�c�ڦN"'7���N���F;MC��T޹�s3�:�m@�n��W�Ղ�h�"r�t��J�
%���%P�f �c\ǻ��bj ���J��1ҡ�Q���S҇ҧR��n�ݤѩn��S���s}a�aWa8�p z�D���MY�j6lڤ�)F�G4X4B�Nb�蝨�8D%Nc>�w����[�W��IwI�d�$�q9�m����r��l�SE��M���l�cWƮ�]M���][�vK�v�Q��=c�H���]����mhC7o�@�.�3f����t{�c4��/N1�}�G�͐�:�}t6v���tv���"gs�S�2�\k��s����U��ǮF�*R�D�(m#"-]%݀�����*zb7?�^��#�Ƣ�ݞ�q�*��k-����
�0��)�+ ޭ}���,�^�|��1��\�El+q��H�II��VJ��mMh�v���,[�h�����c�Zv��Z�u����G[mb���}u������������o��`����+�"�;�u���áh��<����^8��(n���1�1�q t�B�u��o9>w�����q�{�4�L5Wq�g>�e��|��.�._]*������zcW �v����m�n�/=N��� m�X�$N��7<��y]X���Fdco��ʋj���Z�\��R�ơD�����mg�SJS�Ļ�0�֔ԕ8H�I�K�%���9`��Q�U�W�4C$��v�fa�5��nW�,�n��A�ׇvyv�D"�c�B9.�_a��~��1�@�;4w����0�%w��5�}��aoq��x��	���)��f�8-���Tѹ��Ʋ�s�s_���κ.&.�.N.n.�.��`�K"Kk.𽯮�66z_`Ψ(�+�JG0�}SZƭ���m��ƀz���eb�a׮:�2�qP��K���
��Ř��A;��DuE�E6�Q�(I���{@�L��Eqq3�P�C<\�!i՝.�,��V<"� Ɂ�~-i`kmK��(�4ۉ��0[������)�bU�ܦ���v+�ֲ�ۈ�[���_��g� �em��a����9*�MN.=?�^�YL�M�8[;��E˜GB�Lu^ �x����c�2po�\,]\:��qIp�˅���u��l��k\Ϲ^v�����;�O�e�r����+KWH���܂F|���f�CJq���mn7��]���P6��v�g�W����:&�$�eck����f��p���_hn~�F
=���4����{�^���[�]Ş�ǊG�ǉg`�y"N�Ǭ�����)��b�Yf��B��jp���:�ug�}����v9v�17[��Z84t }��0�a$k�g�k:�`TǢ�q\���,�N��KG#�*N���9�BӜ���D�T��|���s��C��h�:.�]�.�.�.�\.�]��U\=]�X��t�s}����Q�-�eZ1E:�f*��%�"5u��&t��L�խ���m9z�n'��q�ѝ{/�hɲp�#mv���b3}��Tl���N�Q�%H$U�=$]%=%W$ul=y�,�ۊ~v���m������_�wu��pD{]L�7tr��_�#���mGK(�UN�Γ�g@���|���s�se��.���c��T�Y�[��I]��1&��r%5� ��3Y�=e��Z�?\@ {��������/(`O�66�l�l��,��fs���3�M���Pr�m6�^�1�y�s����D\D�x'��uqYIeIm���]Җ%�
��3 �MI�����Z{��$(�4(�-�{�|+�UF	��a��ޱ�n��̞��b$a�h?�~����C�_g���4��S�[���3�N�C
{ݙ^k�ח)���DQMh&4���\(��
��ڨ��Sh{/�N��6�6G�tOۜ��l�ms�&������-���H_d(�\,3�ޜ��=�{�����������=�����6U@6ž5OY��X��7?���$�V��N�3���qI�'H�#�YDF����[�HL�������dA�`��Ȩ�_ǣY��.}{{��'M�i�2V.[���+`��YЏ-o]����d�R~�������zT��#D�3���)x[�KA}A]C�`�.��6z���[�G�����.��y��0z����i���зPm`�Q�U�C���J`�'�/Kk����6�	�����R܃M���R� !�o�R�BS�s�t������[F�?�����د����@��2�ې;w�IuG��νebRb$�W��f�\7�m�>Mbg9��O�����{��Tܡ:�9�t�/x�����\	�6��t<@m���Gc�L�=-Ay��� <����Q�CI�\ez?�3U�*�ϕ������~~����	Djǣ�y9j����Q6�O�Q���)������׿�ĽIX��f;_�2ܖ[���W���;����g[^d�t�ŗ�&\����KW.�Εժp�����vr��ar�
;���cV&����r�Ez+g_ee8�|�6��	n��'�r��4��?�ʕ����/���+����&c�����^�r�n9�_ߠ���E|=��r�Y�L����b�l���r�g�ϛse8�쾐;��Z�r�Y~�0����v����� �{�� W.~�?ߜ�^U����c�=]�7q�����_B�n�z����φ�/=��%<����?._��^�~�辟���Ǧ�7����&ן¸e��\)lȭ�ԃ[~��[μ���So���O	���l�ޙ��6R���O�gq�Ǖ�nq�.\)�ʕ.fO��gN�R߆[�nȕ�M�2�_�>����>W;ʕ!��q��Ҋ?NVe��Or�ǝ���;n���\��_��m'��W=�f�Md�aɕ�G_[E-�p��a6����_�d�v�|V�L���I�sYy��l�d1WN�c���,de6�|���U�����s�s���+��	��/C�RX�+�[�������ϩ�T+n�������D�y�9(x��2g3W�ґ�BY'V^��έw��Q���˪��,]�'N����a
����}�j������C��Im�.��?���¯���f����������=��G�AC_��T�ӻٷkk�sb���m^���t��剙;��hd���d��W�mL��78l���oe�����xKr���j�w[�|uk����]<�����/��;��9w�Ś�^��4���#\���}�����q��D��♊U�����q���Q=j&���p�~өZ?�Y�v�
7sDN�}�X����״Y��e�/�J��};�}=d��-�Wn;����^�}��	��12���"l��w��»�s*�]�<s^���v��3iI�сG��s[o
�S=��/W�v+�/[8�͵���;���J9^2�����ǧ����<����߬
���7l�$���Ֆ�ݗ��S\h���>j\�ꗗ�������	����v��iں���N�^+���R�Bvn�)s�y�)'݌unܧ�Sub�i�=:���d��sg_n{���:y���ۦ��h�k�|'�ͫZ�49��G�Jk�����Y����������r���z�O({�fs���G=�8ru��m�Z<�hƉ�/�8�oh�nSV��Ԡ�5���=�j��q�";YV����{��>�EF��6l��A��:4C�����>}�����G�Å� ]���{��ܬ��}���ڵ^�k�>z:p�oSN���7f̂�'�?>�ŧO�[�v͛ܦ͉�/_V�X����˗{�-]��g��'��?�|��������잼cǡ�_���Θ���Q�_���u��������ӧ;�J$�W�x{��C��W��0cmvvR/�����n���g?غA������Y�����ƭ~�m{��e�YU�bW{Ԩyw��s=��ר}��q#�l9�$9yQ�r�j�IM]Ҽ�\R�VK�ڵ[܊�߲�[���/��<0��@gg�W�Fߺ�l`�&C��_ڳU�Uǎ��2(�ݮ�Ϣ�=k�na~�˗z�7o���{�g��eƩS�{��=�ѱ�̶mo���)$$7�ܹ�{Ο�s�ŋ�֬y�����㼼����-F,�T9-m�D�s�?~4���-�m��ы^���x7\�hw�U��/���M�e˾�rw�4�2e�����-,؛�� {��~�޽w�����7n${ZZFZ��*����yS��ŋ�F�9�gV�b�FU��~���������g/���}�e��3������_1b�W�6YQQ�v���f�f���fe��/�9z���:\Xv��H���c��6�<u��
&�Nj�����ϛ�ٹ�u�j.�߾=xoϞ��W�Pg�͛o��8G�D��NN�/_w���͊eʔ�YY���`ѡC=�]��n݋#�z�t�6m�ͬY�/=x`�z�`ŕ��)���������o�NFƤ�W�D�o������9�}�n[׹�7oߖ=��IÓ���2�͆�M����}�eJʄ��m�2���ܪ�ʕ���m;>�ر��rs,���a�r�|i�z���k�gľ}���q�'��$$L&�zؾ��阘5Se��2zz޿�1�T�ʡ��e��چm���cܮ]�k�7m���!Nu�4n�p��w�:���Wm6g����+�/���Y}�zB�ɓ��3g��b޼?\�֭o:~���[�?{�wM�N� k�w�ћ4iJ�%K�˥���edT#����=���y�|l��1��̝��[���W�iөU��_���s�y��N+ �� �\   0 � ��`    � V ��� @/ � � � ,  ��� �) � �  *  O�� �W �	 p  �  �
 t  � � � � � �  �P �-   � @  � �@   �	 X K  c `; P � � � @#   8 , j  9 � h l � ��� �?  � � R `  0 x � 4�� � @=   x � Z ��v �m �2 � � �  M�� @u �( p � � � & @ `4 � � v ��7 �7   � � � 2 @ �  ��H @ � * �  ? � ` � � K�� �# � x � �  � �� �f �, `1 0 �  � b � �Z   8	 4 . . �` � P  8 ��� @] �& P � <  z  � � `% �
 X � 
 @ x ]� �$  
 � �  � �O @Y �! � � < � �+ � �? � X � �� @G � 0 � X  � �q @ 0 � �  k �l �  � �  � �0 �# p � �  ��] � P �
 ��= @ � � � � �  �/ � R �! �    �  n  6 �1 `' p �  * � �/ �U �	 � � � �� �k � � 8
   �7 � � \ � �� � � 0 � t �  /�� �e `) � � , �L ` � � 4 �  7 � p �  + �� �+ `  � �  � �> p h   � �_  �7 �, P  � � �� �   ( � ��Z @m   � ,  g �* � h � Z c�  � @�� ` | 6 ��_ �S �~ � h � ! �9 �< � X | �   @ � > �G @ 	   . �" ` � X � S �� � � x � �  n  � �	 � �  �3 @E �* �  f � @ � �; 0 p � � @M  	  F  �[ @} �) 0 �  � � ;�j �m �' P �	 �  " �	 ( � e  +   8 \ � � �i �, � 0 � � ��~ @ p h � � ��� �    l  �� @
 � h	 � +�m �1   � � � �v �> @ L   ) � � d � � � D  � @ ` 0 8 �  w�| ` P � � ��� �< �. 0 x � : � � ` � H � � �# � � < �� @ � �  { ��  ��1��|�����!����W!�oC�O����ׅ�?����/�������O!��@�׃�O��������d��ϐ���[!�� �} �@�A�?�����������/����w��������!�/@��������S�C��Y���!�@�!��!��C������o�_���������#!��@�W�����/���������;��r�����; ��C�B��	���*��J��]l� �����!�C����?�7�"��L��9��� �� ��@���� �����o��1���!�'B�?��ׇ�����?�!�;�����= �GA�@��A�[B�'@���������������!��W�����!�� �A�����o�?�%����N��_ ��@�gA���A�?��τ��	����7�0�3���I���!��@�[C�����:��z�����Q��r��j���!�+B�� �wB�/��������������k��+��
��x����:���!��C��B�gC�������$��[��6��&���!�_B������w������?������\�)�������F��Ɛ�9��� �@�����
�_���9��!��_ �7@��A�׀��������:��3�����!�WC����C����w��7��?�?�� ��
�=������ �kA�GC�_�������n��u!��B������߼���FxDժ���S㞿:��s���W�>��mw_o���S�����pz�w�~;<���h�S��z���kٔۛ��6�]��ϓJsz|˼{�U��h��U2Z�^����czS��2�>ց~C�fv�qyj���%ߜ�&�Ody'J�����)sC�}������x9a}��b��u�y����Z6cfw��
�9jPΞ>�~����a��	�ؐ)>_kμ�w|���k�.5Hl�{�~�)]b:�m�%Ϻl������%{�B��X�EW��Ϫ�	�xμ�MS����q��D�x{����+$��Y�m��eЂ�o:-6�xW��}^r�ԧ���/����̾x��Rˉ����R��������}���e.�0U֜����ǳ�ݽN���pЦ\�}e�����ap��K��o3���q�غ'�!�F�K5{&�[9a]�n��VR~6Ns���J]����_��]i9�{�+��N���<��_�۞�z���iGe�q�bi�A��̫Ԫ~o��򙋛>t���U�v�:��Ux�8����vU��:�˫�i���=���e#ÿ~�i�(4��^���?��(��<��ح?�}����U�5�['=#�L�ή�>�Xe���V�/�q���QT�x�%��,l�����q�O�����}W'�[y��S��Q�W}�td�K�Z��7Ϯ/��b�o���.�tr�9�+ح|7�܊!��o���m���͝<H�n�K��y�#Z�z�Q���읹-?�sx�E=F�;?cX�+-V�kXekֺ��&f�ϝ�y��3�R��w5{���:�~[�hV|���{��0�}���y����;�dQ��M6�j�|�Ʀnl���)�]�)o���˘�+s���$�=������Oo|y&�R�i�[�����b���5��~տ�����~�L�}�y����;�\���$���˓>W�h��w�n�o^|l�Y��j���]��d��␮��&�UuI?����'l�?|6��f���t��:�ͬ���I��}8�$���w\�WK�9���7�w��:XI�Z�V���Ľ�V�v�U(�fy8��`Xq���m�Gu>8u話WD$��������   ��_�S �+ `- 0 � � � �/ �5 ` 0 � z s �� �. P X  � f y � � p	 h x �  ) @ �O � �  l � �1 @8 � �  c s `&  � � ; � �= � � ( � � + �� � `7 
 4 � /�% � �
 P � ,   "   p �  e �� �G � �  � �  @ @	 X ��� �  ` 0 p  n m �� �	 ��*   � ��� @g �. � � ,� � � 0 . � �R   � �  ^ @ � � � d i � � �
 , � G 	 0 � � � �I � p , �� @> P � � �  O�� @_ `. �	 �  j � � �8 p � � �  k � � x   � �^ �!   �	 � � � �� �V � � � � � �� � �
 � F  � �# �: p � \ 6 6 � � ��� �& � h |  * � � �  �  ��� �N `$ � �  � �� @7    U�I � `2 � < l�g � � p   �' @w � 0  H�� @ � T  � 0  � � �  @   <���h `9 � � �  ! � �	 �  � �k �) � X t j � �L   x	 � > a �| ` � H ,�8   H  R `  � X � � �� �   F � � �b �  | � � �% @ � � ��C �P �  �  ~ �  � �6 �5 p x � z � �  � p � � / �E �	 0 (   � � � p 0 > � / `! �	 ( �� �s �< ` � h�� � 	 @" �  �+ �# p X	  -�� �_ �� �4 �( ` � j ��� @ P 0 � � �� @M �, �'  4 � � � �	 p � � n i @} �2 ` � " `	 �
  � �} �: � � Q �$ � h L �  �� @ `4 p �     ��� @k �* � �  l F 3 � @ `. 0 � �  ) � � � �  � �\ ` ` � � [ � �L   � � � � � �   � � �   @ � L  � �' �-   < �: �E �3 � �  * �   �1 p x l �  I �Y � 8 � � 7�7 � @ � ��� �/ 0 � �  �� �X �   � @�w���_��	�����:��v�����!�'@����� ����v��ې�!�} �{@��������_���� ��,��ː�!������!��!��B�υ�o����%��	�������!�gC�����������G����)��3!�!��B�'B�߇�������
���%�!��]��g��!������?�����#����������!�+@��C������/�����O���i�� ��!��!�kB�_��O�����	�,��_���!��@�����~@����A�ׅ�����������<�,��<�+�����3 ��A�׆���������&����J���!�[@�W�������9��2�������ސ��!���� �����	����*��X��4����� ��C�ׁ���o�?���j��ʐ�m �WA�/����_�<��u��I��s �WB����������? ����`�����S!�[B����_�������	�.��M��3����O!�S!�A����������-����&��6��M!��A��B��!��@��@��!�_A�{@������?����4�������~��!�[C�/��ׁ�����+��t��ǐ�� �������
������]��!���!�;A��A�'A�A��A�߁�O��?	�������u�����֐�J�G�C��l��(�����W �e���ϑ'$�H��|�L���_S>@^��7��5���c�/"�H�|%���ɛ�W#OD����?�x�W�{�G#?Bޑ<?�v���]�k��'?H��|y]�T��)g���|e��(o �IyN�0(� �K�<�
��'S�A��rUFAޚ�:yS�����#IY�4��+��'�G9
�2�3�c�'%�O��|#�M�!(G��r�$G���e�/P�A>���o�ϐ_���2���){ �L9�q���)� H~��0�O�Y(�!�G^�<+yY�t(�!oI��v�A(�!?L>���M(����2�(�������PVC� e���W%N��^�>(K"?L����g(c����'ʁ(+!_N��|?e$�5P�@>�r����)�\��	�ߔ�Pn@y	e1��CS�BY��mQ.@	eN�)Q>E�����&�N�
�U�Q~@Ye"��P�D�e6�Q�F��22�v(��,�r�U(o��2����)'����(_�,�2��(���rʗ(�����O(��\�2�(Ϣ숲-�_(3����ʨ(����?yB���G��$oI>��5��E��o _C^�<&�"���W�� �Kޙ�	y5�D��ȯ��#�G~��y4�#���o'_Nޅ��y�����%OE��r�+ȧQv@����a����	���CQ�@~�|2e�{)WPe�ɯ�7%_O��9�E�O�쁼2y~����/�<�<yR�����7�ߤ�r�(P�G�q�oɟQA�e��)� �F��u�(� �Lޘ��͔c�'N��r��w��������}�ɳ���L���I�o�������)/�܄�	�/(ӡ����(!oK9e5�Pv@9
yU����샲$���)��|�2&�Z({��������SFBY��)� �L���E(� �M����PC��<4e+��P~@����P�D��S�=P�@ �o�딫P^E���P&B�eI�9PfCy�h�)#�l��(ʂ(��\����(!�O�r��(롼���R(3�����(w�|�r1�(����2��(Ӡ��,ʎ(ۢ��23��(/������h��'$�H��|�L���_S>@^��7��5���c�/"�H�|%���ɛ�W#OD����?�x�W�{�G#?Bޑ<?�v���]�k��'?H��|y]�T��)g���|e��(o �IyN�0(� �K�<�
��'S�A��rUFAޚ�:yS�����#IY�4��+��'�G9
�2�3�c�'%�O��|#�M�!(G��r�$G���e�/P�A>���o�ϐ_���2���){ �L9�q���)� H~��0�O�Y(�!�G^�<+yY�t(�!oI��v�A(�!?L>���M(����2�(�������PVC� e���W%N��^�>(K"?L����g(c����'ʁ(+!_N��|?e$�5P�@>�r����)�\��	�ߔ�Pn@y	e1��CS�BY��mQ.@	eN�)Q>E�����&�N�
�U�Q~@Ye"��P�D�e6�Q�F��22�v(��,�r�U(o��2����)'����(_�,�2��(���rʗ(�����O(��\�2�(Ϣ숲-�_(3����ʨ(����� �W$H>�|&yK�A�) /J��|��b�1��w$�D��|�]���Mȫ�'"G~��y<��ȣ�!�H��|;�r�.��ϓ$OD>��.y*���3P^A>���o�7����<'e�M��%�E�r��)� �K��*� oM~��)�z��ϑ��,�|e������|��ȓ��'�N���&��#P�@���?��#K��2�(� NY�7�gȯS�@yg�Ɣ=�o���8�p�ה{�$�K^��'�,�א�#�H���,e:�ݐ��L�|;� �ߐ&Ny�&�OP~A���_P~@Yy[�q(��\���Qȫ��l�|/e�%�&�K��3�1Q�B��@���/'_M��2�(_ �L�yd���P.B��o�g(7�������)[�,��ʶ(���2'ʔ(���r� ��_�\��*ʀ(?�,�2�_(K�́2ʋ(G#�Me;�GQD9�*�7PFy�蔓P�FY���P�B�	ee��P@��K��Q~@y�'��P.G�e�gQvD��/��Q^Gy	eT��PF��>�L�h����\���.����~�l:��!q[����Ń�����*��.w�9��������ы1����7��]�c�3Y�}4}L���ƴ�wß�j�x���x�6�R�f�����ٻNMo��f����H�n�땲a���	Z�]n���'�&[��N��80���(���s�+Ͷ��5�a�������hf����퇪��r`����{ZXLkq\�Z�?���n�e�4�JU��סG��/�K~���X_�z�4=���l/	t�G�?��
]]]�4�G��G���z��zV�.~��xZݪ�V��:1�a�{<~vϥ��;�e��x�J�آ�{�nb��;Vt�������������u�ɹQ��ŷ,�n��Sʞ�p�p�}��;U뿶���Ye�/�y�7i���q�iG�W�?r�������o��ժ��4�3��G�<��I�I0���o�����~�ne9�JfϾ�]���X���B�Ɋ�;j���kݮ�ݪT�Л�����Q=<�֯Ӷ���%�F~��&��|�ҭ1n�uFȗ���W����f��A��>�m-�8���;����(��ӭ�l����Z�xY�ng.L�0�YY���v�MFtk��-�u����FE���^���'��yѢ���~��W?L/鲫�s�~.�M^{���E�_us��Ȕ�O�]�	]5IR���)Fe/9��Xj�2�><����I&�	�1{��`�z6S���wt��_���=���\��Ɋ7in��r|��m�ǗCG�����pJ_�˿��W�6Uu�Q]�����Ǖ��?�w�`n{��SvotZ��^s��/�w�<�r_>����g'��/�d���P�hO��U���'�zCA�ZA`A��qga!�>:��,ܫ�iK������u�{���E�O`G��+}͂(�n�?��f;��u���A������|;	���Q_�}���*��V_�`�WԱ��R}W��Z���Y6Q;�K�~�ϬH}�%ԧ�����|r���;s�T�<ϗ�|���K]~��`��`x���yU���-��37�����ɑ{�.�z�&晟��(�P��D����rɟ�6�`
D�H(��n�~p�6������{��{���$g��M�NX���a��M�6Ǿ�<L�˪G� �}s8}9}Γ��ք
��������.�>����~���H<�þ�<�}�9=��l�-q$�_ H���w����'�%
Z	���B]������qf����ٚ�"k��7���X��m�a�6�<��"���6�$�+ڞ�XO��5�x�����m}V�e���
��/����\�Pd�#��ͲJ��>ZHη)}�z$ku�;�-@���У�%=v.����-'\�ۜ/O��a~�_ϗ9�zo~��T��uJ�:w���|�"h�>�Rv�%zx�'���{}��o��Ůڂ�H�L4~�`}&-揻כ�}�|?�F��?���۩>���8���7A��M"�H4z[�_��U��?�c��-T磭n�,:���}����Y6N���\�q��p�8Vk�Iߝ�����jV��8IX����g
�=[k�>�bE����QZ��u�?/�Kt:#�?��-��^[k�����?�I�|=qn1�����\��ߑj5Һ�J[��8\Y<�;��7	�;Xm���l�'����q�]�6�5��6>��(�̢��&��Ă�y��>�m����z{��C۱��Y�����3��q�M��p?J�N�<�ٲ#��f?>#��6�ޞ������U�Vq?__DT�_��~���,4������p�Rg�:K�]���_c��؃J�U��.��Ӣ�*Z/�離}���=�H͞CK�hUg�e	�+I�~������_qf�G��?o("_v�w>
����^(��j�}��ҙz�n~��И�J&�?i��n�����J��JR%�;�"���6Ε�>ݵ�������:���&�m����u����O���W��z:�sq5nٽW�-�|����Gq�8+�+o=��IOx}�/���J�o\���3�2�#W���T�k�˕��+Õy�P�+���+S�ҏ/���e�<���'�n��|�r[P�h~���s��w<W_��t��U���<�������v�Õ��r�/�/����[C�_�5�q�T�ʕÊ9_�+�������f=9��S���7�	�ƕs��o�zܯi�P�"Ϗ�ʷsU�����^���ޤe1^���!������(��dsF��3]��Z���yjmA�ه-q�0Q����s��Eg�����Q��c��T�j?������b�q���cj�Z���\�i����u�?;�ݛq�֥9W�reT+�lނ�W��\qeEG���<7����N�x\�@���qh�=�֋?>_���o����j|��/��w�+��ƕ�Ŝ�j|�Q	��7_��˽|Ynsbb�c�����F�ó^�/�\�ȲWpP����.q���侪\���]��R���VS���_�h�ux&��D'�����T�Jc��i��♣�|��n�y�<��ϡ��C֞���k��Џ[6���~���ގ�zo]�ҝ�N��qvv�Ow�����Y�a��C���VE�Օ?nגu��n|}���k�G5�^o�|��y>_���^~��ށErgZJ,!u����]�}֧#�\�+{��y��Aۖ������by��q���<��2�ϻ��^z�������ט��?�o�I����ͷo1�.�Ɵ��ߎ?�꺂��c�r_����\Ҽ��b{������ܯ'�_N�Y�~�I��-�o�Ē۩9�������)�iTn^�oh����X����k+�>JZ�{����ZT	�fz3HmTYU㢤��Q��g^r�AC6��â�S5Ƌ�P��W���o?h� AW��a��B݊"����������^�փ��E%�G��Ql.��L�x� R��,؝�W�'�|~2����.�9�.g9r|A�@稞>�E����W��kB�z��H�3
t�͙���N�yE�^P����I��c�����~�|�Ԟ݋�����*���A�
�m<o��q�q���@~�k�Ok�{ z���������g�����#���Xm��KD;h�fz�)Iй��26�Q��=����
�W�8/ׅ�<�g��__S�C�v\�_��"�(Ю�Z���mp��} �ˇ��@<�Z��
�͟�|��ڃ��� �����z���U�&I�z���L*�j�WAվOK�Ӳ���X%ՠm{?��{�8"�'�X]Ŝ���V�^�'�p'��;Jj�hF��۷4z_s���/�7�<?�Q"�y������1F��;`|��ʥ9��ϛ���:b��O�O�x����bmȑ�3OǰR���l�L�߼�����l�����b3Hп\'�u;�t`�"�1��?�O����1KS���_K:��b<��x�����������㱸���ƣf���x�bz5���H�����^�~�c������}'Kמ?���1�o��c��?��4��7���_{�.��{G��R�(6��s�/�5}�*瑭�J����5��Y�9����r��s���������j=���Q{�~� �8��e���}���j);�̪��������:mO�S���[�]Cp۩^��=�ٮ�h�g�j��_�����;ڏ]�7�?�]]$�u}��^�~V}ۿ�������_{>���G�y�H{��{k���d��s��Tc �הq�y���g�%�����ϝ5��qt��?�y�/���	'4_(n\�S�a�i�8�ɇГ:|=�����sN��K�S{O���Ҟ$�:�g����Sr~d�g�����R�qϛ�j��EǷ����|y�dn���[�H�1�R.������[�x�^ ^�A=����{4vf�0��m�n�#�����=���~b6-�(m��S���՗�����ׇe�*]�}<ثaa����r����YҋO������}T���ȗ]����\�~A���|�_�~�C�9�Z�Y-\���S}�»�~��u�,�����WG��׶gq��v��WO�v+�����o�|�����Sݝ�z���^��e[w��.C�(r��_�Ǧ�3���
�yi���c�ߨ�Gg����g��;?��Js>���z_�w0�AP�����ؗ�!��������t�����Qȏ����⮢�z��4�6Ū�~�����^�v_��j��^ّ�(�^�ן��J�?��L��@up^%�����4�W���k��֕�߿Ҿ_��W�T�i�K�ܫ�?�ur�kJ`�眜f~ĝQ��fq�/m���X��x%%|������)��mϿ�bj;��2/�w������2/��������x?s���6^�L����3������k��~�V{�֯~~�3�6_��כ��_O�����%�W�ۯ[����k�?�;HO���j��;�վ������U�u&��X�z_�*�Q�E_�Z�%�,�{��J%� w����nr����g�����+����G�J�;��F]�������Z���9���]���#`���X���c^C����۵���ʵp�����5�*I��|��R��G�{������J����K	_��r�X�Ɨ�J��S���-���_�TI�(���^3=�DT�Qű{O�Ͻ�p�@�z�jd��ۆ��d�OmO���(�������-�G�gl�fT��2A���Xֻ�nޛ�דTPO�_�=&Wk'�����
��ѫo�W߸�N	Q�hYD|T������<��}_��ߪ�٨�+�g{���U����W��&�����0�u��oԚ���N��Ow�yGEQK���պb��_\�<:^՞�����.~�6�r�.�&I�rB=]�����D�LJ�m������>W..Ro�1�`���Sqחb��_9�׽,�se>���?���F�y���K��[^�~���⟜q��G��1��q��.�~ظ�9�8�hn�϶�(�UI��~?z�j��R��㨫��\���?s=����zԷ/��<���_�^�`��ӕ*��͟��8���	w>�׃���Ͻߺ�>�hlf㎯�9IP��=��'|�)7���է�l�4�֗ P�{�S�2�ޅ ��߫P��i5�o]�;�~�����Ք|=1�7��~t]Ž~V���;}�\o=}���V�T;����>i���~����Z��.�ǚ����#s>��J���#���j�y����T��g�<珣�����E�����tey�Jש�+�=����K���J�/S�z\$\yމ+����1��y)W��q����҂__:���?f<�&	�^������ty���//�߫�{�c��Uϡ�5]9�&Ϳ.Ӿ?�n�+:�Ϳ�)�_qL5k�?�m���]��?�tģҽ���������\��F���YEC��X�-�_�k(A9�Y����Fhq�/�K���
�{z�r�����YsyS��rqeJ���"��׆[�i�z���?~e�������k���]?:��
ݿ�>��=�ϴOq�[U���̑л������Ͽf�:^a���+ꯩ���K+M�zU����������֟��ş���^x��߫����}��w���O�+�����Vҵ�#7D;����=���!�ޚ�~��wl�<�����9��=�eyW^�}?y>���{��З[~ʗ���Ǘ�#�x�W�Y�E���t���°L}{��T�}�Q"{g0�Η��R�9ω���7��K|�q�h�T����gܫ���DPPS�l����`�^�F�#J�jԟ����D���>	J���[N�����`��Ћ�,���Զ����K��E�Ꜹ����U}���R�>��D�5Z\�u*�3�U��X��u+�����50�����+��'3�i�,� ��K���D��R��6Ts�m�y?�/Õ	�r�0�o����N�u:�#ܹ6��(7յ'����>7��૱�g.���I�{�/1*!�o\B˄�^�U�je"K�[�u��~:Uk�j�¨�����ּ���P�vU*����G��o��Y�+'�ZE�'?1�鍟�c�Vq�t�V��'���,��* �����r��jJ��٣v(��=Diq�Ӂ^�>���ѦÖ2�?�(���J��a㱫pd�i�nJ�"K�����c�[���0�D�ܭ�ӣ�r�`X�O�ex[%(��2�&�y���TYr�,à^Yj ��}Q�m�#�_�����W��Eފ�k�sJ��l�����2Ar-�#OԊ���'��i8SYzkŝ����y��L�b׈�ӹ;���2�[Q3�*���*�,|���f�^��2�b��#أ�Gg�1/˳�k͂��5~�W⛸�8W�e��P��?_�����Q5!�ѩV�31����tx7:O�qP�J�Q��Xg0��ɕ�wd	eG����0n8���4|rM�¨�!�v��#���_p-�̴L�	�]|���訣4m����`3�4O<�;b�@�����
�e�S�0�E�s���{s]��L�k�k�3O���]^�;�X �+�j�5F ]B�3�	��]�
�U���G=2��	5.���2���Lq6�
�Ϥ�X�ѩKF�\���\��a?E��n:<�4�$=�,=�\�����R����S��s�o<v �ӛ�����(�:�'���bqCr>�8����mehK!ףg�B:�V�)��)t�ִʜ?[\M��
��~�E�^n�eݤ
�_�$V�U����B�>���qB��=~P7�Q�8쫸J�����DWH�L�(SLq���2��M�Y?�q���MaO����,�ʜ?*���)�
��]��P�C�R�vBn��~�|�3j`�>z���/*���jLd���`ͭ+��%��y���yzފ<��ص^au��2��l�{�	� kw����,�&�ԓ)N��)K{&�,S���'��R/���]Y��^t��C3ʫ�YJ��.��Ԇ�޺�h�s��.Vym���q�2<1frۛ{���geH�\Fiz$X��Hfe.�{�gȭdy��}3�Mh��*�u��������/�8��e�4��Y��W��w~�|�wl��TR�&|�{:��i��NtX�<��P�1���)W�8h�r��]^��0���jwoqT#F�j��}�A6����ӣ�G��p�O�a̘��Yu�"K}jA7 ���6��;r���.�O���,c��:t6R\S�ڣK�O��Ȝ�2L6��4�W���3�(�R�X���^p�Ӿ��~�Pk�y�I?E���Lٰ.�gn�S\��ڢl�)�D���#�*.+�p|�����`:w��ՏvT���d��ݷn =���[��4D7 L�WM���~Ui:�]���2簀�Gy5d
/C��*Z_���x�.[�oP-J����Cq��OB�;b\���ফ�-�h��6{��	��k��˝����� Uc�ze��˪kO0�ۅ���ː�rd/1�0!���4��);KN@��O��)����LQ���K��
3���e���������Ld�:&�ڱ�z����|��'�����9�6���4�Nu3�ΧV	`�W�U�t8����U\vp��+��W��):��)�P��ud�\s�0���}���.:Er��m̘��m�F�*:���2Fg��\_�\_'���cg10s7��,��R����z��Å'A�rf2w�ih���k��`���	mk"���VҘ��
�9���5;$��w$��0ޡo�ߌb�ue����B'9�'��R���X�d��oz3��Ð��� ���������,�s?��a��B���H6�AE�rg�9�K�����9���5���W1ԁ�:�}�ÐT�	�e�a29sѤ@�l�5F�sU�2��� �2E~r��#���u6Y��PW z�IL�3;S���r�Eo�z1����e�pO6�9�*�l�[�n�w��,���Lq����/s-����B�%�I��n	�qu6��IVЄ���Q��ke����z�X��c���$�0՞S��w��A`�&��G�ql��؈҇T�5S};�����cM�a���S�.� �Թt��e�:��&���`�35G��!�^ف�g��~X[�3q�	G#�����t�j-/+�|\�)�uV�T:�e�V���}^�(�)� Z�8�L�vdj<-����݂���dP���P���I ��I����[�b{�f���VMe��o5��۬��LP��L`������v��\YizW�:�1NsSR##���,F�Ǡ�"�!`����W t�@p
�zU|[Y�lm����Ê�t����n��@/a.��4����_����	-��WQ�&Usȱ�y4�M�Վ��QI�5{�&Y�O���-��0�W��鐑��b��Ch�W�Oq�_qv�vY�]F+ǰ~�2�)�!��&��3!��4�:hj��@5���JF�G�Lq���$T��o�,U����Y\�CW��b꯴��1U�Sǌ���c�P�
B�����K��R}u��鱫���N�ҽ���,���B&6q�����(�a�gM�YЍ�<����|�f�j������G�t�wd�>A��n����hG�{]8�K�8(}�N�{1,3��M�Od�2�Ў�	K��T��w7at���s���`�2�e�P�^kj�i��1įB��f�����c�V��p�Ĥ�/09��naZ��eJh������� ҇
7��3�_	�I��|A�3)��Mwg�I�Z9a]����䧸�{"�5��n��7�򚤬8Q��hj�nw~��,5_'��q���b�`_��٘[�7��iQ�(D���T�g��NQ㴠i>��@��囟
��iR��FV���5�-P�p �q�-�l���6\����V�6���|sG�(���<�M@W@�y�{��2����0�$_��ڇ�sW��ʰMW��<1҅�)ctǈ��)�%s��9gk�����X�nc�h�;�4�#}�%��j�{�V�e��Վ�j��`�$�{������ez�ܺ��j{l�nP��n`H�b��UJ��u+�
h 2�(쩚SR�:��0�O�nF�{�U���#�;�1�����i�{��ξ�x���řj�:���|��8�CW����`y�,笁�����b��kᑚ���x(2_z�����͂pEf���Ne���z>LK^9�C�<0\�)ab�/Ƴ�Ln��y��k�ǿ܊I`��L73��C�L��̊�S�%~>���io��3<UD m��hZ�6I0LaM�����M�}һ
i�)�`���<rft�+�ҍ�1�qg4�KQ�*p)J-v���)��D>Eq�~��p�1�@"��1V���S�y?U�{3��fNakL莎m��=�Av^PpKS;�(y��a�zm\Ž����8��2��IK�މ��L�Ҵa[yu?�Y?�L�Y�
c�1�@�M�����.�a�{8��4��R=�:�҄5g��9��kk�G�9+؜r�kN;�܇��\#��N?�c����������q_�D�=>i)�����"(�T	�%,	MaBS��ZťnX�[�D��P�"�%��������scQ)kAVQ��,OP'DdQ� t��{g�i����~���>h����s�~�]�������@ah�̦�נ����%X��߽6���	�@��7�	9�`��f��fZt|}"M�&7�]��)~'{W�}ώF�E
@���oP�1qꇤ�9-Hڲ":$�矓@��v�h#�z�i"�@<eA���Ɏ�B5�1�<v�;��;힣J�AG�B��R[���е3�[�O���V�&r
mu�m���
$\	mH�8Ė����	c�{��,u��]^�"��St;z&��FR_;�ˆ:R�eɛY�fy_N�5�/����e3��{����E������r_�nN���yS�r�Ӿ���r��F���i�p_J��})�}ͭ��J�/�N���b��8��.��BW�$"n;N�J;<ʁG�flu,�Ku�m�XR�=�b��Pjf�R�e�Jv�)�K�l��9�w7(r�
���ւ^8�'!�h/d���SlR��@Ђ��%R�f��W��E(\�K����b�b|Vf~V&���h��&K��J�p2	�F�~�p�c�����^�O��Y����p�TՌt�����4>���S�5aϹ?ܟ;*_6N��(5�P|�����MSo\�`2����)���_�gڸ�p���A��Ix�B������p6��+��$�?5o�)TB�/�~ُJ8��v�Y=*���{�����������r'��lǃ�l} �*�m�ܲ�`�00'��Ǻ&���U~6v}��Z��kF�W�;Qƶ��B����˒�L�BZ��_dT���l(�]��s#l��ǉ�;�(�e� � ��7��*����<Ʌ�@�<7~�������-�L*��%�ʗ�g9���"G2�����͂�O�27���>�r\�a(E]�&�!̓C]�"�{���c�x�q6+~f�tl�I������o������j�ռ�=ӆB�ly3�V%�'Ic�Lԍ���Ρu+�+$)��|�/̗	3��TY_˕�e!'H�Ÿ�A��ΓY>���#^�
�>�y�����,�ZI��� ���F�I%2��'�{�.7�.����a���o*����h�� �W=B\'\�+��#��A(刔�Dm(��U�X�đ��Xʒ�R~8Q'o�ް�$��m�<8|�ɿB��3�,A�Yn~Vx3���\�+(1�,N�)��	B��{�����PpR�];�چ�Us>�nJx��W�ƲƮ�y�l(k��e�twcY�h;�A���n���G��Vj�.^f��iu���Ol��F�?��~�E��չ���)��Z������*����^>�ueo�a�+�����>wK����P��y��PE�%�c�8��4둊�X?ȵXc3O��E��hdT��|�	tנ��Jhl?���Ի��d9�}�\�M͠�d;��Ճ����-�� ��gy$���{�m�T9���i�U�LŏFx����?l�Ӑ�1�h���>��Y���Dz�|� ���e����e���_���
���+y���kI"���ż��m��6��m���֫�y[�f�2M�:y�r���L���r� �1�� o²,)vax��'mRR�*(w/W$�]�	˄e�LƖr`2����ŢTo*u�(1u�P$�8�i1K��ԫ��!��8�9��8� f�-�����1"�3U�D�9-'u8)��)���-
(y����t�i6C����eb�2� �\V�3�$����`�?��Χ������E��2�嶇���K�G5�ZOg%ѣ�����y�c1�x�|cd`/�Yz��T^��`�(��Q_@t��D�zG=�N��e´�� D�|C\��4���[4���tݑ�iJ��0i�Q+Z?���T�H��h�@NZA�ad/Z>]l�t���u�u��N�NT����vH�6D��F���iu6ˬ"���q���ƅ���g�r%��7��aJ�o���&��7S9H5�N�:��%���� ;��nU�D R3�B�,������x���y�Mg���*���9���� ��������ꈦ�1�ȣ��_�vC�C��x��V`��!l1UR�
�_t��!/�A�]A��`/�/o-Kc#)}�����V�E�SKQ2Rˎ�v��K��8���-Q6��3��C�v��q��"�S/9�P�U^�EQ�+���R�4)�M����ؓ�w�5]��V7�wd��@��+�� ����} ���O�@4יgYg���ز�b�:�E�p��G�C��ǋ���Rz'o+
--IH�cQ8d� ��)�6T�]"l�7C)Ef� �7�:��[=~�A?m���zc�n,ݻ|t՚~�T�'�薂��,ї��v�bb��a�5�)�{Ƚ���9��߈��������w�\� ��m�������! �%T~ ��rjF�-���U[h'ᄯYR���{z�/a���ت�c��i���P`.>uo���1�r��Å\لh�W]����@T���N}�Jo����[����bmk��0%�(�9��`�p]s��q7Cd�b ���p]J�V9��8�|r_�ɝ��On���"��ۨOn�ztC� ���\���igS/��.�~���p���𺁄ѝ�H������tS��;*��W�e|��,��k�
]j�"�m\v�&�WO�����w�wW�s�q��0s)�}:�Pc(G���|���s) �Jr%М;�G���;@�sT�G����T�|�?B�%�l���v�X5ڕ.��F��
�
:3Ө�.ǣ-оɛ�^��'�*��B+ވ߆���i�]���y��{���y�jͰV%�+^�Ǿ�^�l���C�^��%(\Cm���yc_������>x9ykk�=P���_G������z�k����z��1��R�B�j-6f����f�G�{���|?1�UPʻݲ�? {#y3h!ܫ'�D�b�ފ?��w,��k�«*U�cg���˨�K�w!u�T�op�ڻ�ۺ�
|�f��z�pV֡.�X��ý��V��^�M�@y���)g����n��^�G>��K
ڽK4M�렌�ݫ%���?|�%�s1���![��1�f��˪ج@v�+�`���l9�����
ى�253�˴|e�D�Y���q.Хi2��j�I����iE�*'Y�R��b#n�̰t�����>�`Xh�"�Ƣ��wo�>5��ް���#�׽wڅ���M����"�à�B��`��m�,67��Gш�M����	˺J�OG��Q�)�(�F~�7�))G|���p�ڛ���v�~�=�nfg��/B]dM��)\^�cv��U����^k��,tN#V=�e�_�}��W1�*y)؜;���k�생+������:f?�m�p2��t��7y����f�ݓ@ةʴ!�t�~F�= �3���R�V8�8�����w���$��Ѵh$@��C��9�q��^��D�Z
A��_Ǘ8�ېφa��oDNҜ�.�m&=��֤��N�^X���yF��mR;�̦��' �u�>���r����$�c��Y9��t�!fs����%��=�.:z�Z�b�RI�o��'������)��j�=\���}Q�-�cWJ��[��wb�ٿb�����y��Swbg�%�v`�c-�܌?Y��s���Ƭ�xٝ���',;WR{@xj��7jURa�S[�pK�-G�Y�g3�pdW��%�@���)�����{q�p��$��M�Ø�:H��惜�����M莻M$�q:��<	щz�k�Jkd<[��>�c�)q����[�	X����g��w>�������m�V+pã_apʂ_p}.�!z?H�&�@d�#��|;�u/,�7zZ	�qw��jZ�ٽRfj�8�
J���Ìo�e�|�|ֽ�ծ�H=*���T�BV
��K)�Q"u�)�����}�,�c$#.vG�{	�Nb�v����Ƀ0n'�Tu����ʛ�:*��b���w#����cs�U������j�9b{B;�z;.���ۄeR���X���r��O�������+�$��	˺>���;�2�]*�㘵�]�#Wm��A>B�
���B�ͧ�b�Z����u�w��ƚ2*F�P/1�0&S�O�fX���=��/��������5�+̈́�<>EeM��x����	�z�T���i��B�x)x[�����u-��X�+�z#�Eɔ�YP/6 �<���}f����Ri����~��^��Py"�G��9��rd!'R_�D��A�H-�$Rs⬃Q�����Ca)�He�N��z��(���g��� �`w��`��O��^?ӂm�:{O\fO��x��6�t���e�����ϕO��'�6��j2P�e����)��(��*��3�����~�aG�UI����V�,�|��@z���>�s��Oq$��{���u�O�ۄ��^ �h���x?�����'�x�z��U�~��R���ثX����������+W���AΒ���
�x �0���D(S�^�RwED/��w���/ӎ�z��mֶ�������5D�)F��
)4��F�[qqY�M��N(��&��$��Η�H�>�]��:cw��>��-��\�~�j;�#~�c_��1T{G��<�43���9a��s�5��Ec���~����M
�	�.6���h���8��Fĭ����5W�~���I�s��hSܨ�d�����1\KwN�	�]�y�:�r��j���Q��Β4){���:���>񤩎t�U�~O�~��6n->d(�K��x��D�/�y���K �+�R���~���;*����/t���^��.A���4���**��0N�J<��XL�l��]`#J�k�tUTL��V�
�	�d�5,�W+�ȯ: kͭ��v> %�6#��ܛC�x,����P�>�G��>V���	�zOT�j�s��":�:�{_����v�H�V��,�Uy���yg�3�څ���*��?؂�^G�̱��4��QCGeT2�Ls����'
0�1z��-|[f��a!Ŵz��i�L~���}��?���6������p�/�Ƚ���XX�v����i�¨��'��N��d6�d��I�I��b/f������Q-�bH�/S�h��j'��;����x�Z���������ˊh�h����e/ �,�f4�L����4���ZM0|'M��p���3�yf$���8�e��\��ݖ����4d,��c��+j>[_�N�EE��ݦx@Y)O7|z<ٻ�ᨭ��>vH8�'��h2���Q�^�[G�a�@sTuЍ�u���5]�+�s*��l�f�xi�#iG��MP�o�Fl�Z$��tG��o�K�Q�o�8�N	�#u���FSr�./�UN]/,�)_�ʩ=�"��Js(7S�H���~|�݀=�[�U�IѶ����d+/;��4?��b�.c�oN��ǘf[�ĸ�M�݉Ӽb��4�/���F��ۘ��i��z�͘��w`5��-�-�ԯ�r��\�|G����x��;���뾜�Oy)H�Q���\�#�lc����'3H���g��^�dA{�i',���;��R-���LR�o�1ץR0ن2]�	ۇ�p���\�똿֪�J,Vu(��f�K9��44��e����[3;�6�[a,꬧��m	��R�t�K^�1�5�Ww������ٻ�P-[B�t��T�y��xS��JC�!/�u%�F�#c�Ъߧ�$�����J���=Y�ܻ��Aob���ڳq�eTW���_�/I��R�y�&�Zu����[����m�	ʫ���F���7�iq3�;bnפ��{��A��E`?����Df`���/�~�	؇B)b���O���I3��̀�������	>$3�v̭�dNi>��VP
p��@�˾&��7I����N>b3�6��H��M�ӂ�(��g�'��cqu�.9_F>
�[ jdv��xOd��Fe���d5F=>kŎ &G&y��$oa6�$��w ����E�-�Ћ�IQ��>N����~����5�o­��m��C�^�(op���ql�Ä+��kaő�r��R\�Ǩ'`G������#��ԩ��I�h^n��s[<#��Ѐc��F%>�����G�a ��<2���������&�à��n�I\.E���2(U���� ê��O�a,�#���c��/W?߽�t��HͰ7�*i������	�t7���hp�2�@5�s�Eo���M������� ׀��'CT�ȎR��"V�9��j�o�9 )�c;�;
�����<�/�o�ùn� �{�v�96Ij���5�GN���$i���Ճ�Ӆ�<��&����Ƣ;��A���NM�y!�T_R�����J��4��P,R�\lGU��m�_Soo}�To���ܒ:z�j꧛��JHV�A6CV���ʇZ�IŰ+lǐ˯�x U+=�:{Wծɨ(�A#҅FP3؀�IQ0X�n"�?��+�ިiΟ�i���Pjl�E���d̍�i#;��O�(4�Xy{�q�q^��,1毁�r@�`�zgq�l�\�`�|�=%�F�K���x��큚��������`�׺WOlۻ6ZO�#t���i�-K�2�
a��bї=_�f�X�����U�B�@T�6˪j��G��-Z��a�.kcm����Y����jW����蝣�\8�idbI��K>��iTE�0��D�a)n('�m��1�ŲS��	ˆ�xuT0�X[oMe��ճ�#T�ƍ4%�n�B�0D��+`3M�MA|>퀡�Ô�$��X��o>ѣ ;:�����#���*3I��>���M�IV{�DH��)'��gr�է�Q}��=�ړ��E��P��b	�	Q�����>8�}6L/�Pn�t	�s=�-~����V�ա<Aݥ���?����.����RLa�l�DY%*����g�6u��=>S�@�$�Y�k��w����>��{|�-T�:��ٗj�!��E�.�"n���D�X�*av+n9�}�V{0MQ�̼v��T����k��/��fU�6���7d�UR>ݳ��6AVF�#d�z=m�k�q�|N�6�q*�7u��iF}�T�H��'q^{�ܨ�Q��P���zW�Zm�2�k6�:��:s�vE�s��.+m��>%�)�>��g�3䑣��I��c�	U�1��̽��	�vXѺV��y�x
��d��k�,Ʃ`��>�1R�������\��+�~G���,\SM���L0�`�@`�[@ؙXʊps��g��,ğ�ʦS�C�H���|���	�����-�ȸL�g>@Ղ{;2�=p� ��~���u[hS�n�Y�
��\@���@���o��"<�E��m��A�FB{�x{�[�6y�x�����|.�4[l2ZP.��b�7�Y{����ؑD�>y1Q���&�6,��H"��)��a���%��J�J�)5�a}�j�H!��*��fZm����8���i�p;m�?�ۃ�^g���%D���f�ac#Slț@�.v��C�~3���s�U�pׄzɤ�"����a���)9� F�,ɑ'qJ&��t��~���5}�U8h=�+�����ݬ*��㍫���޺�����弅���6�_r �ҽ���7r;C.me��e#%�Ԯ��sc�����[��,|�)%>:K�!}�P��$�{`'�
A�ϑ�5��G��C�n z�2[�QP+����UձQ �`�9�������`��L
�a��	�� )�{m�+�V[���ˑ�ut�w�\d�L�e@�GZ��u$&�W��'io��B�
�m����G
��*|�+T�j1�YQ�)XD�[������D�C{��[�O�By&r�g#v�qE���z�"���:������6�&��^M����x:�\q����� �n(�@�y,���Zt[)+�R�C�O��	�\	PL2�W�������9qsp1Y?t=Vb:��v�gF4�kx=��Y��z3�u��k�U4ך8�Q|��x$�Zf���4y�>��r�M���� �}��2�Ȩ��7� +Xw}�0�b�w����f�K[����4h4�G��2�m���B���*8��}\X�
�� ;`Q��jvCs�Z|Yˈ�c~��`�ȕ��5��8�'��B?
������r�����/��+�j"��J��,D�s)6?��R��;*_'�7B �}j���<j�'�Jt�H�]�[gE�K�v=��l�;��}y�d���q��6����ȭ9r�C��?#Ə���a�|��:о��@0�x`���0v#�@@N������	|�Uki
[�L����j_�ŧ�xN��O� ШOp�3�/�m�ㆉ�Q�}b�~d�h}��b��!�9����q�U�~�N���7��g��!�je�W !��JظwI�Z��X1��^_���cw�P��C�}�x|<�1d�� �(w��-���ƴ�0�IWb�"�ԕCuZ��D�r���,��%��Ӵ�#��]��M3��4�����\`�c�"�Ӥ�4���V�^��I\!�C>�]ԍ�����
��$�k6l�e��ydqb�2�����V��r�۱�:f�\Y�h� �a=ƣ	4�H�ך�[T�Cx
7[����6Йx{
/!����ͪ�X7Tm� ���F����h��VY��[��JI��C���x�N�i%���уA��M�y��<Ky�v����n��(.؇}��I�P��� �u�+�vK}�F��
��W����pA��{|6v�v��Qs��F��	,���'���Ҙ�pp3��g�`}�JZ��VZ���2���E��u�3"�o%D&X�PM۾*B���C��V5��X^s�Qb;uJ��p�\��\M���j��Q��Կ��nZ䋳�ٷ:�Qg�&�Ssx_����oh:��3CE0��kZ�~����S��>Ys>y��llJ�+������w+D���F]�FG�����Nđ�����+�%����܉YN�>��XBC��9{��"y�/u򉝘&��v�m��A�ƒ�Qc�lB�,��Ã�$Ge�6�����.?k�ۈX�ٲ.
����v�Ĭ��;��%x��o��t}��k��h1͛��:MR_]%W��?�
���pHjh��͑Wz4���ઇ��r�)]��U�v��'�5��ޞ;���`?�WD�.����?���~X�mh�LX�nޚ<�l�"K<�����xƇI�*�X�7��S|��Ж��y�NZP��O>�U��S+8�5X��x�]!IǮ3�	�*�i�j'c���x��Y6��-����Et�P?��p/�.˃���,�")?��=O��k�.���z-|��_</����Bi�w�,�v�}�s;����O�vn��v�;��vW�����f~r�s;g�8�ѷ-��U���������������4�˭���s{�3qn[��˭�m(7~n?����m��O�H���p�?��
�j>_��8�\��d��C��-L4�5*��M�y�м�����Gj�V �[A���ဩwP�;@�Ybdϒ��$�{8@�Ċ���r��R;'�9��+s@��&���kr�q�#9@>�}Ro����F�\. ��J 92 ��	 'e9f�3, �I�8���z�||_�A9r2;7ɔ���v��,��@�Ur��#�,�ο����w��D��LL{�Ei���Gi�J�L?9���[JU��{���~@f#�3����^$���6�~��q_���l�af�dizPx���<���Z�aK�����q�?�\@�9�F�+��>0�5ˍD���I�ޫ����U�{?����p��O�z�uk������_�����	�'�"za0R���[��f�$����z���LNj���o(�w�`.��f?���E�yV,�|��g�|��gos�_�0�y���;��3�}v5����_��c���Z�<�#E�]y�J�>�5���M������jι���9��99�.1�^���w�O̿�6h��f�=�A��>2�R�3L��Z�H��Y�	 �M�<�&a���sM��#��:�ׇ&���}7�`m�~@'�����"Qϋ����Z�@� ��,�Q�rF�~b��� z�Q����c����D/�������	�a���xö�n���ذ���m�_�P�����5�+���9!W�Ӽ$G$P��k���)#��"���s|ՌBӧ
����k�9��%t��Y)�oi2+w��q���8�K��1�Y������Lt�����1���:�0jM��Z�w�@%z�)9�H�R&c^������6[���_�Z,�Ԇ���i��Jfr��C�+�rR5]���ڛ�K���?�f"�E�w��r�/�l�W+*��P<�)O4f�2�N�S.��6� GP��'��,=�e<���3��Ӵ+��s/7���5�G�@����z�r�rm*.�� �>�ʮ�d��~���;&�&���@���C���M��hb��r���I��,��n�(}�D���beb��~Ϧ��?������G�����)��K��9�j���3*ѓ�2*5��bDBn�� Sn�OG��H}�50����Z����g�t>���(�֚󼟉�#��6o��#�L��c�To%��H��6�cs=V)%4�XO�=Vq�)m�����I/f7�6i�\��r�[��A��\�B �S�:*�@[�F��Ux�k&xsӃ����$�GPْ\���X�ܻ�ji��y����m�B����B���&�Xr�O�h*9���$B_;�t�:*!�klt�U�+���q�)�Z��]���z�
���4K3��i#���k�>�C-�4'��Vx;��U�u�H���' \(��sc�]oq��-+��!{�{QW(�9�r^�eY�Xo!Z�yAOʐ�g��30%�m���tb����&X�M��c�/
�gL���j���u�/Q:�/Q��7�R��B��l�%a�8|�c-`S��{A[�;FY�����?!�d�/��w�Q� w����������P B���^��
�XHh1��~(�^���<v/�է|��C:�F�vù_���f���7��>����+{�w���A0=��w}<q���y��=����Ҷ�ǁ��y���&�o�����������֦��J���}�����.Lj5|��\�P���˂��s��M�3ۓ��?�kPm��D�U�ӈfz8��̪L��e}M���K:l�S����S�}f�>��QÀ�~�o�^^��p$�w ���2�f�p���0诨Cͩ�as�|�6�׬6g\/���YJ��`�݌���"5k7�E8��>��Խ-�>�Gi�e?��2y�l-wP1�������W��ѣ�Z�<]@��K��y<�/�y̾P`�;� #��b�����~w��m��-������NˑH|��\���X�:"f�й�ӄ�P�8��z�g�a�#��?�)�pߵ
W�̻��UZ�9�

�����"j�M(̝z�`���1*�o�g�ƨ���O��iM�"�*t� �E�z�WM��Q5����� ��gr<4_�_O�j:Pj��P����5�(��4N~@f#�1�p��i^���W���^�ұ<�)2Ǵ��[_��x��W����+P�"��0b�"޾�+�rg�z��ԎO	҈��q@��G�grH�GGUX!�UZ�5�'����9D&3��.T��#���cE�3=?����M-��qx=�ZZ��8�B���ʎ�S#��Ou�D�<�Y�z�?i�������ց;��௥6��st��@��E0�P�|�����xV��b:kz�u��Fw��g�J��Vx���q�X2��dR\2��d�����?^����"e؞�MN��P�r�+&�͌F~���G��~�fcF ��.�S���]�n*ލ��1��d.2'>�!rd!�2��Bˑω�<!� !�`��W�6)K��@�{[��ub	�� ����([�˨��'#B����zB�H>n�;����[�Za��4��@�(�Vl2&�٬NoAnx��Ǥ@fy>�D\$�'Q@*澠Z2ۣ�NB�cB4?�D]�{ɪ��ݰ�N���|��&�23*����ME�%�����XS=ǊO_�|v�˗����A @!g>,�7am}���q����Ӕ�c�	F�տh�;�/��L"IF!����m���6���W��2)�jC� ������?`]�g!�?�ؿ�[W���k��f�H���������X��"V����T,��qF�)+�ǿ�2�Un9���]��N�Yz�f!���P��^18��u���eG�rnU� ���E�=Oh�d`�	��~���3q3ˬ��e?G����Fd�*�:����`3������dʆ��AԽ��M�pwgw_v��vO�c�l���Ǯ�sys�H��=Om�=���BmQ��ؿ}�͡�:�w�;�]2��c-a�I�d/F��q^�3�(}Y	٨�i΁����>���fb���ǃk]bG���ˢ�+9�,������r��,:����C�X��lK���g���d=oŀ��Uy�J��/�U�+�d�����x��sV���."��`�����6]���c�n��gw���D����)|���::�~�����|�����y:\
�TS�	�:ZG"�Z�9ߚ�m&���y*�JG��4�ܤ���Ak�ͳ�;?���V�V�mIG���g��7��Z����I���saLx�d�,X��ʜm��[���L�T���"����ʇ������ݖg�fW�g�!����y�/HBOB�-s+"���R�y��ӊ��z5P� ����{�x\ /�z5�~���A�LH�G/%I��;W|�$�1���k:E��Ts f6#N������Ӧ�)����ۮ��<�d�fxФ=��]Oz��+�"�b\<�O��t�{��=����3��2%����[Ĥ~�Ń©�n"���gQ�{1�[��`���8fKtd�_VN�k�朼�{}t�P�y���A�s��vt��ѱ���1"K���H��눠�Oٸ�m6�}�������O��}h'3:q$C��g1�d��(�\��P�Ltp9�`�$
�>E�溉^�A�+;b��J�ό�NO.�I������^���C��C��/�΢'��v�#.���F��l���H�28=�|��q��<e�H,���t�
w:~��-�/H2�>�h�" �cXÊ�ְ"�5��}���H��D�˰"�	}yT^��
��"�dq'�.��1��N@��]U\����-�w1��;qܕجkHk���(�h��^�`�#�=��l�����hRQ' �eu�H�c��E��}��1;��z��q�.�0��*Ԃ����8G�\��2��ծFb�h���{�b�(��nId��JJl����Q@��y�#�PA�,�zQD�p���`�B�뀅|���\��yN9��&����˸/�r���
mU�[`Z(���y<Ǖ��D^������V\&��S���;��*�7��X��	��1umgh/����5�kwM��h���,��m�J���x�.a�;���uYVqYVq�kRt=��<�@�E��؋7+���I�v�ϣ�0���1�b͕�i0�Ѱ�_���¾Wr���m��]1Ħ������VԹG{�JL=3��I(DF�q��YJ�W{��G_���_/`)$zd���3�"8��=�Ji�:r���҈�:`'dV����M]!bC�:w�%�L)���j]���Q�w�nt��7y�%D�P#�'p�8/�������O��`��Z|�02��c%$�t�fJ#��|(�W��"*��1�8
��Q�&�S ��	�I�C��;c�i:����Po��>F�
]� ]b<r������ �[���K��W�d�v�G�y(�f4��3Mx�qn�<N�9�q��	6e��;v#d<ݑ��"��^"�UY'jaGJ
�l��N)hzn�H����
jk%��`�goW�%�f�iL=zD�'}���<G�y�c���y|�#h�1��ϧy?�V$�y��f�7�Y���<_�f�|cFt���k�c���kx�G���)d'A,�����,�}	�ˏו.�Q��.0֑y�!�M����4*�
��/�y��,d��Q����P?��cm1��G��LEuJ*W�n��0��K<�kYv{�W�u�p��$DB�b�Kʣd�b�c�K;tj�-1eM>���Q��q��O4f�G���4���k��:�4AϽ������X���E����-���`T�k0�M=y
�-?��0�y�)�W��g4���_�ʔ��b�?Ofϐ����������"�"����pߋ�_�_r��:��< F��g��b�\���q��2�h/�2�3�d]��a/�V\��%�"����g���n-�#�?搫���t���g%��1u��cc"į���x*��j0vw��)Z�,yį�X��I� S��~"1~*������W��������V�lO}ފg��6�*yG��9�rM�YgJ˳���"L�T���5Ɓ����q��8�w�qo%��8~e1��!rt�"�%H��1��W�c��
�#"����
�p��n^����h4��"���"��q���&jj ��,G`�d�.L��*��vT^��=v��.�4�F�?���PN,��
��#�����:��E���g�P�U��s�������"���9� ��%!�5{�&��2��w�!���8f1�3���gV'� � �;�B�Wum
Wd�H���c�c|�j��vq��@Iu����8O<��,�h�����!�?o��hs+�Is�v��-e#fn#H�m����!m��P?�D�v����h�)��FZ,@��5g�uh<��D�R�]��)�*̓労·1��@������9:3�yB~ٛ����;6�.�X�X����<�;�o�=f���o⿙��p���;�����8�M�{]�Ll#�]�>d���tu�"quz�mЯN_��RtG����&܏&^���E�J�䌻J�jt�zgt1�\�"�r���
 k�Pn%��%��>��Q�t,�?�S�R-�\�W�BH��}�,
���;��|[Z�9�oK�a�Ɓ�ɽE]��T����r���fM���ns�9�")Az��#�a79���H#)�2t��s3���������˘�) ��\����	>���~O�d%���u�&��뾊��Rd�9e�C�qp&���i��h&|ZIj����6��D�>ئ�G���sx��I-��9o\P���ґ�}�R>�V����Dȹ���fY9�UA���n&Aj*���)�9&�}��ܻ�:�w�>����+����/��5���"UR���0�}Fl�Ї��c��w����m�ϻ��'�H��o���|u�d�clr����Na�Rk?;�9o_Y�a �%@E�Z3G�3�Рt��7��jH�"SUVKSwVr��J��bu]y�i��j�5IӢ[%$<e-W���-d�-�U��5#Z��Ƶ���F#��� ;��'�7@�:!�'����Vj�k��y�C��+\=CO��2��TJw�T�i���|��ц���11w!�m�����Q��;���.��V��ӽ�.#��{�6��b�J�|�$Ui�g����K>�=E�,��Y���BX�j�^@[���r>���l��[= 8��AP$e`�5��}��kg�5cYq�'���z>VC�`7�7���T�>Bs��>���ez����n��)��̯������RB����H#c֏���
+lPA���7�	�S�]ѯ��Pka�,�~XNj����B���b��?E21o�	�%͝�zp F����M���`�W���y���b�G���P�iU�H��%�����ϰI�{ݓ�&]�c#A�#goW_e��J��s� �1�R�g�$ |
A^ծ��2M�a�ޙ���y�����6S'RX�`p�g���I���nфYi=:����ԑ3p���J�zc�Z����sZzw?��y����;@8��ɮ�;���_��}�M��^�ɟ�����M��I���9��������Npy�(_��LjBb���4���L�����:�2V��'���(iD�q��'�v����7.G�Nv����2t��Rn���(�(���cҒ�`E���|��`eѸ�%u��F�Y�@75^Wql:h�7�Q��G �<@��p �1�]If6ͯH�b�,�x$呤�P/�f�u)HC`Rƣ�x����A������)v�A���rO�Y�u���"�$�����JA�El�]�e��4��+G��y�qd���c��y�82�G&���G&�i���ϱ%M�s|i���ϐܑ\��T��Rki
J�n}-�Z���I)��\��I���bS)�X�r)ڠA���I�:�Dh
?t ����z�PO~/P�f���I|�_6�k�Ud�1.Oxr�O��ta�G�Zx�ǦL�
kG�s/7�4];`���dk��kEeD���!��3Ya��:&XWO��m���ۨ=x�FA���pr��%��E�9W[|�y86?L1ٟ~S�.'���$���Ȣs蘬��t�#<����m p*4��:|�Ymx:���7Z�Z�G����/�Z8;9��_�(����,��%����h3ٲͭX�����'ͺ�'��e;�=��}�����W��G	w��gi�d�����`C��K�=��e�(�ѫ=IqS f��5۟��Py�b��d`�ou|4�\��N��^s|���ڂ��Ѥ���IfmAW	GZ�[.ʴq�,�m�۫�И�}7���`��kEY�6+Tl=e$N���y3H�����/�m��be�Ś��ٚ�k���唡�>�b<����:>�Ij�H����b��臋qIS�Gs�� h]du�G��f1�m��_��8��e8�>h����}çl���Z�����$���"�%�<���4?������4�@�0O�;�N$d_Qno|��u�� %J���b���V�e��*'��xj����m�����*<���!|��G�H��#���G��+r��J:�(wNU^�A�~@���O�o5���k��G%��_��]�{�ys�?fp��u���ߡ��+��/��!x�m��be9���]�-%F�+��_�i�.��� �������S�Ab����QB��Q�?���3�r��6�L�uo�G(��O0B�ৌ2s�>r�Z�4j�#Z0x+�L<ƙ����j�_U���'����S��DFhnN�'�FO�=�h�$�ѓ4�������-�J����\�b5ҏ�Wj%�z�,���|��7�Llל7�M� 8�_���V
�:��zZH���
��D����Hi7��Hʇmt�MN5B�SE��H���-�O�9Ӕ<��g�l}�������y�kX;�V.��8��q�S`~Ff��2e�8$���+(C:
�	o�5�~����mk'2X��RQ�C�t���)i�Q_�K��[Ύ�qS�N�)�����=���K�����A���DpXvy��(��ET"��v7o��ş!8S"%?��r)�y�7k��op�N��=<���}:8@�ܗ膎��项��T����q�r�v��]�/��>=u���#��4Mr����D����il�2s�N�s���q]�V	ڇ��0R/;�mwn�N}%I��:
�q�U�L\o��g�=]�/�Z�v�XBԵ��,q�j��7Q���,�0#��G�M2J�ޠ%�Dq���M���冉HB���M������#l'.ɘ�I�<�?�^��D�1�m��/�0()�5�b���a�헐�x�I�4�"��3����(]�&�x��Ɨ��0�.\�xFf�OC�^�K<ci3R"��F�B���q��Wl����G��)R˧�b`���j�@��1���hax1�R�AS`JY`67��$����r8��
Y$����5ҷ��T��7��qz�7'�Y<^���&�G̀]r��]�
�^?���e�aǅ�'&����r���4���"a��K�e_��`t.�q�6]�k�ݲ�eM�Bh[�L�Z���ļ+}l�HGCՊJD�b��bzQ,^<��ب�$�F�{����#�_�0�_�K@�<jh'��h��n�O�Nu���9�Ɗf ����^`5��`/��*ډlIrxU���vb���<[E�j�c�?���W��B���I�= ۥ�q�{)�c��j9�ô���a�uK;,h���?�3<?Ͼ�����!��T�J4�����ݥ�T^�M帠f����b�ۜ[��X�����H�\�ӯ���΄�P3 �W�����m|�d ,��k�i�!���%rs�$X�YV~��ܩ��#7|z�)�@[���� vJ8�SVF[���C%��H�������6�ӽ64T*�%�O����G�X7�ؙX{��)�bަ��f�<��4�!R���J0&C�@U�ꍒ��ɛ�]����-@��n�8F�\Xܝ��`h³���~6>������758sHk8Jk�G&��G��������y�uI~v�K���$� ��4�᭨{�#8��\g��{+Lؼl Jw"C�`E�*��С���0)��5B*0
��x�{l��%9�*��m���6xq�X�a����Ɔ���J�э{�e9����]��9P� �)��k΍ԣ���M��&my� �°<�b_���Ҹ���X?댔�y�en�.�il��B�	��(�<���`�b�l�u�&I������m46�����Ӝ�8l�����0{��(X
�q�9Z�ۦ9�l����������v���O���� ��I`��&�5�+etk��ӹ.�%b�~gnd)O����Z5y�:�����H�Kr+��`��5��9o[��7�/�سl^o�%�׷�Z
?�ȡ��Do�	ޥ-�5���J�-��]U=�R��v��\���N�Q<፧rrW��(G��g��݌�_Ť�P�#M�K��nW��$`�":�0 8 ��|߾��z�6�_orW
����3�����y@E~OZ�t���c'�Ooz��lX]ygs��/���qܓ*�,
�mp��+G�j�_n=b��Дo���9N*��FP$�2�%&�)��Qg��o����a��B�S�w�����2�/��������R�O��s��<�_���2e@�?1���4�-�ԴR��MM;�W�|b9
��y��M'M;��f��֙���0���i�hȷ�Rn�k��m�Ѧ�p09v�JY�H^�]�m�Lm#Y�cˈ�-(3[J�H�xkhc֌�Nj�϶[��x9w@ט [�w`"�؎m&�$XZ��|� �*��oU��DI���*T
����Z���)�%����U�7%�*6�3K��d�WB��`3�uɎ�vȓ:�?G+����q��A੅J��W=#	[1�U�n&���&���&����,5��ԣ���=�<�ڌ�v��(-y����)�b����c|dWwO��7�Jp/�#@��Kh���W��(��VQ���^S}c��Tw�51���k5өf{t����I9�F]GAI�݇��C<��M�C�x�.�-^�%a�g���,,!�P�x�/�p��x���{��ՅW��<���ל�@#�b���obf�&���^*��Xh�������#���q;��\�4G8�o?cM�M��J�,���ر ;����ZhE�a����g�#篎J���'t�����Q9	��lwǂIJ��g鞗`�|��G�m�-����c����M/���^
 K�M�I����|�Z��u�~ql>&$2U8+�^G�ƾ@��~ӽ��𚄋c˰��`:�8v��8�x���큵���Qy+]�,eo>w�{�����jԯ� %�g����%7Xy3�U�s�WQ�R-�.�X;>�I-ݱP�O��x+�@-��##��v�9�/����Y���m9�����+��OY�W=̀�-5�xَ��ĸ`DO��#��jZ�VXuȏW���젣2JJ�]�Z��5�1���3���Ah�M��\���Q�D���,���S��	�����j�\�WM�_�9�b�,�oף�����z�G���� }Kĵ�b����H��$���U�&�����Er��P:r2dK^�9oǾ�j{=���Jr�.8�,5:����x�]�mg=Ig��M�G�©�Y��})�G���^b{���ph1����dˎ����pku��Q,�9��A8��h���,�4�Ԟ�i?�MX�^���(��2ox�Oŀ9�������:����B�2s��eh�� 3E�x�Ms������lˡ`��ܴ��ڊ��<_;$� �@�v����~Sϝ�/��0��j2���P�)�u��ev�@��[R�}�v6��S��2{�RIJ����ą\'�'�����.�������/�Ki^�����7�l��b�{���� }࣑-�(X��[%��O�&��(�	�U?�k�s�~�A;��յBx� �O�>�rG=�"�[`�Se�MmJ�����Y]�y��h��`
U�LO@�V�4�~�P8T>�칼�,Q��z!�ޛC��U�sծ�m�k�|~���2��h%�+A�`�x[1k��I��.ԏNJG�T���b�78:�/�}S��}��u��qI�[㭏�M�����}�����k\�~�z�(�x�rng���RsNX@cE���q����������xm.�O��OJC���9O@%��%� pM���c�֫cf�������#i�
+�>�Q�>3^�;�Ų�f�=�н�ñ���r�p�M�V5�J�-��L]��~<�6f�o�ڲfĄ�WaS4���ҫi�z]m�st�o��>�e=e�$Nv�9����qT��"����P҅dV�9[1��:��R�o�t�k;=J[��b	N��pϽ���U����'�f3��|������y>3�;N`yH�>I&������O]}�C%0j��-ⶋ���	��8'E�/��%������B\�ئ��G�	O�4g򓄸5g�'`�U�B#�<�!�1cs��q4ۧ���n��m���0�N�:���e��|��7��@Η+��>4��"{�A�.cc�G��1�1mI��>uƼ+C1��X�cc�T%�bp�ؑw�ю\�wO�����q�>�,\ ���ǉ��4��y�P0I�<ƻ��:пo�>:K��~3�l>5X�A�h=����(����� ߟ�9�5��.8���/��Y��7Y_�g� f��UG�[Ƴ��tH뮤9���j�h�J��|=�1D%����J���ф�)QO�a��s��}��Rl�+�z6.���-�hk=Ϝ�[M�-��"�,$�9���fУ1(-�y0!>���˩=
�_\A��
>i3<���J�"�A������{�����Yb��,a�9e�g�9�����!�Y~�1��B�v�s��pΖô|��pSZ��M���8Ή#̙�O�8���s��8ga�OpN�"��EV8g�f�sΗ�}c�pΎ�s�*8Ιܙ6��ι�dc�S5�`��1M���Ў�����ю���qΥ�qNiD�9ζ�9yw�1��,�G��n��!�Y����]�����
9��`ݺ��Uǚk�8�D]�τ��C)�4���+T��ύ�y[4!@�QҔ��%��Z�����.����L���m���Y>�؟�_t�>�[��!�+)M*�,\Ӽ/���o�.t��d+�V���5L?Ւ�����5&�f�w��v�G�t�jzU�d��/.$�����pڽ�P��� ��υ~��íP�Tm����Qߊ�lZZvu���K��o�,�*k�J!N���$��Zu���fxӷ��8���yk�h?��?cy��y:@��d�
�������|��kg�2�,�y�|%?���Ӏ��x~��L[��u�
��fp �c&�"td��U�MG�1/�F������{��b>���B�F�궖ԥC��5s�2�C��,l�#>[V,�ObB����k��G~�
��g�m�ݤ9��U��g�ʯ:p�q�Z�c��i�$�S�.�g��9�M9�[ӎ9.�A{�J�Z���lL@�;�*f��;������E�"}UωO���T��T~�f��̀�fItkS	4ڊ�<�60O�s������.q��3F�x�1�H@Q0qE@��J�/x�"�Okxe:^����=�?1��	�*x9m�{�UTsӜ��񶅀b󻿐���yh�OQ�Q7�z�����a\�5��h�y��j�XKnܡ���P�+ =��q��.�\�a~Unu�y@��Z��^
��o����RG��8:�}~�`��������8�4�j�8�75���AY,&�����WI�^�9�^[�8����sO.B��|l�T$�6Kv?��g8ns��h	o�E`�w�[���Z�����0[o�b���A=������xo�[�Z�h�@��gT䜵�J�T�G���&�^�%�m���K{���1�ED"�VZL����Pe�.��P��I;��lq���)�1u�r
���@��
�]U��i8���\�%3p7=`�f�sCۿZ�����|��lBzׅHGC�au�I�q��ͽ?�V���th8�=�����@Z�Nv��|��w���a5+pPtm�V5/��v���>8�����513�W�#���9['Պ���B�t]QR_�==_N�Hdk��zY�F��}�����/R�s�v����������G8�ٍ��U�j�؍|��(11
v�cDc���O�i�+��x��z�Z���Gqq�Gq�P�q<�OK� �Q��{��D�oSz��bx20J�o!�4�bc�L�3Elӳ��1��|��'���o4��`6��PO�B����P"�i�ZKQ-����j}��q?�k�X�W�s�������ie�qv��v�Z_}�N/�O̲��2 _�Ws[	�ך��?� doלo�#� {���V_#G��G�k�6�W%�7�G�������S ������O��8IJ�I�qN[cKd�-z�D���ϡ�jy*��h!d�(	`.��@�$:�x�Z���漩�&�,�x�a��a+�݌���p�rd�S���І�
@�=���䈂�1� ;�^����.�b�D�.T̉�r�b�H���]�YƓB�������$�n`NW/�%�U^4�����k�o��BG����P�d�{��X	ӆ��g8����r?�.�-��mykE� ���(���؇�4�=؟�������
���B&O �^�	�K�'yE����PƷU����@������_�VӖI�Q�E�"w!E��'�y|:�IH�՜�i\�-��Wq$��w\|#�(ќ[��X[=Ai�9�{�^#���W�"��W��:F����ٳ\D�)3����s�ֿ������(x��,y�\N.�ַq�mE�
E�rU��EK��М�h=0�4q��qV?������Z��ZY*��>���p��Q��vLWO��Tdx�D��>"ǡ�t����	�����ȹqxf��5jV�P0W��a���a�4�c���0�Hk):Tpw92��͔�K2E(1�F���]F7s���>N���*L�,�B���/�o���t#@K�,{+E�(�% Ma)��
J)E�ɒ@T �%QD�y���ʪв�����#
�P�v~��sg����~��J�̜��s��O��p�^H/�S_��s"A����o�`�4�91����&!>�ƽd���=��R|X��#��H�7�a�J��m�8�ZE�m���%(櫏���(�l��t!9�R��� �\D�>A�:�������<y^����E-�[a�t�r3�:`Rk��g<�����x����ٵ����M���ٛ^k��{�kMsj�׊��j�F���s�!P�giNb!���#'՘1Tm�3��2��n)i�ӨR]�7wu�a��nǬ�Kl~l.��I�6�k�$W8*��[	��^��]{�9=~?����&��q+a"����8������^[���9i��R�d$��t��/V1O��667�|W����3D��˔�]�F;�6��%�|w������mT�u�5�8�<� ��M�� �Z�8?����F����b��q��yta��T(&�XgO�S������86T$Um1�[���Em�~�6Ȍ�M��W�T0
�@C�Û���30��\8��@\�{��j��4?k�0bb� #Oǎ-�6�Oa��=x_{���lM/Ϥ@{��+k�$Y���p�
Z��x=�Q�$=��kln�t=�ͅ�z���1�_���W���>����H����@ �z�����.otd�����^{�^{���_kF�;�F�YOO�/�_̬�F߮���~�DC?�Q���i�N���XO�N��R9�*�ɚ�����w'�U�����/��\�t:�>����;��unw�T-R��l6hp&�4��rX��/z	���z�\�N�r�4߼��Mc�m���EZؾ��
-R%Rm}�A��r�h9�u܃�I]�o� 6��8�|m��l��4��q�̵����I��Ocׁ�V1G0H�nL�c{5����$<�Y�4�0`����!p�	�d�`���j�ܴϼ�Q���Ƭ�k���eK>l����5��;����?���;>�(��W �.��N��%-�Gx�`	c��O0/�C��{8W�׽��m���x= ����A/9Ӭ�P�x��k0��� �.e5��؇���x�����-��[e�8�K쮳���᝼E�P̝�c@\�6��$��='*Iq�g3�p7�����v:�O��livu��H��� �Zv�l�gr�HCL������uH�P�T�M�����$��K�K�T� bl$M$�n=�y�S�h�f1]g��2�ܜ�����
e�d@�Ts36{G��G����H�k��Ê�)TX0���'�P!&���w����G��V��_�e�}a����ߖ���O�� 6R�-����4BW@�c$ͷ����a�Y�y�7�w>$_�-;�qԛ�M.�9�Y���\u�E1S�������������ne�hbf=�so���|�p0%�#��0��4���)fg�Q��@~�E�MSGu���)�剄��2^e"�l���;�
�D��l�M�S>�eu�wp>��d�\I�w~J�{�.��~�1�ʶ�ᬋ83�FjYH ���=iq]*7*�T4ggMH�XMEm+�;��6�%:��]%[���Y,�}���G�m	�GS����>����ވ��5�G�c��kY�'��l���N��FQ��=��UR1�2C.x������>3;����t�	�y���V��K�P� #\����B��r�Tt>R=�c�p��@�/:�w��i��#&;�_a��H2r�Y�*���κ4h��7l�ݮR���@�N>������:�m�"Q��8F����!�).�����l�Ѯ{��|���a@���a��h�G�cC��.8@���a5v���LT�q��OCv�/��3�0�����(�)�2<Mg��]�����LSlЅ���uI$	�����SJ��o���A��m��L�U�V9�;�V���JS84��~�0A�Vs��� ��0�[p!��pѲ�T2+,`E����/��;�|������7��gg�Xm�0��Ju��c�zEȦ��0�b&��B{������I��=_�6�K�4�~	�_pb��%����@c����qy�9iZ@��m�؍�]��:m�i�l����u�-2�-m�#fL�
(ťlP��>��n�Ŗ_0�
�V�����{�dPr��!'��L� [��!Kr�i�Ѵ�IZ��Qt��1�T��T4�P��=��ݐ{uR�|R<��b��H56�(�d*JC,�/J�R�lcs��/ϱ�7A���bΜD�K#�'	��EI���
���N�AOv����0Z�Ƣ5<κ_�0L}r�vM�<\ãV���}C����fO�ͮdi)�@%-��������Hr�#9֑��]N��8b������T�w
�c�/�.�2��sh�
�CЛZS��� �B0�|o6��u=�}�� :�q��-��^5vAB>�g�%� u�U���j���)���0�l���	bhD��Lho-B!�G��4�4ي�:S̝'��_r}a��"=�𲀩����-�2tZ`�C{�I�t�ٙǘ�d��6�'{8ߖ���2��1[��H��ׅr�F����p�]:��m�bb�=�0P�6{�6G��eF �]|�����J2Vj�*'] ~Ze���� X%��-�*�bNZ�c��_Ŝ,?U��~J&����Y�������('>҉F��-2V�g ���VJ7�	�t��{3'h����1q�1-E�SF�5�!Ժ;Qt��N=�����7��`}������
��S0_�#��r�N��(&ji���yOѝ��r|�j�	ʏW0`G�Q�A�T�T^U:�l)f��.�xS������r����M�Q�F��T�S���J�tpy,' K:�2�eI���o�#X��������_�a�F���qZ/��]j��M�e����i��^�����R�&˟\݂Q���x�=�o�j�b�f��+�'ı�Z
�,��6Cp�����| �yE���\t߈�6��o�$o�hD,��xv5�Z�Q�z$	W3.Io�ǿŭF)l5�����;Fj`Zώ/�c�(O!T�d���^"�k��<��h�3��KQ64�U�9t�ԻFM1` )�B�<���;4>�����Ln�g��L<�i&�Ldw�Ƚdt��bʌuGJm>���<�}0�޿}��s������&׏䋊ȘH��O9�*��y`�1�`\�����q=��#���� ����F�x\J(�9e����~��������x�}k�y���n�[�n7�a5�;vx���0i�/�v�W��@����T����w̺�d���e%10i�^Q#���N*������d�}��B��w RƦWkC�'"��9�b�l���n2�F ��^����%�E�ԅ ��!��/& )g��!�$H9*�+���#	a��!�ܷ]� �nZ
	t���BZ�Az� �!ۀ��V�	��]m�ֶ&����!P2�^����ׁ�K����� %_�Cᾜ�g��i�oUJ��~���<p�{
co�����to��qfARQT[C�\���{����i8�;߀�=@�$��$=�^� ?�]�Ed�N �BA�� 3B@����A�N �dF(��2Fdd[���'oȜ���@�TA&���v;�r�.�Y*�v�.�������D�:�r�y�
2OY�,^�vd{9�@��,���.W��x���xv��˒A�	�����W�>LEg�_���z�_�W}���a���"Ul�����U��?0���K��5N|�x������i�i5�!����
g���>!8MNg��%8)5�,$8�	΃*����g�>�x}Y'��>��i��I��$�n��"-4��?)(�Xk�s�5���7Oߜ��ti��'����Kp�VἬ�YJp����i�ndh�E ���=����A�:�Eํ����5y��ݤ�r��2��E�[3N�����~|���4F-a��]����������oh��4�G��dঊ����B���J��wo�$�ړ�a ӽ���[{!���~�ޓ6�7:��s@��m����͉�b<tQ�Jd�����͓O>�n��m���q3��^_�PkY�0���<妞 ?�(>��&Q7X�$�K��\��:>����M �@�`0������"�c_�����j6��J�ʏ��8P�3]�!݋��%�ŗ����"
�>�T�BG�d��XFm����0�a_eK;��1<S1�>O®���P�ފYέy���BgQ�����n� g���$t,�2R��y���P����M�pC�%�
��
0����'y}$Ԍ',)�{zzt�y�f������C��i�O�⑶4G�d}s�٪����ּx�՜�  ��{4�I��N+��-�3��Y��ԟ��)�]f�w;�wg�W@ɌT���殘����\u��a��-�g\�g�5wE��o�	�f��.��4�����ɋ�9]��
wͺ5c�x
JJ�54Sɪ�x<��6�F�+������2L��6�e`�wb�^�����x`���5��"�s�p�Ν�8d�vh����L�uuSϨ9�ܘ��������9~\�ϐ�91�l��g$��aw7Q�m�k1:��yD�0���Q��?��;��L��.�_Y��=}��RDb�O�����}#�+c�Ib��ވx,I��C����k1B8�~q���8�#m�<77���*t\3a9pɤ��� �׫��nNʖ⧻k������^]^��
L��r�d���y�AE	(���D)ֳ��ҕ�3�r#�; ��TU�8P����ф1I	�CPv�똈����y�C��5x#�_<6�-F�
,��j���3&^��t��zDފ���$+�� 7r�M�0Y���m ^yI��Z���C��Ck"3����~�7�[ܔNl"��8����D��?G��ֺ��1|�C��U���[x)���7�ix�#@t]j[\�ɟZeoզCA�!V����vi)��ŞX_ד�Bi�u�\��v&�O׭���~�ϗ�g����g�BA��>&l*��UǼs �jx�r�������'y�%B�<�� �9>=��c����iӛ���뭧C�ffܬFf=j�j)Y��u����~#6S@}�xX-�g�m|�	���$LPڀ���W00[���c+æCh����b�����	���9�����I�E���#�S�^g�|kz�[�-����'!�(>2��V��:�(IM�u�&���$�>�۷]�b�ы��a��'�w�
Z��w��X
��~��[�B�����"���b�L�#�Y��ʷy}q�?\��u�f&U�_�XASƢ�8���|�fm��I �nY8}T�z��4p2����4�6�gQ��P�ɾK}���E�[u7eS�ǫ�r��'y&��I&�$�ZlD��贜xZ�b�����|+_XB�z��ÌZ�˳�N��s�������HϺ?z	�t�y4ibs�R���`*��I���b����8�����c�'U�ݷ�ւd�������y��9/�5
�,�5�F5�����s��Z�Gr����U���f�Ԃ�KP7����Q�rHn�n8����`__^�ۃ��ƭ����ܾ<�.Z���"��`�����=Fpy���"R̅���U��S��������E�ki,�^��{)2��ޠ���o������_�:S���um��$y�1(�j�	qz��P#nxt)�n�T�)rY��X���RS�m�^*)I>K[������C|���6>������T���FM�yW3�?��Fb}�/8퍴~�9Z9"4Gq��d��
�c�	�w>S���4�.��[T�^`@�=�ej �)㎻¬t�4 �Gڇ;p0���cFZ�EdxJ����������	�c[:Ư�æ:�yDe���ۼ}�yuԂR^���pu�)�>�����ɡPs���{kp�Ӧ*D3&#�!b!戙�1!�Nl�h�0�����(�ʑ��*�=v8���'ǰ�ɖP6Y�-߰U���� �{MUqO�3���,Ԋ�E�ԅuC4��hZ���+rӊ.����\�պ����N�1��q�z���]�R��#	%o�k��=��'�w����~pP��@�Ϧ���=�ڼe�i`��B��~�w��g�f���>M��n6t�Y�ky�)P6�Vur%��+�7�m� 6��o����/���`L�e3��>RY����]�5o+���e�H�����7�T��.�dʵQ�K�t����[����eS;e�d���`���t�cH���é�ӓT�p��{U��ُm��;᝞�"3/HN:d��(��V��%��.���q,,m�H����wYj�iz?=�&
-ΪV��r�R�/o:��X���Y�x�`oɪ��.of��Sw�׎b4!��D�_�Z3�;������EYu����b�o�7�"���j���Y���3��z�N)�N_�K=�f�Պ�ZV5�ߌupp�{o2�}���[SLϫ167�CM-5�����T&L�q҃4q��.p�bL�,x�R��F�O&?�Y�1��i���@1wg�G�S��ܛ���v����ܣ	���<i��p��ӃIB/P'��� �� c�`�DN�U��LB�Lt@�`܍[٢Q��BݪLմ���f�x#�B�4"�#!W4zƀ��t���G��{1at���?&�� Ŏ�_�W�?ȇ�Q�\S��0��9����D��|~#�q�����P�0�Z@BlO ���o������NB����i0���y��eK>�XJ�(LLa�W��d��U�*��I��"qғ"i�"N�߅W7�.�0�[�AJ����B�ɖ���P�	���2��H5r�~���+�'7�I��:�?�K����[�b�k�j�6S�YkY"��P�/d�'e�n�k=��A�إ��A��>��-�s`�g��߁�;�#_r&#���fo>eU�7]�`�3��r���j[L�h��К��oNCc2nFC=*�\-	��?֫�7�BC�BC����4�-��c��Y�س� �[vk�.�ӣ��Oqz����W-Ԥ������v�D�n�'�����'�������o"5��ҥ�a#k�Ά�����i�j��l�t$f��L+;)7A�.6�]��!}Q٭����j��+�my_������fH[�7I��xB�k*����C�����
����j
-o����C���R���;=�����o� ��RXݨ�|����:���Nν����~���j�6���Q���֏#��G��_u_Օ��e�t��P�}v���4�}\V��^��y�<��w�y0�R�gJk��s�Cb�L�}��Y�����a�.�d�lQ�>	�.��1rj-�׵3�fCu��
�1�+|�[�a��6ԜCp=.��3�Umn�!	�Ѫ�������4L�e�"��Ew���� �wE�>�k�b>n��WA��W5����ԲNyw?Z�´��[:�o���1�Y�S-��G��K��߅��@"�oWa����cEo�X��,�<
k��2X��s:�紼:hNciN���i2	�g	��������l�uG�n4�^6�E~�'c ���
{�Ŷ�÷�-K����}��Wa5�+�y�-��5L�-�9&d-�s��r՚杚�uߖF&���n=Q�,��9ʹv��Nש� V������[�I�*�z��1#C�b�W�rXP�p��_D���B�(דgķA�dLsf%�i�n�G�� /��N
2���\�oX��1���'���_��=vN���s��[@b�
���Av�<�u��n]OE�8}���v�����u�6h�J�,�,;� [չ?a��O-[ջ$U�Az9^|.6���5�b�[����y���Rv���Q�$\�e��=��x_I�ۆ���5��J��+����N�B4`�'�*����3�N�~1�.�1��1���"�:qւL]ܤC����Vj?Z{�TҏF]�F[k2��C\����e:�|C�u�U���n�{&Q��=���Y*I�h��_b���_��}l�d��c�S�畈(V
���F�+x��缮�!/	 �-g�\��m<�Ch����!����)��0d��C������uB�·8��#��}N3|
�ZE�z�!�?,�!�i�HQ3���H��ͧ>஬(���x=�Rܶ�����yx��ϩ��	9�G���	*�>wx3s������i^�������&�D��]�����3��x����@0z�����
�9����DW�4�3Jӂ�l�,LA ]s�=0E*���fJ ]#��@ӊ�t�L	j�H�[��;�
.�`]���t`(j�S@�5�vT�ak�����l��'�Zy�,�t�(�m�`�)o�{sl�@Tʫ��������.��ؓ�T���]�ڕ�o*�S�T��+�j���;ކ~��f�8? }G���NA=O��^���g�a!Bi{I�����u�GS�3��V�
af>)f��x��̮�5���*f3�*<���6`g�%���N8s�Ra���Ao�o^�پz���x��!��7k)�.�ߦ��Rt���ઞ@<�1��&�m�1ג�D��D&��6�����vW�ҙ�um�L/QS���˞������o��Ax뿀��.�/V+��I���~<"�!�qHe�!;}&��?گ��=*PL���@ܘwt,���E�[��F�tj�4�wS���J@��w�0����>Ѣe�̉V)��`�z�b����er}���9�>C�M�g��Y �M���YA<?d5��m��s[��H�xUF�Ö��\ƻWB������~�Z�g|_�l�Ծ�9􎋿��s��{�i1n�n�����d7�_��&P�~a�����E�-�i���Z(X�<'���3ގ-���o��2̡����n�*�|�+�dk�C�7}�Hj%�R��8��%��v<0�ZѪ佫�yL�3>��{�R-�k�i��D4K�/.�q�eqX���j���d��$���϶����jVz~��;��)R&�<*��
���ߓ__�`�m)6i����$= -�V��D�;�A�gd�g=\X��Ot��/~�;��O�?�>��0|C ��ʒ�Fؽ#�v)"�M9�Տ��O��6��v�n�������H�4 Q�&�YN���~�oï��m�)� �=�IS�9, �E"���E�/�H5.��s�>�M���#��v�E�1��	�L-ς��j~CM܎�9�"���ȇ��C���f�j�A|�¦�%�e|�&�fY�2��C�.�3����򥻠��A�u�n��2^O%1�! 3[MY_y�a9�a�������(S�ʝ�j�8H��t�N1����Ũ�'�۬L�jc�xr�������6n�������v���@�"�X��Ry�j��P/SնC\�#$v`�M� �jL�_��:	2�@)>c�`-�0��-x�32pcs���Tf �&�p[�gUc_*>IDڕk�r����:�O@��2���/C*����y�	S��M����-p2��>�dW���˷n#��,9���?��GB�b�)�{pX6�W,�Ph-���v?�P#{7��YX�{c��]�|�叵aN�A&Y?y#a�mA�$���;�ÑQ��X2��&��?�{%�25yNM.�����9�ܟɻ��px��!�]�X�]�}X��OS��}�K�M-��>��XG"�a��3Eh�'�0]� M7�%x����8�{%������$�Q3��vu��$��u�4���5HM=͚����sP��ښAj*�L6��ԥ�&�P!-�@$gD��i]�B���d�N�����9���Y��c8��ln�O�.g
�l=o| ��ޱ��\���(����a��L�"ŝ21gu`����<g�nA�x�Zq�ƍW+�ʫ���\����~���2؋�z)+UI�&&LN�Hx?��{'����o�����<�!�P��w�������m�=��њ��\8���>�웝xס]_�~Av}(������E��b�h���@���5�O>;�F��٫��a�(�#ENZ�>Y��	��;�ػ�Ƙ'�Ɏn�.��T+V�o����t݅���}�����~An�ާH䏀
�?��|��9��?%�/4
�tv%����F��h#��}h]x���F�֖+%�C�_�F��3����N1eI?�8�6Q��}�x#��b�݂�W��g��j���-��y�;�0^������ �]oC;�W��{���٦*С�����.-&m`;\UK��2N�z�`s(���ێߢL#�>�L�hOa��!ٳ[Ql�7c�JŜގ�L\�3�S����,�*�����8���T�è
XT:�˷�Į�6�ҩ؞����Ի���铷���	��?�-1ut���A����L���Yp{���3:z��-��_����o*�Qe� #UA/�G��;������o�%��n��=Tι��D4M"Rji1�N�V�ڥYވ�\P)l�XW��_��b��i_s6 �.��K��1�e��;(ڱA��K���:��W�X�޳�b�vm��6v弘�-��ս�A���Cx(��:��v��l2��F�)/�A	-���A� :(3pFV�HFfU�vf�)]~*���_��죥�(o#���q/I蟾��Xk���?�ĕ��wtQ����c�ނ��x����^�)Д��骳��?"Kz�ډF)#0���N&�ä�S�GM|d��2���&�a������+�4���>��E�����~�@�T9!(9M1��[]�u�-�"��j�p���d+��Ksx��=����ְC�� ��+v�B>jm�x�40�-�{<҆�L���Vo�V=�f�a{�[8t_��KiW 11!C�(g��o[L���m�}��j;��սOq���^��B*ͺ,@��!#� 2B�4D�{´[5E����o�1,��s�ƚ>W7L�Ʃo"6� 6�ݪ�V2l�Ȗ�p8�F6��:�X�d7̓qx#�M�;�w#vA�����Q�F�
mR��g���3�]��P|���G� �(���,l)z����4� ���O�讌0�����:�v'�!5U:_k��¤���U���w@�c��[�hw�kx�U��h�=������$yO"W�%�}cʵ�4���𞜷��Q}G�~�V̵��M��+��w�Ju�b��s�����Q�3Y��
�4u���?��,,�ϸx~�A�����Ǜ0>����P@��ˑ jě�@�Ҹ�?�B!�B구�k���w�6���?�w����3�B�Q\P�c*r�|�a��LF4J(ԣ�E�`'��C+�NQ�I����#v�����jE�hI�p߈�*{�hN='G��o�� �0�p�q�{���J�b�����_�k]���M�9��4�N�����h��!��k|k���ʋ�����׳�]BT6�x9{(�2��^�/u_�5Y�8T_��A����9�l��Ux����C��¡Nmݭ\���̀Y S0�pv7�~ی��f|�P�-x� �p��p��� 'J; ��!\��΋Ǧ���
�NS1������8�A�+�y���J�%n��۔����
�~��qɩd����#���4���D&;l@�Z��U	��;D��gp�P����3B�Y�k0�`�|#9*>�Xc�h�;��ф�rN�j%}�ϰ�n)S�->���� �2�T�u� 5��&0�O�M��kl�_�	|�+�����.�v"H���Lר�3Q�N�8T�� ܈"<�Kv+��L��j��6��<�F�qG��4�ƣw����$�4L����p��8�6c�����B0'���\�.�m�U+h/��AE�<�:PH��t����Y�P�8j?�V�e�AL�6���`��~����:`l��oi��{4���HNL�XM��#t�冄j�5rmU.�2N�!��>���U�A:��Y�p�5����!y����%�,�}��7�蚩h ��㪩j�ḓ�C5�Di�eA3ē-�xT#L#]֪iHf�I����7t(�qyf��g��-��B����[҈R�<��ChX��$����agBׯ��F@�\ӂ�1�<	Cx���@{�:k#w������5�����3��g7��6:���5�]i�y���u� �m^��!&������G*����Mw���|�vB���fZw �?�Z(-�Sz$��.�	�;ժ�h�
�"	ҷ(���"#��H,>��}��W�	(]�$��J���z�l��IћsA���l�;r�������u$�IГ,ޠ�3����z��,����Ҡd����
;�ʌ��H6j�3� b�N��w�F��F������\�X��	��ɀ�aS��z��C8wx@�#O3��nS'��|L1�OA`�|�&O_j\��1o*�uK���U��`̧\5�����J'(��J��Uϙ?Rk[c��Y�fbW�_�D��DӢ�k~P�V����_�D�<�B�mF��LE�H�J�F��{�BX�a�il�*����	��$�:@������'O̍��ty����7�y�Q���!�D!�s���۰�}0�;���(�a�����B�еQ�/&1��d���Wc��	H�)���I�i%~�G�w�pj+��N �l$�@�2�(���Id`��Vi$=F��ڇ�4�K�D�� �+�w5=�����.���wo8��e잡r��O����k��zG��ɵK��''8b�g
۬%A^m? ����1f;��3�������LD�3����!�c��Ft�%ls����q�6�yܜ%������:��!:�㞤���32VD>�^S$�)��R�CdN<�"=��}hb�8� o�v�=C��Ϣ��;�G�"�Aa��=�30�~'&��?򞾇E����*l��$�H�t��;�Z���Ϯi;ڶlwNrHaK	<�j耾����Oe\˒�o�Sօ7k<劳{�'ٯ�[��m˰�-��7�X?Ri��k+z)vз�U8c4���!��y���j�x����៽T#w�A�\���˘���>V�*2�_b�kD$�z��U)�1��`��#�^l����ž�������w����8W��xm<z~=
V�Uє&]��mj�M:�>����&͋EB��YJ��ɋ����壢�3�*�cZW=�e����]f���E06"�R1�?r�����j�6��e�\HJ^����?��.������s�۔�!�-��7�#��@e[�Fx1JM4jԀ��^%�Z�_��Tx#?]�֨��"�Q�lM&���t\)w�P�RnJ��Z�;S� �J�EB!�%�"p� �v@��ҷ?o*�P�4l��8�#1G�X���$e��7A�/j�F=�\��ȍ�"s,�Q!����$��a�Z�W����f��Ą-�Ag���Xݬ{��~��d-7��`H�����0�)vZ�B���$L��^�֒�d��$c?��dܓ|~����N�SI\th��&��1�^��z���K����>���>�]� �~9�����bc���r�s��)�d��(����}���y�p�A׵+G1V�Z����8��y�>=�n@k�'�vY��.T��x���i�y� �앫��G�H6�'�L,�y�U�E��޴�Uu{�����5b���^���
:U�^\F��~Կ
/�����?��kpJ���7�O����i�N{��/��[�ח�
�G�S�x�e����67�C�T��F܃�T��[N�gq9����?\N��VM����ҩ���]�y*���a�6��	K⃵����`m�V~c;�:�UMPg֩K �k�
�ar��L� �Ǯƻ�umR�<�'�_�*9�=�������E��R��zz��rC�+"W��鿲����4� �"G-�z'Y����+[�φϔ by�8�%p�nB�2���>�\USc�w���"@n�	�P'Z4�}`��^ �@�C�(^�V,�mfDS�6Q:��#9��=�}�U��_A����\��6�$_l��E�ʗE���\}��:���4�`>R2��	9���Q�o�}L)�./���P3��j&˽Y�r��Z�D���x�p~�@1�F�t�
/�"ejT訉#���2L����z�g�b1��@���r�Qc��X�*�EsdR�#�����Ю݌k�`�����%c^���������û��.��]z\fS�$,?��Zقw1ӥ�M� �v���K��-�_͖N��	�	c�x���j��������i�$Q�o���i5?��-��*I5T�U�Rv�z*w
:9�?Yy��ts�S(fzUf�I]�z��@��C^H�_���b������	M��i��Ӭ�I>��V��&r����3Dٰ��*p��!��V��~ܼߩ���l�)�_�h�`�n���K�Ů��!q��c�7�3Rt�e�g%	�w��BC5{/8sրB�j���o�;���wWC?����k/K�1�������uC}�6������@o��m\�������n_=�� U	4���ӪE�cM�
}I;->�ד����b�<#8�\4��+�Y�n�Sٖ�P`�-5�򋀿��sva��C���D{�ވX,������S�l�y��}���ڎ�n;� �f��f�z�/���G��N-E��+/�-� ������8���*_��i�������+�'���J�����9E�.%�U�+5��d���f[�M��=>J}|�����u#<װ�����"���2���jJ�L*�v�A��::��F���a�]�`Ha����V�3~�`H�;��8�l#�n8��g��D騳a�#��N٨�rC~�a��ʇ��N�'��o�S��۾e���e|=ë���R0kP4�R�+��L=�d��X�^�כj�G��L>�9���Պ�vG���w�~�5��7F\|g�j!'�ƒz���(zr$����9Lk��]��a}v�*�(�Կ�v��yܙ�nč������]����[q[|[��ܯ�l9h89��n( Xv�̳`��DT3���s�����|�_'��:���yb��:���2\��*�{����#��-;|��,g38�M�$�3��0��T��([�7|=���x���z���Y�I�s��F��a�73��?�b�L�ٯ� ��[���Q��X�3��V�׵���h<>�\�-�f����V}3�Z�ճ����&�� ���:3Ȇ2D�6^��l����>�(���Ka�~�Rؙ/���V�ԯ9=�N߬9�F$��=ow�UJm�ʍ>�V�}�
�����qI����Z?��A�����k1��2\��oԵJ��@�C�ƕ�@�;��|�Žس�������c[/-r8�2v��x�36�W�k�
���-J�/ HcUHW�8 �ܶ���/e�1r�s�o?B5�
쀡�0��dO��Eq�즍�K��T��4�	�e^!�ו���܌/��_xP{a�1�`Q'"��D��A,��;���	l�m%��`��,�!�%�AMg�k>a�>{"��T�ݖ�%1^�^c���Ux-5x�/j� ���1���Vh��Cx���^	���
�� �	x= �'^��~���aŕb��*��1��F�Y��^��j�>y��~��An����𗳙b.c���*���_�d{��L���|	��,������kKX�����sa	�+a	��a	%1/B\�i��>��b����'B�mQ:f5-+�g�%�1yV��g#b������C�0�ϋ�gt�w�U�*
��{���lQ����W��W��W+��y����sA*[p�7���ʺX �$���\OC�uH�dq������n�	�T	MC��D��J�i��5� �2C�O _#�/� i �`�b������dD �P�	`6��֮��)�%��g����/�l��$�o!�g����J��,����,�b��׷Ƽ�$`��`��oU��-�E�`�����q��=ѠAl���f��͊����?�Z����C�n}��XplԆy�I1?~I��b.������4qO��IS(q)���n/�J�)���o��ȩ�-r�Uu���-�o�E�=��,2��0�QB������l��,'M˶A��rCN]x�NY��;q]�y��7�FP�]9e�q��T��R����z@W�h&N�;d`�-���躃8
��`*c�$��V�8��J?��n��#�]C�ބ��#�b����bS��E�����@�ԿTP՚��;�S}6�
�� �='�@pi]X���.��e���5O|�*P-_[�d�ׄ�	1�Iz�OB�!���Nb:�ģl����wdKM��/���`���8�6E�v�+���j���t����S���ӡ�3�`���U<Xdٕ*,��JM�->3�	C2���h>v ��$!�� �T��*@(#�<7��W�ϒ��eI��?�( �����u�
��T�?��a���L:4�-��ޜCo��p";u�?���j��0��C�EU��+���'���i��
�-��Fg;�p��S�fr�� �s����1��<J7?��R���C�k�eK�ٌT����A�����8�\v ��R1�Xvދq���*���?�=�-��6�X�"��
�6���Ý�)�r��R5m��vwS�?������c�ຏ��k&�Z���v-"]˵�(�i�)��Oϥx��T7�o�E�E�a���*e��Md�r�2+�4\�s�+��WB��~�dt���f7�:��F���F7bx%�(	ކ�����dB�a��[h=��l[����9fڇ�����V�H6��KH.���_�\b�_�g]�T:]�Z��	��
e����������G�ҷ��t�}��N��N�꟫j:���'R۩_Y��X�'��Pa�=d�|��
�9�P�P��,/����310��!`�
�����K��!�|���|hx���&���@o��2~����>'�0��W�WT8k48���;��3�INŗ�c*�]�#���Zg���8S\�XF���yO_�<���+��0�gp�r�L�fX���|�D�\·Eu�C�܇|�K� ���r)�s��őz��
{{��a(ͤ�~���M�U�QP��;1�n�@&`P�F�b���q����}�`c�&Y��t��́����HoZrx���k������Oýe��c�ِ�+��z�O��c���O�Z`U:����
��R�@a�h(Yh�F�إIv�;FR���d���;��x�<��؅d��8  ��Q�=��e�䓯G��7�����[Cƻ̰l6�Itc�q�5�'��3�9v�� ��(�i�q> r�&�[��:��]`Z�Dq�v�+����܏�|�S��#����o�g�B���2�A��@gigz�����DЍ�"|�>��_՞4\�ۏ(Au�se<V�؍�)��~$����_rM|��v��y����nïm@W���>��YC��5:����|��E���-�o�}@��oƯ�ۺ�Gm[!�)�5��As�U�;����g4�^]�*0�um�+NH��n�]@k���	�͏Dps��ڕk�`�U�
.�X1��
�ۚX1����p��0xp�b-[ʒg��l��s�$���Y$��w��km�G��
�
����׵#m{c��{��ys3�~ƾW��ExG������ڑf"�|�m�_}7� ��,�a��v S���(�X��[���>���a�������a�?�4X��1�	[.���$�l�M��-�h���\C�Ǥ��5oK��p��m�� y�TQMْߘ&���/�2E�T�����)N"SL�2���(K���ʔ���c&&d�`r���{²��֥�!Rؐ� ����2ݑ���~�簔9�ɋ0��ò[*sZ��Fg
�����?KTkA�5�������¾uEb���0O�К�L����N�)�:����9;K�F�	�U��F�d6`�B]Xw�� 9��=9����wU��{F��2O�Z��}�r���yo�ػT�|����xW�G�������-���W-~��ۨ��|��O��YyS �Ң9����xT�x��*_ru�B����+�`9G!���2ƣ3H��o�y��+o!���j��E�I�����e��[��J���2�'��+�ib ��w�e��p:����|������y��x6-_8��Y���LH�Z~ƫ���|Y1��G,;�Dő3�0��k��cs42�sx����d�$y�h����"�%��oJ�fA����6�39�q��q�6ϸ&�ў��/h�ӪG[����+��U<sV�Ir�OH����o�.S���؆7/��~e�í��0�&=�����K���K���Y\���}�,�@�$V�y@,�b�/�!�I��T�A��S�\�0b)�&��fk��D��M�1&�c��ƘI֤�N��}~���F��F���ӆ���qͬ4�*b �n�N� �&����b�]ǘz�G�cν���xCo�'��m_�|^�����cq>҈�,i?$�H;��SA�Y�2��	��7���j�_B����I���ي[��e��� d�����}�_)g��Q0;�J�>�މ�]����zdY5oKM#��M#��G���F�H�/�w���iC��ӱq�"?��r@<^���.^�.J��}�����H{�����Z�űM�X��`W�,&X�1��nE\�ℚk��ϰ��U:iÆȘ���J���+��Z	�w�$9D��l�ט���^���7qY-�Mn�)���è֘<��ڋ���8؂��L0��
���l&���\��e�䉄U�Vl���	P��X��0�f���x��?(Ǆq�*���@a�S)�^���F��Y��.�[�d�ޠ ̘����:�s����9�{�Ӏ/IeS�2��awd��dc8_X6�{�}���y^$�6���!ejPrq��S9����U0���1��V�1�s*O~�m�R?���f��V߲gZ� #����2�K��!�΁�z���݌¸別��3�����6�f0/{&�����\�9%���R�t9LM�vO�I������+[S���2�U��c��]����]#���nl�>P�1�$r_9cەWp��u�J�b������r��28/J1o��y9������3UX�S��Zo�$r6D�J���/� GC� e��E`r��7�����]Nε�q�B�[Ţ���,-����i Y�ՊU����qL�gf�	��jyE�0���+���Ä<`�I[�b%��V)`�����X�4=.��lpN6WCo kL��&$���W�2�`��z3p���O/Vi2P�G�Az&l�#� +�Oy�?����
���I��8�B��g2>y��3�(�A��3'�Ժˠ��Esj�r���ϠΣx7�psy�/����y#�]����ї����]��H܎��� ��L+�Q\:�u,"0�L*����춦<\|��Q�m�@��fZu�cǫ�|i3�Z��'��q�
�O�#;�}/�����D��V�*���I�yQW�1S5[��E��V<��\ڃ@d���=+Za'
p�V����Rq�}D�:�E���JV6X�~,^ؔ'�z�F�� U�7)��r1r��H���@����Ե|����~c��K]G.�@�^y��mB�'�u��N1�/Y^܎D���i�v�όC�ޣ���Oَna���B������OW=�Kr��Z��a�QA ��@^ަ��XT����m R:ꮬ[��}��&�aFC�i���b�4�A0�k���JgA`���4��ۏ ���cݏc��)���c�`-w����*ݼ����/p��T���;T�D��ژb�1���E�@�_b�� Ӓ_��t��f��*�75��R���M#�V#
eG�G�3��U|F7�	f3Қ�\>�:���3D\�p���� ��dx��J}�S�'"Q�k�d	�n[��`*�N~�g��r"��H(�9�d4�\y6tE#�z}^G�#U�Ug͹�y)�8v�F�M�'��_@?�C�����*D�./�Ė��P9!	��(@k7��I a-9Y�U٬�o;�61&�W�2@TV%x�܁���u�0LF��*3Ozw����XεX��dA�X:���2�S*:�N�~H� �>��{��oE�A^s?wc�^[�����#��J�t*�i��.b��C�RG�A�.�@e����Lo�b�p��XI5O��`�@�Zve��j�s!��k'�R_8��a����:��f`p�s�P�O�匁��#Q\ �$%������(wz���Q���|"q�m�#F�ė��Z�=��V�k�,��U�q\�&|A��!B�8n{�_<�A�a����z�(�<H�G��5 �9�iM`�E2�s�/RG�Y*�EV�� �!'v���p /3L�E/�fA02y���@��������"�^���d��)3�����g�Vt��+�����s�������,s�.�C1T�Z�_�77�!�SO��W�A>Q��*h3;[���o��t�Z̀�/�oj9A5�9�c̀�Kukl !��&3��0�M���ۗ&hE0"�Iܷ�V;;|
�АI���uA-��@���/�l�5Q�v�F����� ��N��I��{#0���?nf��I�ޡS��`�f
�)<aLR<1a��#s̪ߍp3�Q<�d�!�0�O\�v臖��(��!�<W��zՊ\�]�(ފ`5]�g�}��2��]� �-�3�����ޘ�����_2×z{�8̅*��0�P��7�\�� cڳc]� o�&�����eϓ��D;zbo��9�㐾�&�?KE����	hJ&���{bwUh.Lo��2�N�^C�����*�Cl(}�*c��S�5W���x�R��PV`z�M[y��
66	�I]4�@n��ZQ�1��&�WgB�o�`*�4*�mg
�;/�1�Q��l�����w*P`���FCK�{#*���� n��j��;����{��mk�6�=Ŵ&a��,�����T6>4Ѽ,&\���a6&��=��m�az,�Bˇ��I���1��G~��L���gB�\T�0��|9
�/�R;�Tb�wٿ$Z�0\�@u�2���ى4��/�5fVӻ+��q�n#���1܄MR9��$4�ɡؼ�Z=�oN/�m�C��c<>3W��%�]����+��A�N�"'����K)-W]���S�:;w�k�oE$Ԣ&x�^������g��X�|�. �,F�۝?3�ä��]�\�&���k���P��g�������蹀� ��-DU�!�c9X���^�ssxܽ�nM��.�:���@v9�A8�=�N�������{^
Jء�b0��sv)��؉���������z�'�}�6��x�s��j����kw����%f_�y�9�cD�1����%N���	���(��c����"����l��c�[ 8$����CKeL~���FP�*��V�[:MB�d���0as,^�uǄx���jߴ�?�D�v�@�U�z�?���!?"%<�㦾���X��7�y�2� "�.+�q;4!a�&$�$����� ��0�g��16����,8���dK�C�{��F��z�K�Sg�����cO?Q�'��a�$��rS�"�ɿa	g�+5F����Q���07�=�Wg�ue�JV�}O#��O+�E��`�G��ÿ���4�`ib1�]���&�qoŰYշ`���k�SW�f-�)VIwH�7��oM �O`N`,�1�ҌJL�b.�s����\:�)�mݳ�@�/=��8��Dw��IeO���9��QZ��B(��M��r�B�&�s*�,F�y>��������8��6�����4(��E�$vO�A��vGp�p;jp�܏�'��z�����d��(�f�^p���wYFvs���EM��{�G[UD�2we*���zA\6Z*����OƧ�	(J���ϬV��٥~���J�Jk|%��.��l����� 8H����k��'�S�O��6�G`���b�� ���'8C���Z�����ȃ�J�h_>�j���b�Jy�Wf�qb���n�a�!��X]E�e�r M��	�gK�t�!ͱI�S��CӚ{�{X�saXK��hk�!1|h���g�����	��)��Y`�vm����6� '�T�gz����h%��.�C�q�����	N��������?&@���R�0�8Q������t��vڥ}��);��6��N��!�˷;�j��g��avN굀>Aθ�R��<� T8�ݓ� ��#v�
������y�������UUE��R'�V�
�s}P�����	:7�QM�I�JN�gv�{vK�9�=;Q���/�e���"��<���|x<��I��k*G���뼿�8_<�%혞�A���Uj��r��A����)~����7�$����ׄ��]���3�Im�����f8��s�Ṵ�����A�H���w	؏�f��j�EJ�wy����I�H��%?��w.7���м�"`���;t��9�قo�q�n�C	�u�%
h|�Ѡ�/0:1��-H��w&���B���cx�+��+�Iלt[bO���83l�>9r�,9-�uWN[��y~�)�q��z�p$�p�#ITw�����Ȱ?^:�9Ǐ�C�{�|����D`���������>�/p��{Α��M'=��B:�$>���W@�?0�,����V�i7��=>B�y�0@S��UBp�\��8��ad�S�_H;�}h݋!�	�x,���'*��uyy�w�J1}���C%��t[;�29�jن]�~{'�B)�QE&�S��&��e�7B�e�Ѻ	͌��'e[�8�X=�<�#<���Ҷ����5�Ȱ��ʊ�)�N��*2�vgS� �Yì�$�t���u_� _N�����(��L~H� b�Ԅ���2�z�b 4�?8�u�u������;L�zsn����6�5O~��B��,�eߜ��yu��l��l�	��s�l���g^U���!�����Զe����u�F�oe�5�������`��W��ٺ6X�s��Q�k|�3��T�Z�o�߬56x�q��Z���!������v�8Y��vof��3��=d��g�d�3t*��J�z� �F>�	n����`��m)U���&�إJ�b�>�F}ۿ��ߺ�恖Z /�38�ՌCh�]�*m$�΃�b�V�s@^������X���z�Mk���f�O�ϒ����aw�v���3�1������L�9��*�.���J���/<Ԯ��fW�K�b��9%�4����~?V��̫��&򁚉
���4Zr~�-D�t��[��=�BL�/]e����5�V���9a]�j"��0�0�����́�R�� ���g"O�ZE&�����\J�5��I�6)+n�1�̹����@�T�Ŋ�.�$kv䄙(6�YÎ̽�U)jʝ���إ�trԻ�h�̈́���s�J��\�YX����R��K]0�+�̵�j�b��I;Z�{�Z0ֵ�_?Ӣ���v�;�?�P�2A�[�ݗ��_}��+ $k�FnQT@�p���
��,���u��	d���ƥc����FQj�@�cQ7n���?��.ʢ��{Y9*(��jh��$V����.�*�X��캻��fZ�F����=��"�����
<$���e�5:�A�R�����	��}�����������{�kf��暹瞙��sx�m�2�޷G�AӃA�C������z�t��mm��'zㅗ�t�$Z;�=�Bo����1�����ij�},�lZ�X�^ԡ�]�#W���ljMsXg��u65UD�l�bV:!D�v@R�] 5�^�t:�~-���؛>�<}Z��n1���5[W���%W���Ŝ��ҵ�t��y�&M�a\;��L��N���N1)�BK�s����qe���:�E��+M�}|��G�{�$&�.��j��zA����D��w����N�}e�_�&��?\S��mN���0�s����V��/Y̖Оqg�D�T��-�8#�'����~IvSz��G*���Z��{��߳�sq�}h�����������[~�)6"�m*�)&��E#������)�d}M���1���V`�QͰ)<f��3}�=�#�J����M�f�M�������C���v=���2���k6:׬Y�Z��g�k���Z;��Y۸L,�^FǷm�^��΁N�'E�&,�7;P[z��Ȫ��9���k�ժ�������S�;��i���c�?����h1�6���*��>�����y����n�Ƙv���g���y2:/���1ʊ��e�~�Wb���۞,�3��c�}�Hn�u���7]��΁5���9�,���,�3�xe��脾��F2֞����Id����I�$z�Et\	�[#\�{�^`�Y�i���D���w�qΒ^K󟂺5���^~�DO֘(fH#����K�]I^���/77��5N/*o7z�||���5m����L'̋��D1:(���pVDs��
E�ky�0��i����=�WJM��>)ľS{}�vx�55G[:"§( R�X}K�Xc�W�W��z�ЋMJ�6�	�f������N3�e� y�D���@?N2�����I����!�/b�>}})��pwN�Fir�}0ޝI�MbYB.�Jд��u}�����j���Q'�5x��0?Z���ө~n�I��5-l���&�c�t��-O�DOT��6��f�.�)�v�W�լ�@��<��,��nC�m�?�n�����m�tZ,u��9�a_���M�﭂��� �i�����c.7;�q����Ʀ[I~'����Q�MW:V�x��x�ud.���'+��w%��dQ���ρ>�/��,QQS��|�7rV{���%p�}���'zG޴�QbN2^�)I�$o���n�U}#&������"C��
�UYG�%�vFF\������UW����c=�d'Ǻ�k�6��^3J���n-��|��y�� ��m®����;zSXCq���������\+�&��AtoT�{cz�;)���f�,j��A<=~F x-�W#���:#Z8#]���q�dao�������ǝ+���)���f�'Gs�K��hn}�XD,z�W����HK���q��n��
Z֩\.&����x�̚L���Gax���N�5����%�)��WyG)�}�m�싖k�C0��]k����ėict�'}�4/[�\�Q����xΛ�ؼ�fz{ǋ��N���;��n�V��_t�d��^�sб}U�C]�*:~��[�}��S��ay~t@��4ZJ]`��ӕ����7�
�1vm�0m�厅笃�SBi�\p���|��9"�V��PŎ. ��QJ�m66�|��\U6���3w�^���ٮE��V�׆���X�Pҡ�O�i���w�����E���h1��|Ww}?�9�۵����=�WК҂���v���_<�WT�S3�#������i��H��J�)_�@G��}O�H a������b5��'�>�o:��?�E5ŏ�X��cn{,��>�Ҳ�%��>8j���ΙW�����.ڤ������k/9O�9�����93z�>�u2P��cd��rx���B�˵G9�G�T+^+����l�+��+�,.��mX�u��RIy~�OM���������~��+���}��w��	4��ѵ�E�sAH��D�ݡ���;��<O�6�5��e�%>�x ݹl?%<���/�ІM�Ȱ��o�5��a�9�g����Y�k/>��wTL���
5��i~�^���	T��F�b.�7�L���-+�Ĭ3�H�u>���m� ��9�7�1�M�Z�|�_s��M�?'C˿����㩗 �>�w���+���Vٳ9���*�-_^��m��S����*�Ҷ'�mo���q.�a���{�gq�@f8+��0��&���Ɨ%��9w߈tM�F6�p��܌����ȶ�֠�I徙q��4I����'�F7���1~xL�����C���%�9�g�>bnDmsV�3�����ta���S��6뿬un6������:���w��?�9}���<(X�i���apQ0�,Lp�{Ҁ��[o��@{퀟hk�*���dM��i�j�t�?�{�q,�N�Kq�w�W� �R�T�q�_��=��ދP|��;�^׫�
��7�����y�$����ѱ��6�qb )���H2M���v�1Ȋ��O&kc���/��{irM��%|���ē*�q���J�P�R��X��O~�/��c�J~�����>x�Ǌ�*�.�
���бO�ay��T>�]���-� t���&�֋N�9,�%<�K=���5v�LAӋΙ�j�k��9�k��/�f
V�D3%v�)��G���i��z9�`�W�w��^��^q4���ӻ�Eo�W"�i<��]�����x�Eo�DO��~�I�8\֡�ҹ~�����c����Xct�5���{���x|��}�����8!��F��i�־�|~�R],��Q 4� ���jO�ʒI�u�/ĶC�)R1�7�E��L}ē���	L�ퟧb���	e�vBg��d󀮶�ב|�W�g��F/>�t��54�a?�\^�.�G����ю��k!��K&������E��2gQ�T�*���\E}�N�{�E��g���-eTu�e�<�=�7�M/�M��f�7����w=�����A/�E�y��^�"�r��oˉާ���>��:Z�BOT�#��T^�ӟ�Eu�^���K��x�ԧn�[Ƭ�]�Q���.��TSe�(t ��!���%f�Օ����+�'�]E�q�V|�6�y2�]��E�uP��܀l����i�)�Hו��K\G�C;t�P��D��r�I�����צo}?O�,LT��k���O|bIz���>۶�I=�]�d�O����1_b%65
^�)�Z�����GbԙE�S��G+tt���~�5b;<�1�m�B���#��
<�����OK
ĳ(�d�3�<�qub����t��-K��|��U��=�Eqs�ܥ����OϷ��l�n)�j�e�g�}��I e?��۳��x�?�M��Ǌ��S�>��/��ǎ��ǎlw;R:6Ji�哼t�y#�2�CAa�?E���_豽C���;|�н��;]�;D������b{�5i9����\H͏�K�������9ʳ=(g�)?;�(�$e���8N�Y7�a��s=)��즼�7Q�*)�[�ܴ���*}H6����FYG#�Əh�D������-�C���{=lW��w��=���94nat����	Q�Zexmpi�%��"�黸���]�LM��(I����.�K�I��o��E��2��<xO��xa蘃�_d�(L˷�^��5 ������ܪZL�)��~��EWC�E�^cֶ�~44Ti��Hl,�v}�!��>xf�+N�	'�/����~)�<Y�4���F9�{���9�#�#	�J,O�֖~�֕���טå%�*����t���,?���c9��[�XE�����/������;[m��hڜk���&�b���4��+wP�7��|�]�h����Î��|�%����h%=���:�j����
Y�
��F�����m�ISs��gxo���w?���a�JwQWj���I؏<�}�X���^����
�����,uw_�wvw��;�cN���N���w�r��F"��"����Ӝ`���O��>-	�	Ns�ؓ�p�:���yk�#[�o�xWOg�n�Zo���Cޭu��3��������i�I)��s#���&�_ߡ��N�7~E/˫�UG2�(���©�k�Nc��|��D�?4���ch^�=xcS'�x�$���D��dH��a�'k�ɭ9S� I�����]�?�8�;��ŗ��^],���TC������ j�Ĝ�>��!��'AO9�>������rUS�TM�<M���C�s'�=D�N{��rzo=�gs��p�{���FN/�E�NN�qIo��������^����zqz����͓b��HJ8�7>h)F��C�mx��<�MG�IV6q�n/-M��X��xR��;ns�)�(��'W$��bZ�E��h�pw�y[eq$fǄQ�!��nܘ"!�v�?�(�<���GR����j�=9d��/��ލ>�3�^we�k�\���}�;�Y�;F��r�{-���Ш��+|G�s�[ƼF��z��w&�{?X|�f�'_��B���V�Qg��d���~�1��|��Ð�Fi�I:����,�l��}���(�N�O�Ʒa�NHi+/�\{���)�??�6���&�Xn��$-ا\�"�5��u�ã��'}��������|l8&J�?1�<��c�8�����J������σ�&�ذ !�"'ڏ@�Y$��4`��\��ea�]�P��C!�H0gWt�Hg���@o��C3	~�Q����Q���Jtecb����N[�`���©A//��̷}4l���X���s\�ܫݨE'�Sr7��܅G}o�C:�[���Փl����\d�y�E���D������d�p�#ɾ��w�]�&��M���K��C.����@���}�����R�(��y���5�0;:�|�ivZt�� A�������N��aƄ����߻Ŀ�s�6K�s��v'zB[����	g6����m�M�s??/�������0���9����We��lb���÷����)��(��aĶ|�Z�ms����g�]u�Z�^�6m=4�l������ �փ�N4p5f�+�y�L�Ӧ��g���vC�g������4���̬_m���J��l������:f�2��<�Q&	n����&x���	.r|��e��$X�$hp��&�K"x'8�Ep�ͫ����e���e�9��e��{�<�ZP���>��&�OA�~���p�L���ckS0;�e
�%S����0Ǉ	SPʙ��,x�p�����=A��9Av�HN��ۃ�+����r3Ͳw��w��QP��E�Hrp��'ì�H�t��X�9��L*��;���q��q\�'��Mt-UKk�޼����#�Ӄ�9�:�ŃѾ|]��w;IF�w�NFۻ}����1Ӭ���;=Y�M��du�k�r~@���'@�VXݬ�?�d�1�����Л�q�\���{�d5���jꟲ���kr~�(��-J�?%���^��=�qxW�4��|5�wl��&��	���W[�Y�h�3�����[�Z�{\��R�γ8[����R4��U��u�ť!2��?��s����-��:x�����E�ٹ���G��!����f/mS�˥m�v��6sv��͢]W/�O����x��Q��w\i�p'i#��s�0%�5^p��`�{,��Ա�?�����Z�i���k���'�7����i��=^��b�Z��{BbC ����k&rO��N�돎i����V��^M��nc
���7x+ xk=?����9��a�q��B~�V���H4)�Vi�Iٱ�R���kM��|>�K�	Ǵ�Qn�|{�e�����������;��_�<�'�U����'��7��>,�Jl{w�{�t-�&�'_��vm������u��C	�j��"�r)���"tV�5��#c.7�DKD�,y����d�\����D���;�vtU+�|��u��~�ᇂ^��y���0m�+�-��u`ӧ������ԗ�Y�GNq^t��_�+ש��C�#9{��)�U9��H�kn�CR&�Q��=�U��J��:�4Y�0A�pg!F��w�[��]�8�����փ��(�2���z����գ�%��%]�!I��	��7����>n�"�'}W�wh�A�	0�Z���!���E���`sX1E�͎#ۑ�,��y�mѮ��su��0��N�s��!���y�*����Bx3���2߫9��J��6�Ky�xz��d��D�����~�Os�j�X�d��+O�'���K,SGX��`���Iv�5XryB��CzOc�3	¥�'`x�����A�T��=�wr$����H��
����a�z���N�aK�#P㾎�x[/h"�L� ɠwc�=0��"��"�Z�!�a�ͣc�""؟�t�yx)7P	�J�P���U�U+濵���Zm�kᘯm�TpC�B,���ٿ�C��4���u�P��7O]ȿ���A�i�I��;�J��sl�')�XK�0y��2��R���7��?�:��ډ�{{�KStn;���<�]�>e��q겱j{�_R�1�o朌*���5s�G
����H�׼hx�?��+���zN^x�z'<M�EA�lqDQ���T��9�"\�8��Ж�iڪ���b쾗G���(2�}��|?�k�Ca5�֍r�>>����Q�;ƭs�k��c�X�B���(�o�AgW����Y�}.��I��ȯ�` u��[��m>��Ç����b�gv߷�Ĭ���:�5B�Uy�������<�V��%,Բ�G���ud�$�h鉐�e�خ��|J�rvc�Sg��v�93t��~q� h���)�0�m�諦p��̎��:��~Է-m-I����\�y�dk0��/׫�87���I&�1�F$jLS2Jc���bV5H�O��
 �
��x.>b��U��}ß�K'ԉ�Yy��\pw�Ɣo7�t�#�ȏ����t�����%n�?�ycVɨ>EA�5�/��7Q5o���[kW�.Ǚ����|_Ii,�it�4@���#�5R&� O��b����ٴ�$���[��
�f-�����A�Ԑ�z�)��E���ǌK��w[��	�����T1���W�S7��Cѩ��� a�fd j��PtM�t�i�Y݇�?O��^��gu6��8~��c]������4@D����=ݗs(+���y�oN*��u�9ҳ�����y�:
F6���ՇEA��{Fҹ_O���1�+O�,���3[.�O���Y̯ź�A�c�7뵵!9��67�~٥��r�+Ĕ��.����Q��̏ɲ4�TZ�.�g�Ռ��>��6�7AǑ}ڏd��+E������b}`п��e��࿹o��4��Z��X��]�3X��E�tYG���k�?g�\�� Dn�+◔���/�~8ɧV�564!xkz����ƕ'�pk/�������v���Τ���mi-M&G&�|"���=}'�aH��"#5���i�c��]�4��>�{��e(�����^�՗6(��[|��:I/	k���1���/�e�ŏ̉t����w�lw�<>�]>��i?�8�-�km]c6��-qġ�#�&W ��2�u�C/�g~Gi���`��2��;nA���<����D��U-�ӱTD���淣����C�V.]h�U���s�Ο�V�B,=t�Y�O����]p�N���<�!~Y(lZ�t$��"���6-]���ۉ�\�SZ<UU�~��7i����VU�\�N�Z[߽C�\��{g��/>?�����@�o`�w37Βn,����n�� �hb��氹Enw.A��Ǆ"�6|*�0���}L��GuۢerIÿL
�?
%r;RK��C�b�-�䵗m���u�w��J��1�C6ڈ/��Ä8���}qbRD���Bg*��zf���B|�ʠry�� �� ��1��������:_c��A'�4�����P>&J�\ޖ֠/���{�ɜ߽�ѝ���u1�e��Ԭf����D'�#�E�0Q}�I������w��V��[�oo�}�(p. w����w�?����y��x�_(r��UԶ�<��x�/[��o=�]�nwgw�L���[4���ZMQKݐ`Ǩ�$�>m���s��C�.Z{�_r�^���$�C�����%f�gŐ).Į�����wN�lޢ�)mh�-M�K�~/Ѿ�7�3�����/�u�]�� ��!�bI�G�n��߃�~�q������}Ź�d�D$�s��AK�2�A�:T��D����;i����r3Zص��Ij�}
B�߈]�S[r2'm}�54��A2���1�`�uB_$����+��k<�m����c�]���+�O~���tRAժ��̟�r�Y�5}�.lb>���I"�}8��d=r��C��U����q~�����}h��h��Rk����Kk5.���8xK��>���-k!	�ۉ��-�}�z���ۉ��-���#J���m�F�V*��J�^P*���Fo(Ak��7!��gt�2����A�@�e"�΄h5���A7Ƞ;K=�X<�֮�w���֞x>�K�}���������%�'�?<"G9
�b}U�y
��]��6��A�z����V�ە�o�)_T���y�w��z����z2u�PS{*<�BFd�3�a�)� G��Y���!�b5��B�(["�� LTw:c��y>����с��!��P����Jʢ������/�$�p���b��-�|��
����	��GR�K��o/R�O��!b���q��}�U��K��$���ݐ��6�kC���Zk���J��Ե���ڔ�O�Fo�Od	�7 ?�����ߗq��=&x�Z�#�Mn�l�-��,8{\/�!X"���Z��/��$��JD���D
�v�H�=#�h�&�-�]K��$�Ґ@���R�$��6jWe���8K��$_�U�o0	.ȗ��4<��DS���Yʇ*�幠zBU����Zb@m�Ϗ�]��'����u���h�����=!m�����a��-+jЖ=xZ[V�H(K�.y�����+��6M�|�)R$I&lM2;	n�i��2z���h!��[�lo���e5_i���}���SM�/xiJ��UVZ.��J��F��}[2��%�W_�_җH��T�Ѥ���PMG������	����B|�!�= �g.H��GGG�QGC�F��ضlC@�(��>.
����Mg�ה�.M���g��%��S��b��	���41�QکX�!*}�.�Ykw�%;�uQ����{^��Y۞Q�G�S�#�	T�
S����k?�G����LЉr�����p�H������m���-��7��@��;���?�L�9����P?�?��I	T�@��GϕnX��>�s��e+��ʘz�{���>ԗuIS���>��U��)xvC0��W�紊�<Ba���v�0j�6#̀Nl ��C���c7k;����U/˧T&�k;�+����^a��2N(,`�D���zd�J`=���C�6��w�	1�g�,��N�x��¬XX6i��T�t�gݭ�{60��r�V�!X͂�� ���wܣbu�7a�>~,D	c������T�I/�ŕ�~(㎬�� ��ܱ&���!����B�F��±*��X��؎`�)~����JH;�݉�a!�M�o@��nJi��X�_#BB�"}Z���c�H+i���MQE	Z����B́&%�d�P�
^C�B9u�g]q��]S:7���9�4�	ʎ�Eܻ���q����@��<�����u ���Q�]�;ՈrLnU�<�Q��s�,G�q��}
��9�|�x�Q�(��LE���gY)!RC���v��`�ݑ��;�Y�!A����(��놲醲�f���!sa��.��ά�+n�����5�Ha�"���H��w�C �7�3u�h�|�|�:+� ��ۊvκ�sɧ�p�u�?G��p�������DY��yy�<�����m7�uA=uI	���+y���#z}��"��h�y�9�Խo��}ك��W�����=��[�3Z�"x	��#�
ʪ����!�O���(-���/tH����O)��N*݆�P�)ǕY���� �@/��if]��MA�L~��|Y��;Y��c�$�(ⓗ�?�?�ZvmZ'v-�^k��ĩ�����v
&= x�������]��W�g �i��zf���i��'��S��Շ�p9ɞ9�9I�r��%!g?������V�櫜�<�U9���7@7�M�n�qL�6�C
>�O@�zB�zBVz�|��e��6�dx�亪7tU�6u}[��~7t�����B/ti�蝜��@�2�e�"e���
�9����m6|t�6�ԩ^���{�$7\�]�?�q��)�� �ue{S�_�y�J ��e�2L�N�G��^�Lf\nj<�Le�+�����+��5�+���G?��/t/��u�[�v�}2��Y�T'BS!�z�,R�a�\a��2�<A��C��C��A�Z�e��/�NK�NC����Ԯ�/��~�":�ںҩ�:�R������op9
��fO��"�ȣ�e�I]��zk��A}r~��/xF�κ�> ��ր|}ɺ+GY禐���n���YW��:��Y�S�d���+����?��Fh����z��9��K�S��O/=�A�Q�K� ��^�DX�IB����?"u������^BP/���:f�z�����]��<D���+�[�=�i�fB����8�'�t�p�uh�{����BQ�]X�Wܥ%tzg�������@o��myi���e�#d��P'Bo���| ?= ?^v ��n���uB��B_iч�͜}����m���Ah�3�^i9J����r��NE�-��9�.d[y�P����Q%�T�Y�"߆����n�Y��¯d�ۯ_�ual�������2��.~�K��~G���w~M��}��7d��9@���n�|��^�Gw��[�����%���y��.�I��#܆}*�cm���%�;�Jl�����v������K����E�?��x^��8H��ϛ~�;�^'1F�F���s������%��oJ|J�;W�I�t�iGK"��D?���xZ��ߕ�Mb��g%>,1_�^b��[%��x�D��s�eyJ�L�~�5+e~��6]�U�S�H��X/�kg}Kz�#%VK\.�V����%�%.������<y������wy�Y�q�����*��/H|E����j�}��u���x��4���O)g�J\ q����{���O:�Sb?N%1F��oJ�:(1T�_'�O�X-�	�s%�J<��w���|�k�������Se�V�K|L�R�+��#�5�5J�Ab�Į2���J-q���e~���$�w�wHz�%��-�o����5��k���R>�k!'�ey�H:&�\H�\I��O��[�[ܟS&��i�fCfv��~C!�Ŵ��ƬL�A[��X�g����{��J�Y�QƘܙ��rY��(Ɇ���%7��6~�V�=dPv~>c�Y[�EVC���P�	ƙ����O5dY��e����i�&��F3jN�3d�R����� �b�,.�h1�2��l<�')o�9�<�Y�S2�c��Լ���	��i�����͆B��'c������2��A�dȜՊ%�G��z�1K��m6X,�c	�V��U�1>AQ��@�&"%�,��YH)հxC���*�\�(�;R�'$9K�Y�͙�W�m�QP۠B��$c���<����w�}�*�0#�Bl�gZ,�����薊���OZ�*TN`�b���*��bMk�3���'�9�ؤԄ'��}�ٲ,yY��t�i�,�6�9�К�f�i�f��y�������i�!+/'/kZ.�[H@
���e����묙M3�Y�"eZ��`��|^���iYܛi���i�Y���,!!n�\�����A�=�-k��@��k0#�ݠd,(0f���i9�U"BN�4��Yg��S`��e��<F�QD��bc�Ҧ��͢|����
���<я�i��!�4�3�������Fk^�l���$gu'0TF�����"�y�G;�¦$�OM�
.4lJZ�Bg%K��4!bB>�P����s���L�b͟�g�e�O*�A,{�~IF��E�1E�\n������e��EfC����
� ĉ�)�!l��Y�|<-"?���?A���N֧�x�*���y73?�0o-q���b�~��%�$�]n�I�f�'o��$�o!�"���$Gb�Lm�57.?O��ҳ�4���Y<`�}��j1�L0!�fz�b�+�����KI*J�I�f��28��R��&6�t�En����"�hݓ
E{�N(�2���d{���k�1�(_jC����%Eo0sQA���H_���zZ^��܃�M��"i�T��l�IAZ^�AkAZr��4��K�����:�%���0�$�P����g��8[hV��f� A+�HeB���Y�Qt?�0��c�7Ha�S��[�����"�в\��k�AYr%�>�§:�?�b��������{�� ;�Cdl��I.ʷ晜=JBKe��"uLl4�sW���N�<{.t�	P�g�}x�g#�qJ^�J����5h(0Q���,��#{��,2��<���{��Tc�ӝYX.�&	Ş���EVO%G��V�9o:�l(̗TE��a<���ٲ;F����=4���
D�~�~L��"=�32�$����.�*�-WOA�ea��	hN��lT����2�y ������N���w��u,>�bʴf�%��Dy�}TɖmW1��F�7�w��F�V+�#����=-|�MEyΘº�H��ALӍ��lv�%�����B=��>>Ӛ����#��t��^H�M%���W;+3/?s:�T'��{�/Q
�L��ȅ���e5:osV���H.r�$SuT�ȃYvC�{�͙3�֑�:ãߒe���9֟�q�� n�2�S�ӌ�����Li�y\��ӔQATt��Ds���n)�`���+�Y�l/N)Ipڧk�`�J��9�y�[����S�]���<.H��XR-��ū�Eňf\�-�Bn*��2�7�3-�T�dCv^Qc��8#��[5x4�f��������_�)������sT�"p._?p��pΑ�棯�⩑X%�Db����M����Y�R�c%�Kt�,�-���~���3>rW
����$6�S�K̐��X���Wb�Ćr��%�Jd���%�%�H���|H̐����/1VbC��_���}g�|���K��~����ou�C�ɋ��y�C=�T~�pwK��Y����-���%r�3_�\�ryk�?����Զ9�Zwq쁘7����g�_X��������Ȯ���GY���G�X�l�2m����<1qR�-/�9]����[�/��J���%6|��_!�]	[��i�Ϣ�{����Ï�e8g)�d8�$Q��I��:�R=�Z������Z�����_��/D��ѯ�u��oe��eKF�@�mU��K��6�X�k\��U�;�����^U���7�����1�۬bU�����xg-�������w�>�:�|��WT�40z�3xW�|���X��x���*���^Ƭ��د�Nu�p`\��SB~u���� /������	܌k�@��[	0���@�i ��:����6O�~X�� �}}��7�$�I~���˯����;8�cAg)�S�>��pW����;�
~N�}
�:`�Ep�{|]�� �pL�� ����\����g�3Hu|�K�� �� /�����O���B߳���R��x����o+�V�|x����ӟ���F\���+���n9K'T�����J��y��dq�	�@~�� ��̘��6c���x�K�����>䫰x��l����+,
�����Q/�op����
��� ^㯈2�(\~z �q#n0*Pa�K0<H�5�� h�����Iw%p�t��%��8�R.����x��"�8�����`����lo��>'�����rXl�&�����&x���i`TO�V�¿�|������:�-���s�E�yQ�V؀>�~<pv����ҽ�]�w��
[}���x�z�4��ï���M=�{�"�&P)�<��Dm8��nD9 ��aj�����[o�0�w����	x�`��v��g���Xr��vý3Da��|<Z��x�-�GZ��GnS�R�y���p'߮�*�0x�v����#QO��R�ݣP���|���G��6��C�쇋��M���D�_����?�E��L�\��ý ���(O�sz�O�d�H�r�ɢ�~j����x)'@�Y�P����Qz��D���������:5O�)�9t o�$ �O���W��6`�d�.z wM2�ȦH�@K��g.pC����d~�{�{?��]"�E��Qn��8�"�T`�to^��SQ_��<.N�W���ӄ;�Q���s`�t7X�%�03[�%�+G�#�so��碬P�����D9D �0��M�����y�S�
�K}pW��x�@��XZ(��q��B�C��FY���M�I�#f*��Y�@$0�,�g �m�|��n�z�p�L�=`�����m�&���y�+ECu��H�?�ަ�H�I`�l��V`��`�t��>C��q� �J�s���P�O�yP�����H��ȾZ��=��Dn�3_a��v|X�|�Ta��_�~�0�~0�Q&��#�~>>*�hxT���-�< ��dWHw0�1�S�8ٮp[b*�t/y�`���>_.�V��?�.�&.��R��@�Ƨva���?���p}�z�%�]��|q��_	��9��\��~3p�2Qn5�/��t g� ���T)l3���_�	�Y'�/0v��_���p�����Eࠍ"�P`�FA'8a��O���op�k(ĭ �*��q�h�災0T�]
�]Љ�e�2��~K�U����-�G�<��7���>t����n?`����'p�^�<"ݟ��ᛀ%���+����tw'�'�ONz_af*���"]�~����
�; �Xw@�Wp�"����zQ������O�#�3�0�@݇"�8�C�UOA]��GП�6�1�},ʼX���c*G�;���}x�p�?WX����pk���v�`��w {�D�$p�I�n1���h9���d8�z	�4`�&��(����� /��{�"<df?p�y��u��?�����p	m���f�,j��"���-*�ir���D{����%P�bO�">��I�E�ݾ��t5p���8����s	��?�i�wt�はta���E\��/�������*�.H��F � �C60���N
V�z�
ԅ�z��!"|=�P&�|W� �w�_�&��T�E\?`͵*.�u���C"�E��7d�~��}�h
��@��[pY��S	\rh �r�����{��#7Ag n�@;3P�����x!J���Y�FG��ݨ��b���"�y`�P�?��-���@�m­���S|�v��z`�������u4��i����'�xN+�\&�	�������xQ���cD�`�X��$�g���8H'��KDY�����q"�f�-I�C	0 Y��7^��GOT���Ly?�JC<�	�e2�0�3��D;�LW�~���K�?|�n�^<��l��H�~�>;U������J`�{�&�D ߸W�Us/�yB�����D�#@u�l��ҽX4]�k.���t��w�2�ޔ'hf牸���y�>��~QnV��|7x*_�y���B�GUl�	q~?0a���,�)�p)p�iCN*�����1�msT|n���\;7 ����<p�|�E�׀g���l47w?"���]&�FO�#Op;��"�	��O��h��m08��w<��K��=�֋o��p��}�{���~�q�x^�r��|��z�+}��p�$�w�-ó��;��e����2w	�k\Ki.�\�W�������n ƽ$��Z弗�~D[!�|��� ~����	8r5ҁ[<���t��u�Auչ����o����XI$.z��M���+$͕����
�m�wP3��Nȿ�
���e�>^ϫ��a|��M���x��d6�%����5�fZ(5��̓��h�YFZ!4�Ϥ�1c�h,����LZ�5��l��Ϩ;��G�8PC�c�y3r��Ȭ5�yYf�Řc���d��5R�L��P0=��ZF�)2�n��5dZ8��2ܞi)4��>���¼��:ٓ7OR�نBk�uv��?Wn��*�Mb��Ѭ5g��YY�tkd�̂�[�� ���q1?H�ұ���i�S�J����j�Vɍ�c�+����Y���e��k��@`-;Ф��:*�dca��h1�3$"Z�E���/O411�b�*2��=�3f���zsެ�|����w��b 6���ޡ�O�(/Kb�,��s��A��YT�#��d�[-B��l�Y1�#+#�J��9�7A�\~���ɴ�X
\�l��D�7��R�xY��j�&�1ws�(������I�HeVffy��� �<���\�r�a��a��P\�8�f��h�
�8�)�>�D���&wN;��@��,�r����6#4�̈́O\�;�u-g��,<nºC���x��t��3R�gyE4�W�n�5���4ne��� `���f�ݷ�^$b�d-�>1��� W�o�߁<|4\7rzQ��QyYyZ��Y�GI���"��Ix6���21��(�3���Ѻ��(�Ax��|�����QIW��7!I�"�	2d���Y^�W�{����}�/��9g٬<Z���7�zV�R6|l�'�	�jp�dOI���T���h�*��5z���_<�=&#s��X���9)�|/ɤ�6�W�.�\'�"�u�m����a���I�{�-��9r�'����Bߺ䤙57���95��Uw&��^G\��v�������G�d�t������:��v���@<Km�8�2V�.Y�h��*�
E͖��T�*��%�u�G+*�M���ٚ�5�5Qk2֘֔�ټ�fM��6d�fm�ڨ�1kc����צ��][�v�����rי��+Y�h��uK�U��Z�yݶu5���կ;�.�:�ZSYUS[���W�WgT�V����K�U/�^Z]Q]U��z[uM51��E��[zeFen���\.�\\������rs��p]���|%[�:du�j����Q�cVǮ֭֯N_��ڴ���|�ꥫ+VW�޼z���u��W]ݰڱ�i�y���G�#���5�ktk�k�Q
�(�b�Ģ5��,]S��
e��R��~��5k(��(!?�Qx�R�@9�PR%k�]�v�ڊ�U(�mkk�֡쎮mX�X۴��ZV�WR^E�US[���W�WeT�]nޥVW]_}����Q�T}����[�>|�f}����1�c����ק��X��޴�x}��E��_��b}���뷭�Y_��~�����֟_�6�m��A�!rCԆ��t��7�m��Q�1rc�Ƙ����7fl��h�X��d㢍�7.�X��j���6�l��X���Ɔ���M�od��6�l
ߤ��)jȘ�M�M�M�r7�6o*ٴh��MK7�⤶US[���W�WdT�V�*�+J*U,�XZQQQU��b[EME]E}�ъ�
GES��
��oEȊ���+�VĬ�]�[�_��"cE�
ӊ�%+�X�b銊U+6�ض�fE݊�GW4�p�h)Md�V���U��t���2V�2�*^U�jѪū���XU�j�m�jVխ�_utU�*Ǫ�U�W�+ʢS��qey������:Z�P�j�:_����Ѿ}���(iق�g�p�:JoUK��6m޴mSͦ�MG75lrlj�t~)5:v�U�U�T�Wh*"+ڮG�J����+ݭ�����'�r7����*������\h 0Q��2�?�Ϧ�W��~+CV��Ԭ�\�2fe�Jg9�4�,^Y�r���+���XY�r��m+kV֭�_yte�J�ʦ��W:e4�RSYU��Ԫ����+�_���������_�݋M��qK�j;�bb�B�\{�ّ���@�mJҁ�i�y���a�,�de������P�W���������GH՛��~m��Ҽ�VܟcJ�P�WS��ߏ.��cB�5'Gr�sL��ʥ�-y��ѓ5�w�7In�UJ�ҁ�X����
&�>i�p���gE^Ο/�]�}�8v>��0Y.��\�k�T�p� [�ηo�kT,CȌ.���JYW��:)O��H$�����o����Q^��a�vƠl��3�(�Nٿ�{^��2[�Yp�< /|`��*\� ��-Uu���b�}|�p��m�&��Z��7It��۾Iz��ߛ�$Q� �M���C����]`6��%<�0W����;��Ј��@'=�������Y|�����a��W��z~����g��/=����	�ŧL�����=��7?����n��k��k�8t���1{m�c�ھ�u����v�k+�_�l��{���u�m�譶_�l�m^���M��V��V�s�-�h�-t��旷��F��)#N��?=i[��I���N�ⷞ�=�
[�-מ~�M���)��O�n=v��ǳ'm읓���6����X~Ҧ���v<{%���9��-��)�\��Yp�6=���ﰓ��G���+;aی�X�)�z0�=eK��mۥ�� ���M���1�m �H<��q���L���-�5쎓�{�?�|�f?v�vz�I�k���j�~�V�+q�O��O�������B�;nSF��i?8i{	��/|�v��'m8i����-y��TN�cw�z|G,�k?�a�4s�M�~�mZ��l;:�e[��v��~;l��<��gZ�Z�Я��}~�ۛ��mߍ=b��5��_�M��C[ ���Gl���Ķv���f<;g�ж��C�7fؤö�o����-1���A�a۶�ö��a�8����a�߫�ls�셆C����e�ǳ�ö�S�l8d���C������r�.X�mIA���|��>�s�6������aɾZ��ѣ~T]d��k�֏����Q�k�G��^ϧ)k^��x�sƚ猋�;k<�������76�5��U��o�����o=g<�n6N�=k�q�m�l<U}�8��9cb�Yc��g��
�0�<�x���G�=k���C<?q�q��q�#�o��7����	������ɏ��	�n��I�Wn��<��If��t�KS��6t�E�\��ri��
�4�pO�:�҂��9JpYe�k���塊��E�Z��M��_ߩ��0�\�������ۈC�=� ��ZF�:M�Lٲ�)ݞ`�g�;���t"D(W�Ե�V;5�]����_ D�B%�P�:���cc|�q����	q�dhܮ�*��&���󷨪�Vh_����Υ������1�N_�:�sx(S���k]4�q�q��{�*���^w��9�m���.�����:F��5'Ks�4Û	��,��B>Ns�ɸ��9[���� \bX�|j�k�:UΝdZ�r���gLlj3�SY�[��?��[�<��5Co�L�j����tiV7�?���y=$����O��\���s���~^&���{�,<O���B����.�>E�$�n������J#s0�	����c!���S���}2[���{^���ƤD�/�F�^��W��w�@���לEIz���ܯ�{/.�?����<g姱�<�bN>��Y��Rd��ӂn�%��>��)c�dJ\J��^ &g�N)e�-�ɠG���
Z���k?>��K,�ء��~�?�����觶j��U1��O}���ۀ��)h�c ����%�P�-|V�)��8b>�0[loΛe�����O�Oa�oU�y��-P�>˘��e�(� ���l9S~Ƶ��\���2w]|w� ̿�Β�TӾ!��|V<_���Z�{ś�׼>oz�'CԧoIKbb(3�9��p��>l/�|��GåX�u���kʓoV��ɼ���(�~6��Рd�u��?����P�B���^��ڊ�|�.��M��'��Uz}��\��[�<�V��J�?��2��{���r�׻����šϴ���V7�k1��͑4��Vї������;J�@�����Y���,���:ڳ65�w�"=��$h�Tv�=����F�:�9���i��x�
a�\k�y\�% D|��+�l��ߞЬ����K�����/���bC��~_����u�����b������iї��%b�˱ӎ�2p�٥��FV|�����s��^���;�S�<�Wb9���Q��ʜ�o<�����{�������g�}[���?^�<�q��ݏeW��]�����S��[�fʻ�*J�z�밃)o����R���Vگ��Y�TT��]�����:�Ѳ�n��o�����z��p���s-���r����+���K���6ۜ���k�T�K]a�j���9�E�v~_ԥuS�;��GlH�7�]��-���Ӹ}R �&Ԛ��Ļ|#oW����y�3�"�"�� �?p0e�Sy�������^��|����,c��%:��W�Q�YQ~;�Z�M��x���*4ށ���-ip>Rgf	"
�g�Υ�#�鼊g�~�6��!��Q���mو㖤�
�!�ڲ!��V$��֏f�~��#y���R�i��TP<��(�.�8������V���TL�7#������Sm-g����eA��1w�_�v���Obe���������-3�����I���m>��g"����Ւ[꿫�li�8�m�ih`�;S�	����Q��|M���-��r�J5��yg	���#�J�1b����IJ6��L.�Ӂd+���D9˭-Y��I�y���כ�I\&�K���^Ȕ�y(�S8�W��������[VP��Ғp����A����K%���f\%���L��S�ǽe�ϪU����)\�g��KL���)C��\P�w�R�Sf�����oL1�f�G� �;��ק癲�E\�@sS-�m�`.y�Z�ߎW����aO��D�SjnzW���$����)�ΑER2�D;�֘n�����{=!I�g~ȚM��r��h�N�ז�������@N�����i;���wk���	��4�b2�\@�U�e"�֭���
�K%	��Z\�����+�w��;��S�̳�8}�6\o�;�Z�)��zҡ��]#6��LOˡ�$�]�^��ٻMlQW.��|tf���+ٻm�*\-eR̬�yGk�:vׯ��BJҼ(�i��S��S����~Wj�����t��i뿚�y���w��Z��_���)��֔�C��=�i�㟍�;�l6���狷w��Y�]�4���hq��~p�O�ml�����]�����Fl��������������uy:PQ|����b��g��|�+�����q���=WIv�����gtQN�3�w��v�݆�j��j��2���tFZ�"���p;���$��q��D�=Ϥi � -T)P�h��� RR,	EiI[I@h+
#B�P[Ӳ�Qw}?W��Uw]���JA���U�E�TX�R�2�9��Lf�h��h��̽����{'�7G���jvw�g������'`*#�g&n��킮`�
�'����|U���z%��vωß�~_\��=�k���?�g=y�:���p���{�\O��6��g����_��Qb>Q����8�u:;F����/�+��\��Y�kb_����ͳ�;^{˟�䁽�T�_��/�+�}߃�Y/x� ��Է��yOӽkwL�ٗ5,��u�D�e@"���pq,C�I��c�+X���������X[�b4�Du��U�Ƀ:�K�]#�h�.zIK�C��s�EɅ��䛘��O�ș-W��"���,��@��?��Ճ����w�$W�j���5��Ʋwf����U�Z1��E�e\���o����X��]�J8�2�9��\�2�
������H��؜2�%�H�b��R�x��Uh��_Si�'�6N��"�~�i�¥����m#�����4��Z��Ĭ�`���%O�d���R�$D0��0�B�y���L�S���৹�����qi���>�k^:w��k��X"<�\ZD�j�槻��9$�[���\�i,9�ֻn�9V����/�ϵ�i�Ox#�_�*��8����_�>CF�>��U�	F=�	��)�,�ϸ� ���*\��s%|R�r��mx���/����x>�}�����=(��s�����>(�|�k��+>��/Zy�s�_KF�)�����c����?-`�O��Yix�5*�-q���C���_z���s��?>�_�Wl�.?4���>�&ތ_7����z�����H??9<������q��v�CK�a����sn����9?N<�.M4-��ts�rΚ����3�}��7�����eQB-)�v���b����vəR��U/�����	�֏~/����>/��*�q.@+^���ҥ��E��G��2ˮ���.#��Ͼ�����s|�����>m���-,�z>�=Si�n��e� ]������'m*��d��z�g�g�4�����a/�d�g����ۯ�e#;�m�$��U��f���H�����w�@8]{��Ol�-V��ګ�Ր	G<M�s�����w�c����i|�i�,����tW����������o�����'i}�0�����R�z5 ��V��q��?t�_��������m/G�c�G,����O�+����A�F����YY�4����1�_˔�F��'C��2�edg,���R����>��l�y��8/',���K��D�k��S���|�z��Oܺ��3��1�t�P{2����{*���֎��?��ש����̦Sc3����	��[�	y���P�G�=�B��O#�&ᬩm`��E� u��ek�.Rt?��(�SKug=]MY)�����Zα>��XQ[wk�i;Q�i��o
�ۮ���
_^�p}��r�Ϭ����s~��&��k��0��Y��v��c:k�0⟋�2�*��^�y�a�(K�k�>��ݕ�Ôl�Zj��%�ڽ�����g:���M͈�[.%�N�qQ#|���*�ӭp�j��bh�F+3���.[?�vO��/��*���ǣrDlm:�cO�OQA��E��[��g?�a��:U�l���*�̨{{'6��i缒��ߌOm﷌g^�J�k��g|8�)���u��pT*�O%��uN���v��N%��ޞ,��4�����=������11���y~|V������63���7��o2��	F{A_�[x>��=o��kT�p�܆���!���O�<L���<<�8��؏�{y���N�<쬽�y؝�����;G�����ޓ�?��M{�'�'�w_s���\��%`�����2�9��{?{�!o�7�Ȼ�',b�-V<�n��Ѓ��1;q�y�=dY��F6���àϋ[O�ף��Ė��50�P�f,3�*��id\���穇���s��SW3O=�v�S��y�?r����ep��m���bޒ�B��M��\}\�����������a����榻�W�8{]���]l|_���#���k��H�ܫ���$&>�F��3�\�P���hn@4��m�[!��R�D^��������ݥ��_�z��^w����2�_���Hxk���{�:=y�wO|_�������
/��h�%<wb�=%K��3�T�;r"��?�ȯ�9=��jW����Y��I{���s���*�$��1?y�'�����"�/���Q糖H֜[m������ڜЄe����m�y�C���>xV�p�/(�DV��o������/�g��}�kj���j���I�O�O<���ϒyK�j��B��%�X��{��9ɤ�_�v�'�΋�v�vg^�s>�WϜ�|Ԉ���2�"��,&��S�b=��D���zqB<O�ߥJ��Z�H�wt[ڔ�������ϋz�R�����e��7��2���=(�c��D��՝�E��&�Ӷ��7�R�ӑܯ�cn� ��c,�a���İ���7�3�,�z2\}I��zt�ѪbW4z�;�uQ�J����z�����}����G7+���r]�Pl�)�=�������)�6���W�[��ץ/Q��Z����>N�����tB��^����kg`���p�Z"z��5D�7j���y�hK���#h������q.�lb������$χ�d9�W@�k�e{�M�9��bf�D�WA��xb��X�PCv�$�����2;e1eJ�rn&pL�{Y���ݵ����.��Y�'/��^����8��k��L��j���➱��g���v�������M��M������*	�[�g�y=��$^/'(����lXO}��j�誄�M�1�Z���ѽ��jv������+:�_AW��9�cM��ۭ������J��ي�+�����;��}Z�׻��/�k<xݣ�S���u/1�8���u5��O;	�O����L8�x0J��X��P��F��fp�Kɫ��[���tʽI܏3>|p�ݏ�ܽ,���B�Ox���q�=��~���k$X��n�L&z��>&���%'q�f�<N�ߦh��E�����t-y:0߄��LӐTo���% w����2O����y?�C��F�>I�旚^��,�,�2��X��ϰ8�|p�>�[c�=�7�gR�z�����y�`��ΆOk�3�������y`�yaݷӯ�X�jg��h0���N���-�
}K��������� ����v�;�o���ۿSK4ƼG'>���S�����>��&^�5ޟ�8�ɬ��ŧ��a�纲V�k����5��h��)��Ny�~ū~����m��Wg�����Er��cV�ͫ���i��_qr�����������:t_~L��̣ܵ�f�?��Wq�a9���E~���zI��ڙ?�e��O3�%5���9U �jF��fg���g�99v��ޯ�(�>�����`�(�}0����g����w�|���\	z�⯌��סܑ7X�����_"�Hw�$�.N�?��&�A��é���x�T�D���
>D0&�=n���£���©����xԁ�@<14 ��0k'q��fI�cV#O��]����GG�m�T��ѼB���rt�G}OU�r&���}�~�?w����q>���7���`�Fř�J�¡H"���a4�*���n��7�Ԥ8�g{˖��ՠ&�)�:.���^�|=��޸�u���lwǠ�������1�_㺧�ϒ��n����^�WA�9��E����������̽�z��6���9qL�x��ws�3u��1F9�2[əK��C��$z���$�_ѐ"�n����M�v<����+�}���Ð?��央��w���5?8*��}Z�;�'�E�^���t5C�/���}���߶���dwo���c�V}�E?���;g�z���bθ�ʐ���ğ���_���L�m}L|>ͤ����,���&�~��?�¾��wJ6��k����4����L,�rZ��bג�+n�dv�$�7u�ʿU]'񾟫u2��a�35�~�tГ�g��:�5�m0�Hx�_��vU�N+s,
\ς��հ�g�����t���g�̟��#g"vn/$���Su�B��?UO�Ͽ��L���'�_�"��e�\��}�l ßRN=�(~ϣ�;z�����Q�;�}I'���#��y���A�u�"'3���;�w����4g������Ld��>���s�B;����]�{�0#�����LRՎ�L[�\Z��(�7�+~������뎜¬�b�潝�A䴐x�ݰ�hD�Գ:�_���m;Ȅ���~_�_2��*-D��~���4�$�0�Q%�T�c�tMk]���BWz�]����_N5�'nI�M���/�=��2����_�ٕz�R�Bb2����x�Q2�?-/�N����	GYt��}�e���F�t�����H妒�"�%4�� V�Y.���F��7��UF��-���J�{�����S[�p�t�%����`�~���=�����q�)�'�f1Qy.��D�B�Jy���xe�:2K��؞���v��c����}ޱ��9�S.=��Lz����V����;��;���qݍ/"�_�Pآ��+UNF�7�k�ۉ�P�]2ڎ翉/������fv�Ȇ-��4{��z�����#|�;&��F�:�����(4������&�ى&�@~���.{����ݒѳy��)��\ó/7�e&��2��M��PfU�)��U�v���O���D�m�qwn�$>5����/���(��Λ�DS!�����4G�{a��o���M3�U��;a.ɝ�3�*9y�-Gϱ^�zNw�5�� u/��ٺ�����<ٱ��o�S����c�[��2�K7^[��~�a<{��n�Tݬ�;��U&޶�����rre�Y^4�-��P����a �_2����֞W;�*�s��8�|o��&^zmǉ���;��3�%g�e��q\��f�������R�6{S�6q��<�7I[��6:��7Zj���;����,��_�Pb��	%�B�m�&VX�g���a�$�ksXx�[z��۫����H)�a�l��%�[�'�28�*g�a��E�M���\���qg ��ie�p|�ko�K]�m��0�@z���&�b�Ɨ�ګ�T����e(d���k{r�z\�[����mo���ź�ɲ��*�ko^\K����;�o���a���֝�v�x���Z��]�qx	3Ԉ�\��F�+ ]>�=���#̽������9,�K{�=��.���>�-]��khJk�7��!)򡻱/n���Dxwҳ;��J�[�f�@��ۭ[|��ֆS����uv���Kz�W\#��1��q�.��/�##�ޕ����,���R@s���G6+Z���WZ��!V�پ��[xt���ʂgxC��d*G-n`�4�uP���Ɵ,��Y����)m����0��`�}<\̃��4���~�KY4?ݽC��֓!�HK����]�@=�J;j���ڛfK�dq�έ6�ˁL9�.lr�*g�4X�5���"��f�o�{�r@Gn0�۠����Z'�Ky�C���E<,g�����fVa�� �p�1� ;U��?��P4jY�dn�q�ݞ��y�����T,.�G�z���,�n�R�@���>#�i��5��lKc�?���3[�+ Dí"�D9�RG���z��z _�l����M�`v��t�&�HUΨ��/�g�옜��i?k��8�py~��p_}GGaG�?��b�l��Q��8{D�B�� `Mk�#�]��5HVҡͮۛ:�����џ�_d[U)"8,��ނ@��
�+gؠ<��U���fB�x�谆JLD[Qтm#����̙\�8P�{#A�"4�%���x�c�~��=������j�&x0ږ\�<��MHB�`���RZB��� |1��P���{�?6h�
�1|���~1�������b����Mz�j<��
5¯f���#%�Ƭ�i�LdW���@;��K���Ɲ~��cP�e�=�Ӂ�L�V�[@���s�6�f��[F�7d���M{�jZ�U�����T��H-)y�&�`�	w��m���Z�n4WP�F9r >l�d���"g<|�`������|�����Џ��d_����� {�do�2��V�7��Z1���}��(#C��v���<��;p^��j^�4p�1�����E���#�>|�0��h)-���2a0t�W�
Z��!��UY�9��;�w�5ֻ���k�?o�����>�/EYz�a	��>|��~O��?�_\�퍇/�1�I�gwJk�U�P#6
��e��_�x/�x�zKp��8�
a�a-*��]����rƣl
J�� ��7��^Y�r������~n�N�g
��H�`+�ޜ�O�؈W��gKm��8<�hi�)�v�ZV�o��C�ᴀ5���8Û�~��T��N+j���y\���1���<qck��V!,���r� <�����L>4y��%A��C�`���"���`��%���7�,\,8�B���,�C��_0�#0�g�eo
����)h�Bp��f��#!�>��/�A��AuU
�U�AFy���mi�s������HK5��.�I/����n�}b a��pcA�bN ),~j� ��>�]�N{���a��[��3{����=�8{�qq�{���ǫ�� �^zł�E\��� ��˻�
�F������D�t�rW�}@ݍ�`�P�zI��{n�g9�癩�����Q)0NP���<vYx)Bx� �����D�v���M
�LT�joi}�Cu�1R�+�M(S�^DrFvi_�i�kI��G&��L$Q<򋇨|h�N��J���o`a��P���A���z*���p��"�~]�ͱBC���5"gd��-���hTn�Ȃ���d=�'��W�cG<��M�i�Ë�G��I��~�Qtp��m��,4k�S���q#����	6���j�v~yXQ�	���n��t��49%4�,�>^s,lQ��D�&J�>��O��T��6�AݵE�%T��*�
<i�f�3��c���$�eC�� �sKs��M7�*yx:<�!p�u52+�*��8]�7����}a䖞be&��<U��(%`�@����]�p���� :���@/x�
�))͠�T����|h���c�@�ݛ�!�� �]�Zt�Ǉ�w�ё��n�����p;��υ���C�3:��*S��* �	�G�*`�Y .��C �7C�	�&�N��9k`�g�4����@/��%%�ᴆ�RPJ�_;�A *���z;�Xl_�,�^�O)�[KWTVJ3i���e_r��|r�ڪ4� �|�$�W�8��:۟./����
xN���re����<h#�*w.6;��Zz�y�^�� �r��@��q�y�F�&�k�G�ʹS	|��'{�7��ҭ�?y�>Pmo����B�m�"L�4X�1��;Y=
� )�[*�8ܣq�t��p6���+{FL~��ps���jɟ�5:,@K����U��ľ�M�ԞR.�9���Z
��[aA�u�9e�P�ov��uˬ�֝f����ط �5Q��"˻O���\DҼ�#xE��(�3 �M���f�So^>��Vi@1x�K��\ہ�p/@�`6��3�47D�ai1�psʡ�(bzU�L�o�.`&��$o�2���r`�-r�R��#���@"n Gdˁ,2j�݈��a9���tt_uM��q��y� \�Z%R3��ٜ��jN)ɤ��4ve��(�<��D��S��f�fs[��V\✫ˏ(������P�C���*����b&(z^���yb���k�p����溌�ɈD}<�t�p蹽��:��5��z�Z����p����\��g��q{\���)�� �7(TfFw�Elo��qX�9��4�7�A��͟�^8�x�Q� d|�����e9N�[�0�����u̎���mu�{�	�J�}��?e;�۔��u&+.M��P4WW&�r�m+�FV'���� �X�zi\ �vpK�4�ruQ1ěu:�dQ�?,�[ᶰ2;T�#+sAv	+���Gq\M4��H�Z��|&���Xܞ���,.��|Y����l����-f��fo�F�<鞞Ԙ.P��\��a�%5��.5ܡ��>��6}(�,z��_�l���	��e4 =�&{�:��=ġ����%^w��;�(MsO��[%�:�%�9�%��=@��?�F����g�cyn����(T08��y�Tב��!��p�@���݅��Y�U�s�͏F��Յ����Gi�tFɦ	"5�E|t/�x`E@�9�-9b��Gv�{�C�����2r(9�X�$nǊ}Bw��
��[.���E�2`��͇�.D[3;`�E'�`1r	_Ҩ���b���� :��V��=
��"�J�g.�ZpA.�4��a7r���F�rC�A�s��Ҝ��������F>�?�%��˲E>4���'���r�]�@��DG��m�ܒ��!��Yz�&��a�d� ��N��a�HF�><!�s��G���ԩ(����r��ԸR��"9 ��$qI��7T��vy- �T��[�&�a(oc��;n�"=�<+���{��T��`��Q�0>���b�$����&���E6кV�
�:��+Z@֦íL eT`�����L�Xd���6�d�t�DV���XEk&=�ҁ�qL����������F^��t��t�W����r���'}��3�%=��a�v����wxNg��ʲ��?��I��Y�e�?�� ���ed�t�T�l`�����x�*ci`Aș�ZIN��*#g�OYp�M�%�`7WZ<R���3jh�(�,���ZrKG?�>� ���q�Y)�8��ş"&U�A�C��%���Y�rA�?�#=4'��~�N?l�ǭ�&�@QL$v����b)H�+t
ҫI�H�h(c6�P&�=��뒃Պu�B�۽s�Q8�7�w�q�)$�"}�L���fz]}�{�Pu@�S�>`����^��g�Zk��}�����������T���/�6����4x���yO���W����-N�0��s�q�O�#���ȃ׫�<h�CWU�Ӱ`<!�jN�G�h���TB�J0V2a!�����-���Kބ�S���	�W�������˧WN	����>�{½'<js���S�^v�'�z�t!�C������+��	�cl&0��u ;~X��}gA遴�����&x�}��3Bu�׈`Y[�B��r�҄������ #Lw�M�G�S��N�Vf=�3Ƨ7b�R«!ꍥW�jR��OvM���pB�ί�r��ޚ�rI��c��� |C7���g�;0�����\���u�-�ﴻ��[|��U��$r�Z`u�������W�׬Yr��ƨ�PN�����_҂�NH_���z�P"9��,i"���J���R����{�z��'�A�Q��c��B���1R�.pt��r	�%9�.::���!ǡyhEq���C��x9�؊�uU��8�N	���� VjJB�?S�;y������V�{c�@�V���6,BW�Q���>�z��K��\aK
��'d'�y�?c�P��3a~�N����l0�:��}y=:�g�Żj�^�Z��
>.Tm'�Oڢ`����_AXPP��v�Vq�2�w�-��#��I�oH���	M�d6�-(�[�k�%=ę��OY��`Sn��K$4Ր���]�L�BL�`ڄ��� �7�*갌��rK��F�E9[�!��*�F�Dξs`6���4��:o�f~�zd����O�Ёҿt�}ؿ{E
��{�C,.�Y��H�8 ���9��?���
9�(Nm"���\t؀E��XP��q��t=4����-ҵP�9f���h�n�^&�+H���c��PGǫl��F���߯�Y�3�b[�2�������	�*���w� �	�Ls��9.)H��������,���>�̪mp�HFO�6X�*C��F$����tUz6�}S��k &��f��m�G�n�@��l7�X�GCs���1�1.;F���y�t�a,�8bw�*<�4"�K�4Z����cvu��G�í�ۃ�@�V�
��ۏ3j��w��N��˸��z7�נ+�+y}�I_#/���nO^{+�5�����V�w�aٰ7�InN�<�\�74����𷇙kjN�����)4�*�-t�y�Y�ڽ�����/�����K!�Z��Fܮ���u��|5o�y�ݥ{�b���Aj9�(�銪1�j�Vm���32���Ȓ��'<H����#s�Y@���,��Me����'�����d�f��*����q�tÓM�bۍ�p#$���"��:�A��U��U}�9�ۇ4W���3�mz�]Ժ3�2}EFO�g�zM�?�̶�,��4�8��rm�\k�� �mDu:\*� qs�@Z�QH4��H㏓�v�|��!Ǣ��E���p/�dB��jbK��T?*��,�;�c����Ă�t�գ�������8�SP���͸��L�@	r4"):�:��b���h��!��&�]��ĥ�I�Fd�
g�=dÜƿ(��#���%���@�b}Va{Z��,pX���t�IH-pd�3ȥ��f����[Q��on�P���b�\.�B��O�g�??Ϳo��P��eޒ��*�/E��J�/�����p[ښ�p��R���c<���>X=kb��C��c�h/tt,-8��ѺU��t5�3�������4��6z9G�u#��7^}��n���ʧ�7��6�
t�Q)�����W���­��~�e�ۗ�*���Y�����$��x��%�V	�@���,ˠ�0`�5�;O�E&�B����K�o���hW��^�":2���N���%OA��f��d���$|�r:AM�)���z��_DC��-�X���c�ld�����fԶ����&��x���kٟ�v@���i�� V�0;�i�V����;�à�5Rt��ӌY9ގ߁i.�3���P������Ξ�tlY�(?|���ӂz�]�����񘳒�9+́~���(�����p�X�.�K�>lO�W�R:�.��Y��X:�D^���ħr�\�} �����L��9
�}�jh�F;!��܄��M�q	1=F���(��\b�l�&잮?�ԟRևs�>�=
x�Ҝ?���BuNguF��V�O'��8m�a��X���v�T����
��(�v��J��o0бz7F:&d�r�n�gP�in�/O��2��b��T�^fc���1�#bJ���r�\+C�1��$�g+k�u�x����m0���I���5��5����(�5��%�1�KÚ�5�Ű�k8_i��K0;N��C������E���պ <H68��	)�7�Ҍ�^�p!�W0%��c��WZ{�`�m��d��d�:ɋ�o��4ͯK��ȵfo?�=�,Z�]2�4\�'!�����Z�
��:����,a]�ITw�R���^�����������Ĕmg�����mF��`N��9�[��9���� �$����i��-b=��[���a�����&�~��(����� ��D�@7�p6� =r��-��?�Db�˻���}��8 �����;�%}Byj��A��(������ɘ��p>NS
?��1�,~ὧca�Rx��;�����C���SO�T�{6'�$.�a���d��5<L!�cRZ�I�:�*����}���n�9���	����suH���b��[;��+}=���@|��Y��b�A�z���yno.����7)��=%��!�Σ۳������:(��O�Ϫ�;ڕ���"��	!�b�[��x�f����? Z���r�!JP������V$�@Z���OA�t�-ĘL(F���	���Qz���Jh��W�9��"p�D��F���*b�h��v��-�3D�E�#X0��"�X���2�K
Rx<�o�����Y��׸x���Y)�������~�T��7�I��ל��m� ��w(�f:,���q{�ٰ{+þ� V2	o��z޺��ՐP��b.#�$�q.iq�`�D#5��ݑ.����u�F��R�ז�v��}��P�=�\Y�L�1͉J.��&�7���A�s1�z~��R�!nǴ����坆��x� =4B{��%��.v������N{������1��n3�n���P��Q�[�E��7ui�n�i�ؔֈ^Mw3=����p�DW���ՠ�
/��L�?�Tσ��O��([L�/�HI�/�D��QJ�kg3� 0���������-�����D�=@���lO�
��$;�5z�;ǩ��	&���{85L��7�?�8u�2�Y):��*u>@F��6����,�����9�0�]73��&�&F*��mg�xZ�����$����j���v̤��E����ڬJݤV@yTx���_��/�����=X�?�1CZ��8J���R�Y^��˘�L�t�AC*5�=��p���n<����I͹��H.���
����5�je�Z��Z#�V�"'c+ds(��Oژr��U����gȽ���%��L�6)�����wH�d����7��<�;�˲��b�y��g���.9oR����ji�h�G��:i�N���nX���ܘ��,����MCUL�dE%:�m"��@*�rx��ܣ��k�9͍�;p����� ��C+-,g�"�kl��fC���]�]L����>'��S���_�>�`��ɂ�4���A�bb�-�Gy�_��}�

�ɓ&]hk|?����应[��pR�,�ZX�����oF�&.D�qQ���c:����tT�]�`�0��<V�V ��m��5�����IW�	�q��f��0��p%|K�}�d�fqͩ�X�3��9�0�I(Ǡ?,��I.���[L�`�W9��(�6��?�n����Q.�����H.���x\�>ʪ��֊�=��&�5���75��=�:ݕ���t��~а�ᒾĝ$gq����#Mi��9��M)����QR��3�ˑ.�7Ce%�f%���"�`�6�r���(n|�+�JbB$�܌���S"�	�|tS����p���,���]p�� ������u(N�#��f��'�=zҠ�	9k�`���׈�;u�J�'�e���>�����[4����i\���ܐ�H�]���D�U㾌E��έ��@�;��]��
�{�L�i��W��o�F��f9u��P�#�/�*æ��/��=gns����= �S<Rٷ����CBf5<�) Y���P��Ֆ�7�r���rQ��1��~���L���Ћ���U
��o���2�@7���Q{47|�(��>��4I͉�v�1�ո*|z�e�GW+����~ԛ�})ؠf�,rŸ(N�J�"�;bJ̰ .�W�]o�"' ��m E���e���(m�D{��=�>&�h���*=���4��
��S\ҕGA�Yi��TB�nI�,�������i�2��v�$6S7(3e��)J��� n
��l~��<[��eh�x���
`���D�p��l���$S,�,�$��?4e�Xb.���f���[3a��d
%fyz�<%GLi.ʡ�+R�M��uAKj��oY�`�'UY������U5���)���!}��8�������Y��t*�MB�f�+�*�����"�i��11%T�d�h�Ϗ�zFM� y��'I���1v59Sr�-1\� ������υ��`2�X�#���/�&[q�[^������Z�`�u�Y�#�3,�	�#���,~1�ˣ-[��B8C�!Z �k���B�9����8aU�a���x|�1���_��<Ņ��k���{�������ZX�	�L ����!%��$�(Q����m.!�!=�-	��>��v �Ut6|	�5It�NX��>��^��]��C�5� ���$վ��[P��Up��>��B��?Rt��#(�0.$��4�ޗ��q��@~�k;�qG?��8c���P���JZ+}��JwPP���b�`],^��������z�(wK�_�"ۥ�V\��� �BN��%I�IRl��cԩ�5���٭�	�7\ZI*ј�HK��!Xv�YT��3���"��������PV��75�p_<̂�r+49
��:����������&sB�;�����*9����1���Ǻ�žS;�f-r�R����~��F4���2�Xu6���N��8�!��}�NR�������tl���'K���R����ߍCP�Ε,�����|���� �%��>����.�ͪc_���h�p�X�j�?��b�Հ����ܲk�����sq���O����|���b�	��a>4Ea��CV�i��������3�pn@O�`�@$��%���Y.yY������i�5Q*�M�w�zka^X�U{�>|KT�ߌ��VP��GI���i��Hu
�:i�a�=�ޢ+s��l�/+���	pA��*{f�o���Zͭ�ޜ���q�%��TZ6^�������s�N�~\����G�,,��=$�aD�?.>!$\��$�����p�G	�0��#a�'���}�M$\�_�q�)C�>�M���&X�k��܂���J{KAu沁�&&(e
=] ��M�\\X���kܫ:�9�-5q�t0�$@9L�=T�#�x�pM'z�BS2E�h[�ٖX<҃�D��PY�Xn��aSv��<��
@�\O�=h��,����}ZM�5/_紵#�����h��O����~�uǶ���>#m�]�m����Bu�F(�7X[��`�YY�	�����������=yy���[���&���Nn�qK5���e���c�q|t',�/��cK��"����҆(�L�1秣Z�Җ���8�5�$(��"�w�ʛ$�[!p ���S�3�
�ei�"�T�@+�4�d���x֬�̳�E�	L�9紦9��f�"!Z�';.�뚊h�\iH��]uE�t+�wO̊D����oc��㳩yٺ�az��Q�a�>n�G]=�v��侚=��(��y�'7Kg�K?�C�u�X��Q�GĴ��A�f�]�U��֞d�/��,�����f�_Rv`k��-�1O {�0`4[��qd!g��yͣ����6]C������xO�-m���*Fۛ
Vc��n�,ֶe��[��M�}��j��L#�����u��K�M��Q�O�����ͭ'v&k�IN�����8K���2�-�w�S�i
{=??�K5Wo.|Oq��i�Q��֓iD�D�v�H���῞D#j|��{4��>�(��.�P_-��T��T֜b�ҖLC���ڜ��r���eU�[-�GQ �.�/L�QU;:�G�C����_&4O��,�&� '�eK�>f�[�p]�S�*���&���'��怸���8��P� �)*U��XBӧI�@[��ѧ	R_��=�ŋb=r��CU������&��e6|?�}(/��nkU��9g2��N��No�@ �S����n-��4S�d
�|I�, ѸGZ�-�k�R���6���!�Ԏ�q=�R_3�aj_���s9Q��(N�g2;4%tC&��ۮ!�,��ڕ��hA\݁�9f��aA7f�mL·����2�������2l�`�r��@&K�w0�HӨ"��a��]cyN�� �e�fsD'�LC����T�A�/󀅅gc�`U\�3梁�S�qnj�^�-��f���Þ�$��б��:Ü(�8�|�9z�o6���1�i�u�����?��l���q��=z�G�|s�o�]�t���S;�/���8�&��-;:�4Q��њ(�~R�Q�xh�2�l����8��ݜ�n�u�H�X8͕q�s��,��gIԱ+��ϴ#&�P���\1~�#GP�+�����EG�o�������ϝX�$����sÜ�EG&�@�c�|'m1�X/�Be%�a%C6K�-�2�\���ㅕ���"i�"#l3��,�F����Ae+-�)��G��"�nLj����ŴƝ�A�gY�Wc�x=<�svrY��H)Z<t�!��R=��5����h��4,��F[Eg	;�D;/`<�1^�1�����SS������nשa¶X�{�	9S1KC��X����Tѳ�Ц��iV���{�1{*�Y�>"��]�������9�ɯ��z�х���e~��Bey�Ȫ�΍r5`f��������%H\��R��ED�^���a��/Th�f`��2�L�RJͅ���v�2D�רjգ�k���+l�-�>1 <�θ�QrK	ShZ�hAD����ρ֪��a�];�N��u�=t��-T�S���@pGp�,m�N�G�����x"�x1Ў������'��ȡ2E��؁�J�oud��P�=}ɳ���j�l�2<��ۮM�x5��\���6��į�C�:A���R���(�W������{��[8�u�?�]Meq�yx�t����n�3�0�B������Gpw0���}C{�a֮�ɣ�}K'+�Q�"��Rvٌ��F6ө�}<�"u�˛��vԘ;���bY4+��@;M��7Qի�$�I�X�c��7�B��q�OW�	�.�e@�M�S.|u����6����ن`R��r���D~(�f��$���y!���0����В�gm���f��7��U(����\���/��|g�+�����
])'�*�x��T�g�Rv�=+���VJ�B)��+��{B7ԑ��[���f0�v�U6�FوtJ���ɲ[X���=Y�a,���{�Z��Q����zc3�����c���e�P��Uy�x�~i`��i�.���Ԧw�jWo���A?[<�9���Xf�)�g�('��\1N܇�f�	��WN��ӻ۹�F���%Թ����W:�g�j���-�d��f<�Jƪ���U$Ux~��q&� ����v�jL��#M�5�G{�<_����;��^v[�i�nfZ��GzZ�h��
}�p�y:�!��ܹ��Z_k�ztSr����M�7V<Z�C��Z�>\�I�	�@�C�V��O7��E������m(��I_��_J�߬x]*�Q��U�tv��X��ˎDH����ȹP�=�ˁ#��服÷7�p�yj����Z�Vi�̀w��].L*��.�u��(��ťa���]�XJΦ�m��1"da�}
����Xn�o=_V7G�S�딜��P|s.9����R��g�Q�� \y���\�:JֲG��]6�qg@��&R�
X�땞]�	��P����Y�Ej��b�eGI��a��ҰH�{�a����z}���7Ta�w�_�ˡ�K���
�i�o�~IOXc��d�*��Uv��x�HT�Qͫ���̘�f.��u�>�9�7M��1ATs��H]T�8�94ݢi�oifaH3[�|Hi~�Ei��
i>��4�� ������[�[����Q͙�f�Gz�S��Q'��Dym5[���@y$��2�t �ڲĢ쨼�,L���ԭ,���e�k�eymQIm�M,��NIj��[Im�^��&Mzɘ�6O�.QR۹�&���*�a�_IhcH"8l@X������*y#��.����v�:��&�ل*<�X����MIm�*�m �5i[���R�b.��J&PP���֨_�u��M4��:�|0�Ir y�v �rx�t�GE�蹽�_C���z�����2�����ʑ�q�0t}(+�3��CY��w�y�ݜb��p��I%8�1e .
�MC�
'T���� ��I�o�z�P]+T�CeuB�
)�]6�T|�Gj鯟�����w-�]ǣ7'�2멧�
����ۨiK��ߗ�]��>)KM+�u�ы�;��DQ��dQ�#��9���w�-B&�%ZBk��]㽆�{d�K?��qH�]��}x�f�V�\Ȕf܉���u�2�g:y��M
�5��=`���^��R�S��dQ�2�.�ŭ��qA����x
�M�-X[��L��C5Ώ�=�<\�V�L�B������H�$��T���KJ$��u��֠?��3�L���X|Nk�G���hcĸ�Ԯ���ʸ6	B�/[��;�^�Τ^Tx��p���u,լ���Ez�5NMMO[���ۊ� �'i����y@��:�җR�ۜ�LO
�'�F�n��<bV"�R�������V�J��w����@��/b�u���oث��!�SQ�e��z���Y/��gI�`\`���[��$�xmy�҈�&u~�Q���V�d�҉���Q%X���{R�o+��D��#��	�����u"i���f;<�^J�LR/���6&*�t��8�N�U�i���&C���RFl��!��4
�6���cdܔ��u%�u��^��j�׊i�͎v����FT�8P��ѡ��=���V�q��y���#)���Hc6+zͺ�3�%_(�~]���[��!�I��ͺR���l7�J�~��^���iƦVz��h��)�ɓ�����Ziß9.�PkUϸ����1��v������j)TQ=5��s�:"}�.��>�|�)���w)�>�1�J��i��hI��L����H�/b��<���T�횉�4�՛�n'���%}��v�WlOk��nr?�V�R�Zk�..�-b�%�s��_D台��ohB8�^/��L)�]�Ґ�Lia�Њ�0X��v��m�'D�]�FcO� BzX���8C��+�	=I=�5`��.X�K�����O@OX`�zݴ�u��R���6��v�K%�O����	x�Q�Wh���4��)A�8��UtHtL5p�(C9Y��q�e�be��c&���$�~O�ъ�j�Nŕ �7�R}����C���BY�X�"�x�}��Ư�`���Lw�+�����K�٦,��4^G�^��Z�Q�x�ҭ���Z��ɂ@{ ��a��B�"7Rx)�aa~S� G<��Z��ۘ����7����xr����f�k�7s��j����ѠX�;�2)n79i.�;Џ�q��2����h�?� o�`_��+�t�+�����'7-�Z��fdVP�%�%�zX9"����`��cH�4S���2�8��<޽�Qz��wl_Lڐr�M[�֣��7����7�#�l.�Î��@�-�
���f�5��1k�Je��z*�{?W�_��.E���Y�}�s5T�4���UB�^��@iZ�l��w��^0�Z�p��)eN���VCŢP��Π"�X.%��Q��-�г���	�n���%�`L�-�*�T�v�sIO�й��UF��i����!�����z$����q3��߲��
�?�ڡMu�8Z��GmZE7������4�RB5��~K��J�VN���e��@�����vi̻������HgS��o���唤V!F����\���Z ؞�O��_�#hth�k�tڧR���~
�F iFM�(�ʩ��A^�4W%��ʱ?oR����,ַ����'�C
�����:؊/6)��
�ң�C�2ȕ��$�,���g��o�ګo�R�'�������eU�2����� q�4�y�0m�с.*}�2���&sq��jB��П0���3��`�m$I�iwh\�
%p�q+�o����]�hi�3�%m�l�de��i`g�^ٽN1&��a��(�x�z3�x�2��ކ_�7j
Ay7ֽH��ܓ��˪D��=TZ9�<�6Y�н�>C�0ni	@.���_�5���gtx�i�$ � �NoҼ6���T@y|�@��Ť�w��oo) c5�m��������)��5�)�0g��.�٩�(s��ٶq~'ӗ;�1}����E���%Ź�Kua���
ё
$���J�3E-b�G^fGD��������K�L3�_.߀��6�J0_.�N3_,RŽx
X��I��N��s�a���������F��=����5��XE�cĆQ�H�p��"^MږF��M������d�'��	���n��R͠XH�|A�W�6����U*�ނ"A*�_@j6e��Y�1pi��G+:�0k��Ͻ��y�F��H��%03�*���q��Ќ��F~�tQ/N�R�b�7[�ڸ֯��A9�B.W%;��p�-S�d@�F��6y���#:d ��u�.��~m��*�.��	�p��A}4f�9l��f�T.X��_^�ֈo^���WZ�;論�~�����Q*�|m�f�Z�����uAZ�@�� �A�T����נ\�"[A�@q����������OR���@�W���>Ҍt�����_Tuu�l>�O�	LV�t�Ǭ�r�E �w�.Mz��d�E��q���j\1�j
h��ǳңCѕ��G܄�.^$���Eg�,���t{���q�quhO'����T*�a�Y͹Y}��阢�yf�����d������Z����Be��1�PzPZ�i+sYRGZc��2���P=�1I�7(���4_r Q+������t0T�8�юH��ǁ����,ә/8���<���݋	&(�C�w\��~�w�.}�����|��x|C��^Cm �{�HxJ����搟A;}�OP���B��,���W8�2�8�3�����;���$�P�g ���T��c(�G;������ك���gXX�Ut��3�Z�������/o�ׄz���H���ǔ�4X^ʹ�0���竨���gƛ��v���.�#�%���nv�q	T_��TՈ�.����t@ڰ�ช�<���/>J�1��?��t�Zo�Z/2�\�]��T:(�^C©�A��$V폓#-N2�3,�I�dQN��~'�a�9��/?ׅ��/�}�N��i�f&�9d{=��<J�Dҋ>&�p�A�v�A�Ф\54:�Й��W����P�gx(|�ǻ.O���{#�ZJ�ǚ����E�g�K�h'�ʂ���{��	�Ki�z�lLn��0�"^/�(��r1xj,��GHo�D�x�k�������S�0��vb:�<�����7�'6���V.}�7GIL�g��Q�`L�F.����3�Kк�Տ�+h�N����<!JoD��>JEa��`�Ք`/͗j���ae/DMu����0	�%��7���kѨ��Rl�0��q�mFDoiP4t֮�XG=�!S�q�J:��%�f��^�Lʂ1���
�m.����b�E<݃�\r�8�5đו�t�{��=�x�d����Fa���t�rVAe��?��E}n�(��(��;�M� ]��b�'���L�
��e�bY:��@��56ՙ�r��<�"�l���M�r`�8�\0ی-(H�/��lo�k;L���i	j|�b�F�q[l�����k�%���������P��������L�|��Cp���X����C`Ԭ�+�CpZn=���P�+����Cpv���km|�E��y��D塇���)�#1H}�Hb<E�!�B]�9�%��V��wW�n�+<o#����/���*�lk�f��8"V��8��D���b;��h��r[T�7��O�4�?]��_�:�	��;�+;߿3��I&E�5�#��,OV��i��c�3��"Na�=��<���8�|��9�VS��+�E0c����_Usl#NaJFK�^5zx�֗� ;x������5^j�=t/�nS��	�[�~�2"O����ʮ��5�r���;,�D�I +����u%����YQ5�j��PTPf�|vK���׮��9}U��_ѭ��~>���<�6����,s��8���[�aM��=�7 ��mI��wa�v�i���n��T,T�V�=����1c۔�C�4d����ۮ!pFx��MK�TL6�'L���E�J�P}�P(&)<jt�<��w�V�~����7������H%�c�3�a_G��G�S�w��P�����ҥ��l����՚V=���V��<$ս�DH��;�*,80�����5J�̧��d!�6�ԝ�^K_���W���Q'��F�~u��$8sisT��s8zM��fgm��%�-%�ޡ+[�,W��Rt�2��c'YL'`��^n��uD�} 2��U���9y��-�p0��G?���<�mq�-ؔ)�T^�z�w����g�B%�,,�4e[�~���9+W2��pK�o���۔se��t<�R�����j�EBR�SFީ��R�n�8a<�W:_E�A�ˤ,�������VCu�߉Hi��n0��kf	3RcC����^�E�c�y�������趓]�B�w��u����t�+t���F��ꮟ�]_�+��]_�������R@<�������Fl)�����Z����~�
7�F��FD�cLm�������wЛY(�(-�J�Ev�xc�����`��x�x�4aM%�5�ͳS���G�	�0' ���2G=�\�D3����s�Ѻ_�o��=��PP{	�-�SW�P]U`��$V����4�m/$:���v�ဤ�<#_�Ɓ8C¶�fܲ��lp��C�3�b��b�/�;��-u��'�5��-,9 ��z�O��7�s��Ѽ^f��.� HmZ��[�����-ʔ�R3r��b
�Jg>/��uM=ǒ�4��Z����v}a����:���=_�d_-�S*1*���̘�2�T��>�U�>O�R[��~j�U5ipE�:���L'��yBa�-�����Hs��Y����5xWH�`ګ0�,�6����[ܟg�b��@u�G�L8�#�	�Vf�]Z���,1_Ȕ^8�� ����ml�R�O�i�(C�*B�����_��ۀa�)�X3�i4Ę���Ļٛ�G{��@�B�b���Q����e������B*(��.Y1i:�_�q\�ۈT��2 	���0oa3����C��;G0�r2�-g����ס�v?9�����HNr�~�fiؾ��@�l�Uq�C��	_'q\Z#�C�]{c[)�zoe��!kp�N��!���!�R�T�s?t����i�Jŏ+�\�N�-�xB���M*סo�>�o-�nr���ߥ�� ��*J��b�c�=l#oR�!?=F���r�/[�.�u	ہ;�,�+Z�ΰVxͤ��Ʀ�t��d�q���ae���BӇ̧F���ѱ�tR��d�'���/[Ύ�W��N+JEy��Q�^�*y��ѯq����l��"��&`���=o�ݬ�>��ޭ��YZכ�h6=�	��'���j9���a�}y@5W�șYجI"=)/w��g<j��^[9��+}f�|�vF����*zᗰ�z
�R��H[��4�lg[j0Q�S�r���	N@�������7U^�'mh�� Q�-�ZBk@��R�bJ$A���UH�)-Դ����n��������{u
�(�(�u~�`��aZ�+EJ��������$�x_�$�>�y��s����kȃs����v�2�{X��|�w������VJ����/��
��)��k �5ǧ�Uhp��yڏ<��?��d����Z^'�TV9��]�9t�(�y�[���s�HTY����H�vN�ӘK�.�1�].�W��1'��uO��L�Oe8R{���ץ<3J\�9����9����H��,�~�
r1�������~�L1�0 )�>5o5J��s���2}����Ŭ�*M���o��n"aOrUZD��:(�96��W�O��n(���҆9�π�����NV�ǝ��{��85x�̆X�p�|�1C*�b&5�ST/�����BsB�O�T��� PjԒ`h��;Aܳ5R�J��gM��;n�C)x;�)v�|;���N���st�����(A��z	1�~y�
�`\�:f���(i�P(�6ϡ��#w �����S؉K+�OK��d�[F���YA'0���>�|�Ku#���.�Ų�=y��1h�.����a��U�-��lj!� �~ٛ�QfL4��	3�b����јb]9`:LP ���-dP8E���{00�,��Ĉ�*�*���Z0:���7!�X2��%�J<D��~L�H���čX%{o��d�41j��m���ڛ�ᯇڲ7/D���B�{��.�**[�ȮPي�`�p-�Uge��u�S��Q`T 5��� �)W��EmFX�9�oő����,g��<ظ��->�E�u#�Ǝjt���L3����޾��/\ݷ�1�������Exh��$ѡ��H^��$"b�=�o��!��N�[��p H��YY_���(�u�����AI:r'vJ54�
�Є�_�<�����=�|�'}
^�tK�d��?`mfN����лX�tFeπ���̨�,'���A��I(:�l�6�A�)[�m]b��le4߇t���p�J,��*�?#	���ڝ|���,.�����%c�ЇWb�C~���H��FIՅ~�m���ꨰ���u�9�Z]͝�áa�����?d���3������4D�����L�PI������K�nܚ�V$C/��~�r�i#"<9�^�aM��]�E>�шjP���S5'&���9x���C�ɞ�"̣������'��������{���do��h�����Nw�F&���B3S��mz�����κIl;��C�O~:P���URF���Z���j�o��f2�sH��U>��[䧀Zί�l��FU�E�`.~��t�O��pN�t0������KuN�����~'ŕ�&0x���e7����a� ��R�|9�;5P��"���w�C�j F$|�����ؓ��h���!r��4�7�S�}�;���?T�A��u�h���̞���.ѥ�"9��7&R �س�YL��]��v ��\�,ۯ�'�Yz�<�I4K/I������o����6���Tt�:�vpep�*Hg��������TJ�	:�ܵ�#vںz�	���U��G�4۝W%���/�\���4��z�^NK�ɷ?�I,���D�\���rN�(�kJ���M^�#p�U����+N��2zN��,��8���tYV�̳j�9��im�d^��,-�����Z��������G��d��$;v�&Ku����N�x�+p �.F�����lXb�]�}U��*6�U4�N����Ke�]a;u�(�j�>*��T9ݰ�EE�<��3��+�=�(�Ȑc��uJ�ǣ��Xʉ��� �ߏ��#9۾���ZQH�y���Dچ��h��UL2XD+B_Y:;�o��f�z'&��n�����H/��_�}`�yN�G�$&���g(�^~�rY3%t�o����d��1܉1rM�8�x�[�����\O�آ_ڌ����DD��-å ���PP����l�'}��^�*mx	I���>D�&����۰�_~�F�Ɗ����_E��"�HR�UA���>�,D:�m��T��f�n�bw���ߥ�
�|�li������d^���Xʔ��~���0C��=��@�X)��ʙ�_as�Xs���c�?���?����R��SM��QY�Gp�0qc��� -���%NÑ���VYAi���M���"�r��,����č�lpK|U�x��ru�V��Y��a�0H�����P$w���ξ��gߺ����"2��"⮈ӑ��x���y�x���p@.|�Xg�h_�%����A7�l����R�;�%u�d��{U��j=�j.�jzE�,��њ�vm�__���{�b���fR8$P/�0؇�Ϯ��N�1{ר�|��Y���"R��?����eI�ؓ�3u��
�ap������DDB���1:��S�H4Q�`YU�S����Sb�'��)�LO�e�!x=�Sd�R\��Q�̂��Q,�6T�j�q���KϤz3bmg���@F�~0l�q*��-'�_Mut(�Ϊ�:x�X�)C�V]�Lس�2�,������ݒ������S�6��.��1��I��ҎT�p��і �9��X�B~���`�\��?�!�vpԒ%mD�+�m���G�{����`b��UcL��m�� GqD7*x�F��.��c8��}ȯ�01�����R���p$I�79�S���ȏѯ��S�+��P]�Z�"�����G��$�J���'l�;@����� 0ǃ=u��0�q
�ŲfI�`�{!]����6�o[6Ȉ6`\��ZO��*?@s�L��|�;ȸ\�{D��JNQ����|iO*�J��gtc��t�n�s0bJx�".��gogx֒���m���U�Y�P"�={��Y->�5�ߩ��8�`A��qn6��%'S�ϊ���gy�l��ɱ��Ԥ�uA���[i�V��@��õ�6�(XK�
C�*�>P�?�����T�#�!M�ԕr�c�-���������'ݢ�i��bx��n2��0~���1{�3��{%�`J��/(f�C�7�/Wy������;�����m�ٵ,l
�C����e���Σ2��JO7�e4�N�H�@��ːG*v�hOR���Ph�u���mN�,d�(��%�m�2�@�5�ʘ�az�a �DVd�>��X�6"��n����{�	��x����L�(#O�Y�"$�|�CJ����I'>s[F�9^�!���
�(�Q&[�~�R:;8T��I��=�K6��/�;��m�� Ӫ���������>!��"3�=_��,߬�a`hJ�1�ds�@�,D�!��>��$�8�6�q�S4����D�+�s����D�w��(���b�ÑӛW���l{'�Z��g��Ў��I�خI\���e��),������V��?l����?����|Z'_��X�)��dI81C|0D�ޗn���FZ�[[3~]7D����r���P�[tj�͵�iE�
=t�S&�2�*����ay�C�㎢l޲>�|����g�{�'�"+�'ڼ%K�,����2��*Vs�E�m�?��IsLg�vT�E�[b�純��(OU����UiN��-�r#s(�r;	�S�cS��I:�ѭa�I���>�5�n#���������p�f&I���,@�(W����V[{4ty��6�]�5�u�˚޻�RÃ��x���[>ZoU�9~��c O���L���+�k�
 0L�ao�g��/�L�?3	��m��1|nwC6�/[ _���X��Z��5Q���la�jX�X����T����5ͧ����6St�s;�b�,�P18C�l�xMt��6L�@?��xH�슾���Ű)C���AEО��L�x5n۶ѭ��ȻAi�`�O��ob��ץ�2INܫ(����v]�׮0�n4@���Cq � L���x.o�������*�[+no��Z>��cI�&�?(XW�K��x��3�0���n�'`]�^�)b�B���J+����"�P�}߈�� sF���!3���Q��#Q�+Ȓu�>�X*���S���_�ĞB�S�)��n�Qn��H0S���D��=��)\�%��jb?��'L�&r�E����R�������=�b������� �4 p�� �cI����|k J^-�L#E�˂b�p5�^�rb7[M�\u�ܢ���<=m�D��,���E�2�#���
�X�N�EXa5 M�f�,�L|�&� 61���/������U���h����=�NC�`��i��4���c���%��sV�l�+�Noh��/+�t��h^���΍ْ[Ѽ�?$1��m�)�=�(/(u+:��l��1V_nP앐b�J_�Tb2��2��{�bO Y�+�t/�͊���Ά�K��`ِ`��B�g#�0�����:s�\�K�,���L4U�AI�
��k�����y�<j]
�ֈ��j�����ެ��@G7g �}�N��{�M>���[a�� �X�)R6-�bi<�����2\sJt:�_���t����Éot��E�m�l��4�^��P�����?��ݨ�J\��[��.K��.:�-x���g�Q���N�A�!�F*�d3�<�������סHN�d[@ҳQ�S���U�{��|(H�c-�i��K��mpܛ��f���+�y$�L���o��wĜd_3Q�6��bb)����jMf�@�M~q/vP��6m���!�B�J�[H��E@���{��vaw�Cc;�N�mDesB�F��E��_� �w��lҿ?c�+�;����){d�4ݩ�(�� �y4M��Z�ȽKeg%��_�G�(Jw�C�����r�^�@�]�l���2�&	]<݋T��]Bd���|#����h��6*��(j�xLt[G��z����{Y������j^E���4'��!^>���+�+fl�uq���@�,���=�-V���PqH@��O~6�st{@�7��u�T�؉L���'��b�5�g�Pw��rS&�Gd��8�#3i����2��0���h�`��r�Ku
�R�[\Bu���A)�y�z�㥍d�?B�L&s�Q�/�n���)�E)(`�\q�K�2��5���h��u���>>�}��:�ao�Y��c����Q{5����,�(��H����e^�>2iy	4���ߡxx�M�g������h��4�F��zk�BWK&�kܬ��E��BU�Ң�����Bo5�hV#��o7�zbr�Ī�L�^�Pu�Q�B����� ���>G�B�����XY3]��i��!j+7�'��qPq$f���:_p�O�$�<��Ѻ�:�\�B����Jf�.�q"���K �޳;����Ɏ�K+�K{k��V/��vҬ�F{�ʼ�(]�/�������X�9:L|��J�(y��XOV�JH���:�S��E�b`�m�Z��CU
�f��*U���:���c>[���k��� �&����?jn�]�g�h<ڵ�Fj�;��v�a���� w�P�jr'���x;���fj�C��3ēB�[�8�Lэ�In�ƍ<���c�*�*��2��Iz����NE� ����YFÑ;tM,�&C{K�%�Dg8�<4���+{��<Ȋ�N��d1F�)P�
PK'��M�y��C�ɓ�A���9�;�/�v�2��D'�®R�ny� �ֵ�܇�'.Μj�*_��)�߅Ǔ2Be��XTE���%��E��R�o�+�׊ŵ�+���rȯ�j=+��v �coY�a�3���;D���cmFh�ݒ�D~��#aD!�Ʀ��Pwy��I8֩�X�%Q����������}�Nɘ%-UE-
x��ۅ��B}��!?�3�;�0h��˛ZU�t�[`\�ן�{:9S����2QTDqHe�Ы ��k����D	"��Rޒt��_jP�����%��R\�n�ԩ�G�4���5���SJ�]��h��펵�a%?lI��3�Y��<�����.O���Z�&5��SK�����hmUj�3�4�E�~38����Q��m��$������a�f���K&�< 7�7�C��ZQ��?aoQ�lt'tR����O��c�Vʲ7�'C��f|̝��ߺ�boz]?�*ގغ"����N��8� a�/䑴��EH�f�5E\���\��HgJA���nً3ܲ�\l����ow�F`�3��чD�y���n�&eM�H%���NT�Fn@/˿����å��n<�3ArozwG�p��&�P��l���{�o7����m��=N���������k_��k�5������d���m�#b����	�:���u����
����GJ���=|�N���!wVs$�Oָ"y3c<
�O�2XN�N��Ό:V���*��~�q���������J���B��48���bk���b!��p*�<��60�8�v��x&�d�y(A>����7*ھ�h�RÄD���O�y�bZ�����$Z$��Sc���N:���l�D۲�A��u�]�<��a�~Q�]� �+;B|+�\��32�{K�bk��p��
ĲBс�)\m,#�B�*)u.uɿ\����XڛhD$Bؤl�YU�`a8|��L�"J�l(T��S��<�v;�~aJ˟e�Q�����XI.��R�YTg��w��j1D���v���-�y�����-��}܅SԻp�mj���n5����%�ѵ}��j+0h<��Lh;�ŸA���1��iwV����g9NN{�arO�w���f���P豁��/�π�LI� ���zZ�J[�Q�� ���\��[��@&�x1�VC�\$'A��ս��i����C���t��U���:A���l;�=,�s��x˖S�*�&��tt�sQ�Y�l���	*�
L��":�p�ޅ�3q�a�)5��\�3%��0տ���n�ߞ����L�N8�ջ¾��Y�q�v��xbO�_m0�;S�b����l����Jq⃕�9:!��S�1�|��������|��S0�*�Se�|���;*z����[���J��^92�����M�g&z�����da��[���x�^��{��G�f<��ݷ���7Ӎ�r+K,�z��	k��Y}��r];�5�[�x�$y6���n����!}Xŧ�F٫�lR3��/��R��&d�z���.�r��NP���ʹ��P�b ��)p��~�
QOB��U��[��U�0,{׽j�+2u�2hQ5��h*v����L���� U��ۼ�#���$%�E�(
�홀���V�+�@��K�;��<�%��r�G�ą4����0���o&�Q������"�����ѷ�6"fJ��z;�o�z��<��;��S��3�k�[�����TVM��j[�J8�c��.Q|'}�a�x l��c0�Vg����K51�b�L�6�wO�+�ٍgd��L��Lҏ���/��j���w���mrՑ����*r�1�����X�����Q/";Fu>cu�O��D ��HϷ���aȌ�Gi��1���u&��b�'ov&��B�w�1u:���uߛt���#K�,o
L)�7����B:����ƛj�GwSmX���M��l*m��u�PaUʹy�A��ꐠ�v����Y�~_�@J
��Y�jX���t�|��q�eN��m[rדF�̂J��	��B_�:�iT�
Ӝ�u&5fq��Sx��bO!��M��p؅րA@��L����f,&l&b`�4L�X����[��ܞ�}'Xȟf�4���n�����f��#%�OP|��νQ�?z����)l�,݋� |�͗k2�
�v�{��-l�G:�6�1�P����oc�G,�É��z�v����zU��Lb���Є���������A��5�k���(j:�gj��W �b�ж�d��d��6�n^�6���p.�( ۉ�%;�|�E(LqK�Sp�/tw���3��<�f�pR���W|q�.�w�L�&v�,==S{����b�� �ȫnʀ,�iJ��;���G}?9��5()j����nC��h�z.�ĥ�a��߽�V�S��_h4JĔ��	��r=;���'��U'�Z� ���xi'.�X[����9/�<����ej�XaԐM�7G��dN����+��2`����Q��X����2~�ǰ,J'P�5��O�kC~w-�G��FL�r�n?�D8ӝQ[��F�)���y���K{�o�$�,��L��x�{U�G�4`�O#�~�=�ٻ<%�4T�^iι���X��&͘z�'>�R���\�C�<Ʃ&W��	5K6���-�<�v�>2��[E���-K�2M���_1Q�K��a>q?�&�,'�y���AM7�-���N)�ZD0�]����QU�='khb*5�˧~�/慯����^*�C��J�W��b�&F�B�{Mud6��a���ҶHU���G��{�;������Y/�C��,]m2�*�p�ɈA��d�d޻�[]6>��ȍ4"?j���q�H<�x������aa6|�P}8'1���d�	Ȧf!�I�۽O�����-(�%I{�O�ՀC>�?3�5���^�gf9)��)������/[��o3�cG��ϰ^tJ���u3����l�k��bRVY�U������˪Lʏ��.���Ӱ
������L��H����u�D�h��d�v��;Ӳj=עvg7���;8��BT�Q���>�j>�V�*�vC���Ќ��28ܝdM�C�b�|���-y�)rA@��#�Ҋa��C0���*�TS���E;`�w���kKs"��˯�vB���Cu�Aϋ~��쭱�UZ'��!S"yG������ֈ_9S�$ze� ��b�,�]c�,ĬK�C'��^h��s�|e�Ӕ�H{�H?X�D�2�'��>�A��:���;䧓N�d�0l	�7>�s��������h2�<s�V��`���i��|\�������[<�b..��3DP�	me�*�5p��#g��6���{?l�l��ƛL��ib�ː=%δ�1���˭���7�f�L�v{����|��i?}�ٛ�B�k�x����>L���z���	8�����iP@�kQS�"'觵���
\��(��ýϳ;���ᆁE�/�}�,���Q�D_|��oe.a������}��N�f@������"%:#�م�u��Y8��U�r���]�ś�WlYv�	A.˞a�c����p6�����n
���R��z�K�%}uJ{o���'H�4ԩ��9�y[�U�[	��$Rk���w�&[H���N�"V�s���ۇ�m�Xy>���1�VAߎ·mޮ��a޽0>�ep/�h�"R$�"�Jk�-�����3b}<!E.�Ȟ��)R7�Ay󶦕}���ms\���n�ć� QyU�{��9�;� �T�UL�:��h���f��h�%p�P���ފr�d	ŋ]���_�0o<�6Ǡ�#d�>���k~�f`�MxG?�����h}�3OM����Tj�<C�K̥���i|��i|)Orw(<�jk���.<��)LJgo�Fm�����%��B�SԀO�8"�qx?�N6����
nR��$8�ߡqY36�� ��2����p����]�^�xQ܂ �;W������,���.���5�5�^��כL7ވ�a{[-n	��f&��C�e7��(47��i�~C�qR}�g&�`?�����Rǔ"�$%�ڢ�*��QQ��Uf����)j�@Mڌ��?�:�E��×�k��-�7q7�����/��l��J����h$\j?����X ���	�A�
4�7�����d㐚�"H�~��M�5�u�)ut�4�p�'b�V��P���8�����]G��N����ĺ�ڛ1��\w������h*{3�#��Fp��ތ#I[}��j�t>����$�S���2u�+��7���-vI�$�/q�9\C�=C���vb�J�ٛf��{���q7���a[Y/��~�Klg_jHV���X\*����7|xƠ�4��K�Q<�X�� 3�rEt�pME<�~fƩ0_ ��6�qS�Q��.���{���ǂ"RO��w>�;�ܘ���l��+�5]	E�u+�k�Oz
OLd��Y�׳1���0El|���|�5�������͗���b@��,��ǹ-Hcc����((H�g������_c��,�w{�&��
|r"�e@�K�2L�.�6��e�#�����Y W3�|��m���/��[-Dl���0c��T�_b�ᙩ	���p~;��fj�q��Y��&i4��� ��G�0�*/���TƘuIz��n�N� �W���j�|�We�9���u �&ތ=�]�1bL�Hy��*n܂�Ց�UC�HV�D����=�\�&���M�3-0&
��eڢ�űM<�Y���eo���r���|j� ���A^{���N��=lc�[�^��K���ΧA��j\2�W���c�=�#����ӝJ.#x�r8�/��n��J��*���1���K�wFFD�[|�l'�=��_�\S��e��]��|�w����G������I�0�ݿ4k��({͙�G60N�5���� O�`��� �4 6
hX��xt��x�^�kori���7V�;I�#���sށ	^�oC�N���q����R��|T[�����Z7NW�Z
�E��
f�WU��iM}6�P��
My��qs��~¸,�.E92п�>���9�I�,4��M�{Q����2���G���q|����]$�ӊ���z�>�Ij�w�T�����B	�3C����@0<�FLg{����hv
�#��2��Yl�¬�B��=&x10s��/\����u����?c����R�W+�k={��Y�ro?����0X�ˡyK��4��S�j����k�8y� �M��m�f�L��2R	�|R���?a(_�=<kJzO����d9(~�T���4����#��UZ���cw��#�t�%뮒*�Ȁ�!`Lf.�l�̡�R�����H6qy���-���cxyWYCOSy����&ҫ�OC�ľI�����*����U�:��#�F0�NWQ�8�)]g������0��wV����_����i/z	����N��K�>@-#�=-�%�3��ra���8��b��>�{�"��1Y ЩIټ�ͯ�o��U�mó0��B����֕z�%T��0��
�4h�"�ǢQ<�3*�+,�}�,���-+C��T�^�v빱i!��Z�(bGP
�x�:W:?u�&%Z�E)�gp���2!)P0/�Xo 
5#	�U1<~Ƭ�(�z�7_h(������A�=	�h^hso 6k 6�"�3�:	b�����X���"O^�A��OH�(�z�7N�`��@��o�@L�3�0�3�P�4b)�T%�BO�@��_h �'W�N���y�gt��fCڪ>���vnb���,zVW/cڞ:�5�)-�_����U��ƺ���{������ٜdw�Щ�83��"���@�f���#R�a��V�{���;H�65.��B�^]��w81۱fl�J�������:j���}��Y\�ڱel'��k�v�>�x�Nj�����>��L�hjǑ��F};��0��R��\����������};6��,j'D��qs��p�#?������f];Ok������ڹ*��w;�� 1�qelg����Z;WR;ۼ�Τ�������1j�0c;_�t�|��wL�ߨ���˦>۹Zmg�S����z��G�H��lObA:`5u{UP�wLF��3A�!�����C3����P��`5�Yo6K����oq�� ���:������{��G����W!}$~/?<�<p�ʝN@F���fgr�K�ч�k&E��W�P5v:됿Zt�,�^�x(��>�W�`���'m��s`;�׹� ���D� ƜLZ�E��986�P*4�BCe$/&%B�d��Lh�!?:��[�iь_��l�ˍH25"�F*�A>S3��x�]�Of�'��%�w	�=���������x�{����概��w����~p�i<�i�������hq����@y]@��(_���&F���竤ץd�n;��u��vA�F�� y$A�󅜳h�
������ ٙH�X�,�<w��@�0�(�):k0%�B�uL��`^��`F�`�9������B��`Z���G���^I�����%cTXu�j�Ur�]R�p�ԱL1����s�
��`�SL��V������[�w����,�e!Lq�����{�3c
n(�����̥H���<y�9+�0�j�����:V�W.E�7�E�M��u�ة��{*���g���`�uz��q��^�B��q�a��C���Ҫ�hN[.�:�M��]O��,�2k���qwgF��g<�@'��G��$4v+���&L�SZo�7MBn`��O���=ܼɟ.�F'�SQ��C=9
=�m��s��m�8�d�*MA����	SJ뻣��ym�Y����,�d+ l�E��/(���f����	��2�C!q��,���K�DH,�a0ə���3���h�2�"�[���B������ǫ���6i�&�����,u�H�q� 
����#�2Ț(�޼]�>F	���~�!�o�S��	糁
9�V>P��K�ZC)�œX.��9$,��.�֏�/=�FMb��@�1iI��J[p��܊P�]�}B}�P�%�G#��n3���󤁐e���<w%�R�1�h_hO�	��X:z�n�U��P�D�|�?p%��#K�cb��>��_��\et7�H&�!���L�vx�]+�E�BڮD���^$C
�ӫS�!��UiJ�L������W0O���� ]�'$MD�O�yNt?\�=� ����C�o*�\�O����d��_�9�^d�`�R��P	Lo�p����@{���aOA@�/���"z��&�$x��[�Z�[�L�2�$��W�e��x�b�<}��r�x}���8�M�Q�ӌ���GR�x�(\Ja/
}�Wj}1�� |��f �`���E��p��Ҥ�?^��{�6�L�@s���L��Z� �R��`�ګ\Z��pt3Q�ZR�c���:���j��A�դE3�\��m�;�k�pg�Q����]����Lm/Tډ��f����B19� ��U���%��s�&̟�ąi�f���2�{Jv/�i�A��sq����w��:J% �R��=�LjK)ѝt�l�$F!D�9�!�=�Wv�.�=n��U�e,U��j2{0Y��]��eF�`��J��qNǿ'��ݢ1�ݔ�N�L/r���,�A94��K�jȬs,e��? \!?�y��-"�U=��#��G$�N�؀TT��`���O��/h�be�>z�X�#�Ps��U�75�i�)�͟���a{�h��ɿ��@j���d%$&��ǌ�q'�����?E����JL�@v��BRQ��5T�K0��؞B"��4>�Cxh���5̐�%�pn K�՞7��a0�������]�����$Y�"mfz1�^��х�OwF9��l���X��M�z��L���;zm0��z��%sq�հ�>�eü#)R�yT~N0�5����,����X���}y!�wC�j��5b��T��f���Os���s�ğ�Q	��,��4xh�^_w��P����^O�&�~N�NE�� h1~�P,�+Fw��#�����ﰝ�PN@�)ѓ!m��|����� U�S�=������&0�'o[5BV����jW�������m�j�y��5v4`�gd��bܴEU���@��f�MF��xH�����9���kCu�0��r�
C�M�>}�Ri����'��Κu�64|r o���K)K(�1���
M�gI�P�k`�U|`�yb0�gT��{���|��߄M�#W�6��fݫ����-k/�y��Sz��M�oE�Za@b0t�'z�Q��&(�����?�M@�,]d�R%��I	a�x�#�-SQ�)ɧ�EN:�E&t�x_nk�߸<SܪL$M�_3HQv ��mາVf�GU���t�W����=��|�T>��4^�a4��ʜ�; �)~7q��03� Y��y�Wq��K2�m)��_3ʯ�)�{��^5�I:�7J�8�jA�氍����Uc�[̃��L�N�Zʶ�Y�L���2>�K5����L��d�T�ˏ
�	 ?�-��nvt�S�Cǐ���u�&�a5�[R��Oz�Vȋ���Z(���؋��	�ª�V��7'�6��� ��<7ǀV�O�jŏ��ڮ�G�yuh��K�B�T�S&M8Z��*����t#���y:T�fn�G�j>�?.�ݪW'o�@��y>��%���-�j�S-��G�(Z �ZQ�� 6�[�i�/�iO�9$�&f&���&�by�ְ���,�^\����I]��+a�*v bmbnF���Y��̝4�!?��o�u�G~^�|jB3T����n�P;M@Dkb�s�[�F�����5��4�%5�M@e��hJGS��"���Q� �F^�S�p*�x6۰�a��7�=�w�^w���y��K���#j�#����n���}��t���\�_����U#���i[��#����m�2?m�k��mI�ʩ����mKә��-�ʼ-2mKf�JA���t���i��y���i����{9�?���?���Y��@}�o��D��MJ%�&=r�~����M*�&�rTۡ̐T���)��Μ�O1͟P���0�n��#�Kژ��_�-&�/�?��Toe��E)�[Px��Wg�nؖ�4>���6*SG� fI?4p꒦9YU4��^�.:Lb{�b��m$o)�lӂm��ԫf!ɺ2����䙻����]��8s{��g��������3G5��[b�g���S�s�ty[��ӑ	~�7V���|U��0��t��^���Y�`O�52`fl��sz�L��k�4�+���	����ƞE� �XO�ɁY.i���N�� 3Rp�n���r���R#B,uDG�
��/c{��yJ�<����sPL�S��.�j�����-��p=l<�K��H>e�Ō��Vj���f��n�����W�" pa�9Ӈ�@K�0�����U�^-͕q��m��i,Ck��p��a����س6�R��5�SO#n����A��ro�"�h���Y
��y�0��Y-,w<��2`���и��Vs/C#�&����@Ov�(�N��s�`8�\oί6cDFas!�Eq�^Q���a�O)��p_�,�M>%�!���˩ߵ�e�L�#j�ī�@�P���caf^1!
CG���� :a�|jI>���{0�w}.�]�jҧ�!/�-4�68��Y���O3@}[��P��Յ;mG�Ȁ��\3�.�}8��Gl�͢It��`��
_�� ��eC�>�{[·��z�>����<��O>W[~��5����[���-��V<��M)��͠�7\�}��I��uBr��s�:���_C�����������P�3�T�3�/C9BN���D��)Vb^5�a�"���?�[���[.ȮaQ���Ty1�[Q�1]�X�i��Z_M�s&����J�׶�^��=�L���V"�/X�����0�/aGa��~e��	�h��~����ap�W���5߹�j���vw&.g�3p�������(;QT�!u)��[CW���%Z/����3{y-�Gee���1��� �F.��Cld���
���紞rꏺ��6}O��M� Y2���D�a��p��)�v�q�s�i�i�$��q����,����M�q�9��w��̿���Dδ����ˤ��*ʤko��ԋ��!��;r���VM6��d��Ť�s���N�����[%_׉�#`2Eu��֦H��<E�A��5�9j�a� �~;J���~��4=�2lm��	B`.s�I�:�~JZm�97r����/j	�1\�b��=
�,Ĭ֚����[���h1�QW����(DO��-�r�Wp�B��X����(����*�y��E�:Х�_�l�:�����a���7p�}m9k��bW^A����8�N���(�j:9�|�姒|�  U��$��Je&��u3�.�%�Ν�t�|{"�}j�j��Y�'�M^�:��I��t݊���eph�]r�q�^I���hP���m_�'�S���'��hp	ݴ!j ��� v�s*����D�<~v��xJ� ������=
�4@�0�Ϛd�`��x�;�K~H[]h3kc&3u�3��s0���ѬQ���}��,n��"�5\�y��6m^�p`4�(A=�[K�۫��jra������f45'Uh��S����=��+�|�,`�Z0[�˿�݇(�s�(,�e�YO3��=gGr=����=����6�Y����� ?	t����D�:g��KMp��:'"�"yd{r�o7����8�u��-�5�/0���-b=*s��ϴZ�P�u��]�����;�B�K�v{>�}K�"V>��_0�������o(Da�������0�����^���������z� (��8�}n�;w��5)
Fk;Г��_�������զ�%<8q��V@�˪�ee���������%�0eU'��@�AT���#L�D��_�FϾya��%���So�;�C9VQJ��. � �8�Կ�����ŷ2�,x]���5 
���N�g���*�;����Z����%��Úc��A�%�P��mT?Gl��6��W�:�?l�1Ԥ��s���[ْ\J������6e�T���������jt�#Ň��J�d���(٦�?˭d�S�v��/����7!�|u���毪@>�W�s�w��W>�u�#����B�J��P�S�&xk0{88�,���PG�L����eCP�%IP6q���*AU�@����o��*���9�A19�?l	_+Tv�6����݀B�"�C�)"�@Я��w�E�yZ5�x(q��=��B1Fy���|���(�;�د�{�̀��k�d���'��a�>Q@|6�a�[S4�]c�\�[�k�o���,�l�!�ᣌcv�ѯFFua�oc�5H\��D��FH�io������͝ ��U���\
��n��Jǚ��Tb~^6�J��NT/N�U��׏H^�|���t�95�
���0�v �7A�ґ�*IX�*��FG]�ʘQ�Jq��7���8&�ȇ�EoŇ��-����5����������
�h/�b-Gz�s��:�z�s��:�Z��^��k��z��n�u��k:�B���Ǹ��6'WplO����)"����3���=����_%��lf߭z-�N��#�U /X(� �BX�0���Ai�,_�d�>�\��},5�w߶K�Éa8'{��lm�l�	IK�M���9�&��?�ք��&(�+ʺ�F���w��_8{�_*��c����D����4��K��~�'���^����J|�5=�'4x�0�rވ��גo����g�g4|	�Zn��FƋz�_��9�g�g̲	3��?d�ܿ>���	^*�ܮ��+~�)s�*|�]���*�	��@�jp�MLO�3'��U �UI �������>0�>����z���0�ʳ?�e�����n}���!g{��8s]���{#u'��ԕ�a]������e<ZA/u�P]��;]�؞5LA/u�T�;��B]��X�* �����+U�Jx.�O������?*�[|💿�C��[1X��V!������a`��522��{�X���8$�f9e�������g�QXn�!��n�H?�ٛa�={������gc��*%zq8��ɠ;�L�O��Xo���i%?1sd����披��kʕ�-�S���yZ�M7i�Ç&xT�2r��b5IsJ����n�z[�'h]�V�f�x���a���X�9ꗪl����V������7�z��ܝ�������zMd>�·kE�n9{�[�t�I�'�f�J���6-+{����V�k-�Z�
O�c���фF�+��$S�{F�Z�Y�6;���j�S��"m�L���Eeoy-�Q��������0�X��-[�?^t�V�W�N����L�}x&�4Z��G��M-GC!��r�}��O�q�#�Y�&�7kV${V�p��ź�XNhF�P��ĊZ�Y���̌�g���w�S|N��sڨTxCC�"]P˱�W̣��Q(<�2w�8w��݅6w��*�����Z$ְ�T�?V��M%Ч��`�
�N23�J��ѣ`��%�e'\�2j�W��͕0~���s+8�[CJZ�p�:�-4���-!��f
����.�sƉ/JN�K8����M�x�Y7���w�H��6�Z�&<zƐ��Y�#�F�{"��)Z�7�a�����E����%�n�,�2GswɈ�`�,��W�T� ���4	��|���!~!��J����?�RNaUōP��.���da&��9�,X=�ߨ9}�#�UE(J
��Ε:���
�@\������.���(���u+��]�|Y��.�?�a��K�rKr��J]�%�U�i�<��*w�*�Vy��`G����u��a�t��O+5_�Uo�~�,S+���=���g�]�Q�:�����XV���{�"����Be{$'�b��ۼf�`9yaD�Y�Z���v��ڈi@�*Q��E�wߢn�k9$�ŮN��|�W8�6![6X����o�۸��gg������3�D��G�����p�����I�v .�����T%jJ�J��������S߇N���N~���a�m��W���7��e�1�6�q��)��Yc���U�g�֬5E,��ۆw�a�m��~��>:�s�ބ�����m_����R;�yg���&��<J��
�諺��e�b�Tl�ZL���+f�bN���b�p�?Uߗ�{o�x�6�*Î�	09�Gv99h?�䶊�҂.�a�V%f��]Za�U���_�6���y���H@1&��;���b�jL�����J���ݪ*�Ql3�;�� 믡�zq�ʖ��6`k�R��oL�ޅ��:���U� uܯ�׬D����hN8;����1y��+��>,~���[�Βx���(�����:M��J �B�w��
U췃��A=q�H�~����ܒ�},.��S@J�җ\{S1�cO�U���"�i�y>7L�fd������:�n�Dw j����y��A1YF5��LRȆ$���֣ ����EM�n1��@��^����p�DH� bNx`��=�%�!�"�Z`���AS#!2�%��$�kN0H�mT<d�u�j�[��e���$�"�@	��*�X�J�.~�� 2� ���f�7S�訕�	�����i�?����n��9�O��n���hϑ������B<�?��HnȮ;�Ȭ���ژ������/���Z4�d�ѡ�q�.�4�N�R���!"]2��}���"����*�����c�Ke�1�n�&B^�2J����hn������hKS����' sK�������=�(������kVd;��ّ�=cN���9�ь�գ9�f?���Ѽ��@�ǘ)L��=$zE5O��N�{L�����@/xNG-ag�JaS��.q�c4Y5A�j8װ�����)����,������\y>��B4Ĉ���v�W�����=�` N���;����\8�9h[���c�gsy�g�I`�`�����%&���`���ߩSE3���:�@����eλ�?+����c���N��a��
�P��+�b�Y�(��R�>����#<f]��M?7��80�W��ˁJ��[%�fe�+�<X�pm�!4�&w��l�߁��χ��n��x*���폢��6SJ�Un��vV��C�J��F]ǃ��2b���`ٱ.�=�2�u�'��I8o~����w�U���OCQ�&�^�!�]k��(s���<�?�ݣ�S><6�ழ�C�I�u.O�o`����}]G��^0����d�[U?���1�)c�Sz�Kd���?����W�O��3xԄ��I,�}d���U����<�f�/U��ғ���*o�K
<�V���]A2�[u�U�}�Q��x�ԝ%(�:Ɯ��-���ҜU�ŹV��(��+���A���ۻ���*�r�=�(��j�_P�{�!4X���j��:`^ᢈ�~W�mj�b��������y����ἐsi�Y^�n���#sw#I�iU�C��n��o0:�1X�R=�5��(/��ʙ0n_����i�!��o��~�IfL�'.�ԡz�����@�i��$~/��6 ��������RFw婳�Ȋ����6i�~�;�1�C���i�QT���6j\��yZt��jt��(Z=T��m�����c��g�h��A��r�ܯ�8��c���=�&�u���d�A5�A����r�[�{=
���/����ny��q�
����ǧ��u����f�gž �R�}�(̓L������B?�Z��o��dw���]a�����M�ju��R���*�'b;���`㚠\���e�V�A[D��נM���j�/*-�Do��/G�J��� ��~y�g�3O.�G�ڑ�G|u�S:-�D��䪕�k��7Ȧ���`����'Wܙi&�[��$Ţ.���"�t�ϊk �q�_���`�4�ə^��D�ޠ(��P@�@���S�$/��(T��?"q�:5��M�PkcovP�����P��S�ٛ^��$$pSUp�����y��|�"���h�C�sC"�H�2��6j�-�eBx�zH~tS�x�Y�����JK�`�y�Y�/��v[r��J���  ��3���Kej��@���5K���o�����iO��c�տ�����8yxح_�8�lb���f<����Պ�/��R��y�E_������`萆&�U+^�1oS�΃짝��aU���U�VVz�Z���L<����s������:�tU4����7F�r貾<��GI�c
�By�i,�ȅUhe��,�G)�G7%�h���c��1!�N�g�Ih�L�>��a����;�����/3C�e�pD/d=�Q�b����!(;aR�z=��~�zy�&蓮Gyc?����ɖH�������}*�R �w�t<��bY���*U��,P��A�wa�֔�(�՜�ָ��=JlI w����	��?��+��<j@ؾ��+�;m���BW�B;|��}��;a;t�+�5���)�m^�a���}٘��ػ( O�E����j�c����)��-w'� �P�wp�v
Ѹ;����	���z��0��$Rd�� ��Z��c{�s�my�~�{H��vF`�I+��Π�Fm���@C�`F.I'	�5��v��/`�Py���"9l���[<'쏵�ˠ��ρ��X��i���K�.]ܭ3n�\(�u�Gx��s�t��P����ݣ��C���{�`�m��z<)�hocn|SN�EB�&�v�j�(n�m~2K͏gw0���,uG�Q���.\���.��K�#&�25�mR�.Q@W.U�Z�i��ȑf��r�M-����6�Z�VA:jy�|��TbZ3�������l�KP�E�wp�(LX�@���k�ܔr�!D��7O���6�a׷�OM��O=J[�sɹ����Q��h�q޿@�&R�M����>
��c�CK������>ʎ���R��p-�@rK����7���Y�^H~+m|��#!-�m��/��q�ͯ��m���K9�6�M��_4�6��Na�EX`�0�^yH�^.T� T/�	�uBuD�����"].5�j�EjX�ϓ[���$(�>������l�4�����Oݟג���OA��Q2�s��A3�2�y8���y穇�os]Dmi���HeU(tl"��Z�7�����v�%e.U��=p��_��(��KD�p	J���G�j�F��#_S��ݚ�w�l�X~Q�|VYAM�6d��7��|�إ���>���Aj8��%�cB�O��Z����D�p������F���;.��w�^����)W�F�h��Z{��a?�
e�����@"�ͳP{L�#�N����3�.De!�!D����'��i#~���	ېL8@dB}V�6b��L���	�~���m'2��3#�0^#.��I2a�:�߂����L�E2�4z\�vE���s������B�1 ��7:`1X�F���d�@\+w�Vc�Csk����^@�5�
�V��[	���ѹyR�����/eTYb?Z���J|PUe�M��L�ߡ	oW�A���3	o��%jK��izI����¾���#~J��\���z�z���V�>Da���S��Q�� %O�v�Zl��|�OX�-U���!8W�pn��NV߉��7)�l֨=^ۂb�����-+�cx���\J��������ˇ������rE�p5��A-J���\�Z��I�0K��q;��@#w�9m��j�q�/o��qM|>�uԈ��f�Jʪ�ʪ�?C�n���<��pi�Gk�G�0�?�w���ё�#a��_����# �b���;e�yP1��l�s�wǟ�'��Ӊ.�<!�]��EU�.�*dHV�4��Z�{�}L�{O����fH6)>Kz�IZ�K�~�Vm��O7��r��h���?B
BM�e
g1�#����e�Y;;���$���f�i�����oo���:$q~W�-�<>��xM��c�jh}R�j��VD�'�)��ҵ��9����$��7Q��,/�7aA�I��D�p.|���t��ߧ��Fo;�ѽ�ݤ�3$I!8Q�F�&J��u"��F��_��t�6�A��$əBq�c�yF����IXf����~���Ev�"_s*������Ӄ����BT�)���a�k㉇�2	�q��=i��d��r�Cfſ ��m�7��T�x���D�9�(�Ԇqy��:�7�i�+2���.1݁?"�Z�9�[n����w�`0�U���^x��"��"���:�L���Ӊ*�~�A�_/��_��ӪD"�=�s����\�m�q�p� �^l��F�6��jU�4��Y����0�B���e
��|�����J��k$�{�v�c~�GI�Dm#r�V��r����Ȝs��uI?��=�Q]��Z�:z���Ԁj6?���.WƎ��ǎީd�*nHؔ:+\�ۺ�Ԥ�XtGa��DOz�W届��?e��4�~\��]���?;:+��=�<�Cg�YS}�t��X*��/��Ә�?�L'���Qhϝ'o݆X?O��DĴ�N5���_�O�+�.=BD��;������T��l��^z^S��a�����굆VRC%�Аx15d�7K&C$S�1Ͳ���z�5Ͳ����]U�8&β����̺��Zۘ���Q����LP�8�}��8�G�,�O�10��tD��?�����D?s{�g������G��`+�K�벬���W������!DGeB���t8�w(�[�� ��}ӄ��L^S��2��9���X�ԬN:���q�4�(A��<�� ��}XpRBhq��$�o�-T:��\D���y�vt�����ϫ�_�;hX��ąUx"�S�X���M����!��.���p���l�!�("��;� K�Ўln�`�gd��/.�!�;�?zkr8;�K��R!ڷ��~��<�����Q~vi�~Ǉ�]�����;�6���;�tv�mq�߿��5Bm�uok���mw��}�u^�������h��;���׹(�?��Uo�q�yzHkm#������S��[(�eFw�s���}R�慳T�`���ބ��.�N��k3ЋP/����=�
;LQGP�EK�2Q���u~�1UԚ�f��LM�(vi	��O�RJ�7���M��
[�l��1��r(�Z��P�����������OMl�,���O��gJ�m����=����<Y;1V�2�jL��B��q�S�9�>4�cp��^�y
�eIs]���X�,]�5B��`A�Km/��/��/���B�� �?�C�&��h�������MVY��6� �,X�JŪ([�7���hK����Ҧ��Yڢ�ŴJ|���2�����2***BA�����(�3.�F2P�6�9�]�tq���?�����M�w���{�?�~f$��.��� �}� ~� 2�0�U4["������0�@�|�:��v����.S��Z�?�3|)���@�>�b̑6��%[�W�!'�*~o�)���C��gz.���!n3Z/��vṲ��k�ƪ��|���<GJ�g�'��c�u]s\?_����� O�o~��7v&GJ4�h������DVd�D����#�xd9��t�M��zw��4�"k��%�%Q�lW�׆���V��Xϊ���xQ\���ǋX/��1m�po?���_�>�D4�R��1�ja��Y�w]F7�]@�M��q��((Ǎ�.�6���%��?#:&�\�2i=�V������շ�zR����s.j�%��<�m��ځv����sy�J��S�J=��$�쌅��?�{+��ㄌ�P�k:�Bؿ���K�r������-�W(���ɀ酪q�	f��>�����Ӷ4��Ӌ�'b�v|�6r�3n�\&4�(Ԥ,�AF�|���Co؜L��*��@�y�7�9�7�OA��J��XLbY�?<e��<�K�t� }A��k�G�q/��$o{T�T ���#����4K	��i����/܋���iV�����-��8	��Nq~�'ċ%E��yh��-�t=[$��.�|�L�i�bcXHx;	�Ն����'؇Ky�������꠳+���@���'O��#Em��q|�Oºqgb|mĪ����X��q��u��a��bH�~:X���\�]G��߁����/�^";�6 S�F��o����e�G�H{r�Y�! ������W��G��
[�C��.bp��&\<�_#���o���!�K)z���@7܍��������6��b�y���Z~��8N�����&��`��^���n�,?H�UA<Ce͚u��;(}h��όԤq���̜@ȵz�-N���N����2�1� s"�oBa���G���f*RH'f�����9��|@P�!)),A��&FB1�'l��F]��o{��2�n��0�p3�t��m��д�-]��:b��G��������k�YOԋ�xW�#;(2��%�/��|H� v�`��nM�@��=�m�]A�%��9`x�
[�/"4S Ȼ��@c!���]��aI_�>�آ�#���P�~^>`��b����G�O��3�nv���Y4b<����A����xq�-�Ċ�I+L*�x��$궜n<����1�&w�z��p�p�;x�`xS �*>lgU�9q�_�و��m���n����Ěcb6̓���{��q���~��x_$\�yo�s�]62P��資��+��A7�m<��Bse�rl�؍J�����a�,	L3l�8F�W,A<�
l��>h�2]���K�I�ob#]������GF�D���d衷z���G�H���q�7�3�Ehyp��@�_<��r�}�z�~���k�4T��!����G�<�~�g�_��Q�p�^��u��������q��}�>�k��S����!��_��"��M��{���}B���x���7̢*��_��=�J�1�$�AU�1��?ZO6�vn��\GĝQUQEv��lG�6ه�|��#p��v��t�ib��yE���IQ��c�N>E��
����e��F�Af!��1d�����z��nF��#x�4�{�zaiy�Di�wL���=�w�y
5 �$���؁�Tk (\w~b&DJ�ɰqle���< e��X�b4��]ӎ�]�����HO)6�Gk{�b���1�"��&�X���8.�ʺAk��f.k�(jź�,�C�I��g��X��@%�g���H��D��Yg	; 5���,U�}��
|L�xQH�������}�^3��iG�x�/���5S�ė!���A�;8��{�b�T��Y��Ԏ��Q��L�hx���HH'x�٦�0����.�w�f��r����Ia�B!�=ׇ�G#��1:B9�|������szRs11"-~��@��&ȯ�2Wy��K�m�rX0�ť�%��`A���蔲�@�'���UpQ�F~B��
�����K��H�l~�<� �u>�S÷��,!��oe�Z����E\��Ö��w�S�؀r�Z3�P��XR�bA�.4�+��,O��?����5��i@���(&���I�;f��{�*��D�U��z�@�#@���(� 
���g	ܫ��،<�{�I�`�Dr���a��V��Q����M6�����0l<�K�F0p�`�"�=0�I�y%�=H��Ey/�H謁Ĭ��,���=�H>��yEU��;�Shk��c1�~�{
3#��K!kq���+��:�U�]|�uriys"ȅ�8��
q��H�:x�H��o˳�/|�,��ITU�G�w��]*q��g�f��M��G�oLc��a�����IM
L�[_FG��9A���ki���Vņ�c���Y})q��ɾԉ�=O��������9q�O<#�{�<����/����,�1K��ً�-Ր��K��-�]/���⠭����/5��y��/n=���¶�o23s��G171|�˒������%R*B+
��8��wK�y�#����K�̐0�u�~����W/L�Pv�c�Q>3�I���s��9"�[Wv�n� w��z�Yt���x��G�[t��z��JV�Ën�=�^t;G��<
�}a�A.}}-\��Z��u�5�֑G�����x��Z@��^�~��<���ژ\ ����9�������$=��",��xU6 ��6K�ci���� ,��ɔ/sb_��<;
v7Jʵ���<ԮU�0F��ޟ	�t'�kX��p?��܌�]�'���c�g��$'���y\m/j=�2�9�֓�-�W�ۙ�^|�E&����1Y��,�mYY�a^�8��(�6�b�t1j1
P�.���hh����꿁�ɹ�, �q��PVt������?��w�?�{Yb���VA%��A	�[�{��ؑfyF�Y�D�"e4���_�B��a�z��Q�$�f�� ��̏�O۷ogH)	�@�+[�D���Qp�W(�� �߲Z���z��D��������(GT�#>~E��,T�7��yL8����;$P�\�X8�b�IH%�O4��T�2�ϒF�R�����'_D�0H��B����ש]<ڽ��y�`�O1w'D�H��xr�� �X�����l�#��c20�3�/n]0C����P��y1 5M�<">�+���>�l��AyI���j6ø5�K��`2d��RU���ǫ�t���{t��Z��߹ ��G@?}�lO�KL46sk����!X{ �f��܃��}�z0�j�5���+ �yЈ�y�)}F`�n���4��lϝ�Hn2 6�Q��(�<CYU�g8>��M_�ZD�X�@�EP�_p5��	��\)&7]���g]����D����Z�G�M�t4��;���Ѷ:�����n'��Fo{�^`o��b��=���{,}�����W�0��ec�g$�2|�M��ɾ�it{G�vCoa7t|��N�n?��ӛ�ao���`\�i��1���_V�����@f�kW�אY�Ƅ�?�0$�������0ϊڳ�?�F&7�,��RE��23T��1!ؐ/�)95�Se�Q�i	��܈�f�(�	�S��=�w:ܱL�+#*>;�?{.��|��}��D��<&�tҚ� d4<*5玌�q��c�OA2�?� �{����muZ���`*�-r���[��7t��P�	�9��"wV�I�d����BI��C�P�k�ě� L:��tށ��/��Qy�P�q�����L����)��oP��ȭ?��`0����pl+����#�üW����{e�d�pb1��sr�]��� �c*p�:��5($��mPY�^t���$���ޜ'(���|��F#�-N&t��Z�.��h�ha���YR�V�~���-�P�.��c4�Y����tt��: \I�;|��xk�砾��9�%$�p�m��N�DF��3�'�������j�H�S�k��/&I�g�����@A:5��6��O��$��	����8����Ӂ�����BS$�.��
2��ˁO7������!eWA)�i�uL&u�n����F��|ԭ박9 U�I[��l��V�p����R��M��a�b[b�� �?�����.��x zq2,�ʫ���/ �T�O<� �4���nj����������=��l��Ɂ��(��3���;I�nt��z�vow�=A���.�m_uL����&�j1���u�ݺӸ��x�w�z�72q��x���(�_�+���K�m<"�#e�em����p�/Gr�Q�Q�{I��ޫѱ�x���A|�2ѳ�[�(\]ދ�����'AQfV�/��|Y��ܫ��(���.�qӏ�o�0Mc�4����9�>�f�=��b �bV�"�n��V�;z%cq�]�HTlK=|�Wѝ��Ť+`&�.��xq��J���<�^EUv��f�q�'BJ�b������R��q_�3N��������_�����YFp�O�'����oB����xȀ��F�6�c�Fe�X/���-L�'�ȑ�G���y�Jhp��4�WU��B�"	sؿ�rD4�B�����tW���"��{��,��^���!��N�����k��jqfXa)��Wt;����$�yϟ��ݏw_���2�pF����x�+[C�Dƫv��G�Z���rݘsD1�0�*�	��]I��g�)�
'}�YV0̢�-B����*#�y7�}Dm��eMcwMU��յ��y"yJP�%��
7����
w)� ��F���qvh[J��ú\F����&T�H��~��� ��/^<��q������ �\��w-~�?P���-m���e%��&01v�o�.�����X�T�qB����@BYa��`���DV����m�:�^|��|*��� R/{�kM����V��;�V������X��(!,F��w��n�x���^�/��_�m��y�����{� Dt�m1E��KY���p9��	|m�&r�t�wI��!�n��E�u?�?^E���ě!|u/�\,\���]�c�r��G��� �\�P?��-W��⁯���w��
·�{;E��*��7��h7��-��L�S _�\XF6�R��`}���g�N�z���I��M<# �)0
���6�S����OXn�VW1����r^�h �_#'����9ݒr�W��5�
6�!L��$�n�욐����!+ؐ�態3-,��*��$Q��KIƍ����
��1���L��>�	�""7���[m�֫n �|!��OjP�G����]ӂj�l���AJ�X�}�?����X�A|�*AR%�8��fr�O�u+̀>#�y�/äo��G��$Ͽ9����[F(R&#�E�l/�N��N3��e�j-#���9l=)�&��@2�����,/�u���CԮDr���b�R�s��l0�y��ǉf��2���r.������d�'���S��/��F(y#g!�Dbȑ[����J4肨	䅦;�ao-��_�E��`�\���R��BgFq�i"��E,)�G�7��
��x�u����+r���ST5����./�������{>�{�@@by���sכy�'��S��6���s���&Q������I�L���^>,U@�X�������]�M�G���"��{���l�!7 ����/O��]/e���0�BTz� 5�k3p�*`NO������I�3���ʛ[,
6d3�}6�5�UQ~�����4�XD֒m���L��[�d�|��1|�I�\�/7ٗ���N��1v[�Qc���G�i�C^�pt�4:� �����ǟ��V�Q>�(CǇ�����@h�K�Ť���w��ܲq�r�r��BAUVn�/0���6�<I���V���*�FE��T� ��31U����y���9K�(w�wu厨��^YMj#�/zwcr���Ne�^Psy�]��f'd���	΀�e��9�u?!и4A�ζ\~г˿���wA���/�Y�U!n�y�,��m������ �������87�P6��5c����c�f&g��{cO�br�D����$_�ɗ���Lõ�=}kc�sS�%a+���x��r��G���/}�/g�Z90`�Z�%ޢ`v3l�\3PO|�%��8ς������6�����Zh��!3����܂s7��
��R�׸������S?��-J���7.�FMۜ�E6;J}#�yH%uEiB-�@*���b�7�I����<;�y�P�`��� ''��YT�!���g�ܫ`eL�6"���ěQ>	�	4��_���u�+�o�� #s��&�����{�{>�39q���G�psw���n�Α���lN��{�o�o�ؗ�8 .2�,1����� ��}��]��|�˛-m�"�j��ת��"i1�����u_�D��8���5S�ڗ)���U`�`;�.� (���W�6i���H������,��h�7U�rl*�N�)�-��'�O�-���|M8����=�������eK���BT>mk$��������x�ITQ��	\���H{�����?�P����*��k%HŸ�E�^2d�#�g��C�d4(�irV>���ף4<u=(�{��s��^𐅔�\ �A���L�8;�~ſ9/�,�|�¯b����3�n��S�6����C@)[��{�5���;d&ț9M����ӆ�`��DV�?CmT!W�01x<�-�d1�%v�#c��3��8�4.V��X�o��Ϡ��csNvD�-�q@�H��3϶©j��HO+UR��ϰ����.a�x�Z`Я)`}�=�e�%��17�L�)w�/CR�kT�= ��q<ѐH�X;JY���wz�/#�HY(����Vۈ�$ɷz�o�d�1��e�H���Yy�Y��r��pt8�W�ꑎ���%M���?�5��x����_SF&�o\I�����P�G�����D�@�������*O�:�`�(���5�����@���`�%I�g�G��c~�X����b%���d򊪑�0��}K~UQ%�į(��{^Q5��+�>��+����,�N3y�U	�G�]u~����T�e�ll�v���]��(�?	�������FA��J4�~aV��+����CDFB(z�ƚ�y������-Bq��h��Q�'�_/q)1�^1W(1&p?}��a�-��}Tzޝ�K�Zk»�I�I��t)*G|)q�<!�8g�{�%	@��q�[�M�V��ɓ���<(�BKy2�%A�#�8%�j�-^hd�fǪ��F6`$����CB��-�)�_�}�pz+C��իa� ��J\�������{9#/7*=	���ז3�Q�Fg�gdtG����s��v�� *�Cᷰ�́���V{˽�.�q��B�<�e9b�ލ��}[Ql�FK�rfT�Q��|���A%6���xQ�;6�ʺޯ��C�yٌ>��M4^|k����,Ş_��Mn���oMJ�I�:l2�ў;]m�v�$��I=�G��|�:�\�zz�D�E=��	�A�⼧�D���u�����wn��ek����5bʭڳ
Z1ƻc��b�&���bg+�?�I(Auۡ1��=��2R,���	�H!�\���ۼk�HMhXٗI$��I>�
(o=��؃��~�X��(��=װ���b���F�]\t���T��c�%t{U��ܗ��-�-��J%P�Y�^�N�D�g E#�)�ϭ%�"��D��ȣ��6~����nW�	����g�ˠ��S�5�^�fb����'�\j�KU�����l':f��n��;��}�mE���]���yG�t�r[���s%����'P���1��(�������|/�UF|vӷŶ͌��Jk����n��<+���]L�n�D�Ķ��$-n<;����α|��,}�7}W�7}GR��D��5�ּ0��C2ta��w���ۓ|�Ҝ�NCLG�<&����U�v�)�x�a(e�w���J2�ͳ��������0��~�J�ž}�mi�%��e�g� (�4&�� h�À؃�o���rV��58�e(�G������9�b='�uK�sBX�R�8�a[���MA�I\ۊ(�u))�'=�'����նUâ��2^p�	\9�K�E{��].}��+���>9���3�S�`�f�C� lӜ.�m�?��	�7����s��U?�y�W�;qC1��+$�66�c��z�ѱ��q A{��'IAn��K I^��]{E�\wc��|gH�;���s#�����4*F��9G��`��� �C�}�����u�`|P��Z�7;z�4Ǝ̆��\��'9zɭ٣�>���^ N}�'2�%m�e�Ў��H?�~����l=Y٪���f��N��7l}��kmĥE�[���;���H�艔����I�VkF��/.�;�y��g|��`���VV ȟ$5VRD�딀���]uĶ�A`�I86OOv�5���F�2��LF<3� f6��!���KȘi�o�7PҙiP!X�ĳMO��F���M
�˟5]}g�@`��G�w��P���̟?���~�����mi/jG���MW�� �A�7殀��}?^��d�}]�v�d�1r�Ji�� ����l@����M���&�:�*��:��f2��-E��
�����!W9�*�?�'Δ8��W7����W�:k�U^�f�%���
3����W��+Կ�O��;��_?a���w����*�pgJ����6��icJ���ص��w����f�/��G���&0�����G��nnz愡�
�i��]�g������qN�#PY�v��z��c���Ey�/Sq��M�Z�9䵂{P��Ϛ��s�J�DUĬ�� ��Aȶ����#�?�/4[7��Z���3��xy�����J�,�9��I8�R@A	���Q*Hv��	jU��{�N��и�9 �\[V�17�q#�O���ʝ���I?�ۘ��T �b�Nl����/xB�����;���K�	�cse9��B\�`F���	Àb[&ɝ��u�R��G���|��Ж%2������pȾ x��g/O�xc���;OD��!ϣeT�~\~^�_�l�t	�`�"�d n��,���-(`�2{��ތ1��<v�,�^�6T��fSQLF��s�(7a�_F"4�7H��S~��t��]�(v=L3;k"]lE��� ����i���3s$v��^���r�YX��|v13G����.�e�|q~��7�O�˖iw�î�'P1ۚ�C�_���eG+ߎ�=���n(�sj�� �f�y9*]0��BC��O^[��b�b!	Ј���E�R��>�e���ܭż����ۜ@���uy�i#d�J�o��jh���DT�ǳr��"J8U���˰�O�Z�ѿGBC���k��D���'��SEq�Ld%�v_4lsΝQ�_Z^{d1����1Fã����I���B|9o@%�o�$H�fI��,�V�e����uPqPԗ�y'�Ɉ��(o�$�͕�q���A[��1,fBk7���N4������:�-�6��ub98Ο>9��m7>O?�+(b��G����Dw5��W/�n5��v}�4��!�8�ؖ���#1^�m��Al�!Cǆ"����S4	������0:��ѬM�dd[K�W�ę�����3׵e��z�%��;�+�E��zR�N����詗�t>�F#�+�\�;�î�r�D��G�{�� E3m�@������BSR5�,��:�z m���ǟ�-�`��%ZDWy�ӷ��f	�$+�0|�"� �}���0_0���E�9ݾ9=ƣ�/U.�L��m0<ջĞ�t��r?���On:6w��"�4�]E�A�y{�x�.�G챭B���aR��o�7�띏w����c�o@�I]v������$�l���!%?���ws��f&5�!a�����7�WC�'���/D�~Lz�(U�C�p�*�u[���Ұ�X&�˗*����0m����@����*\=�oܣZ
#��L�x��,x�Y��Y���_,�7�;���h:�z$��4*Oƶ� U�`l+��C�hU��(��R!�2'~S�L�(h����
��� ��W�f�C�g�/C¤�w�8�ަ����k?QK���c3��yxm��[���ç�ўa�[�=�u)�������o�̗�hX�M���q���90�.���o��\�m�\.i�qYس�ɞ�  ��3QZ����w���-�a\��P�O�8�0D��7��L�&��dL�.�%��6X�@Le{6�*�$��C��i��&^��Z��������� ��D|�ـ.U��ބ�����	4��V�sZ/���]���B�6����ҷ�Xa�Ʊ���R>�ȫ<�4tq�an���A\�>�t�~n.
q/7"%Ɉ�^����Z)b[�y\��Cj�2?��l�&T����^dQE�F��}IX�m��f���m�9��~0Vt�2�ygx��8x��y�����*�]�
(.��������Z�5�ad=����`(�f�O%+t90E)���E��<������b �r�0��'݋�)�
E��в���7�|d��� VqL��,_��=��&KCуS�t3�#/H�G�����9�b2��Ra�'��y�hK�n�/�s;��$��hwum&!�|$��.;�Mɻ{��c��0�����e{ΛU2��;�˃a��RI!��|:x{RM!g��0�M��8�SiT�N�&1��,k���Ux��!�"v���SW�Qv��I��%-�W�]��
k7�����?*�^5��!ˆ�.G� բ�)��,�نhNT)`]�2�����]��տ�
�=��ב>K�*��]{S�@�H
��H���B��x��!����}��6i��s��s�/�w�p�x/f�����A3H.^a2)��؍�WD��Sh9�s6;���#F����D�}Cy��Fb���D& �x��7�لwd�!����|)b�8�ð�=Hd�F���xA��sm�_����h�ήY�|�f?������0�x�Ύ�?�����e�V�m	^���\�k�9���0C�|��\����.��?��H!JS�t�
��0J������m��vow۬8�X��%�5Ɵ0xm�N�w1�a8:�($���_�L��
]�T�D�/����K���#�E�k�$!Vi�_�_�(�n�D��R��ټ��u�x�%q~�� U!z)D�4`�����;a�7
K΋��=p7���`b���[��ă��7�Pb���_��6�R�=��O���h�
�/#������x�����Qa�B|�{�a�`�TaPԟ��%N�n�t�5�P-�Į?ǃ��I��h�Lzş5�s9Q�����h>{���j'Gm����<S��1�k�xE�U��ǂ
�Z~�����5Pޟ��_��/zAE� ����s�m�3�p����G�!d�jր��������v``|�|C�$J�J%C��͂�~������ӿ*YE��0�֭л�r.�ɷ���I}������1�}�t'�C}pRX��>tI�"��Y��Nǘ�/X#��5��x��Y��%uBUb�Q��=j�����&B����x�;���Y_����=l���B����.�}{���q|'ݲ�d��ZT\���Y.Q�;������2�ρb�a�EL��^�햺�{C].�r	z�&ˣ�� Qvb ΂��K���>O�7��Uj?Y]���*�,����wGt0]�b<�l��������s!� ԙ%,��*Y�es��d��k`�r�r��r�$�/��&.N��Jқ�>�\�n��݂�~Y ��@�|���8]�4�ؕ��'ت�m��?�j�v���i��(q:�]���\�"Pi�FX�ᦵdL��3Cش3gpZe��0zX`�����FNO^Ȟ�r)�?�Oρo�8�="w��@�@�A&{���`��s[8��&��{�-��O���@�s�F�����:v�S�S�%���/
�VrJ����r�i�@·<�":�3z{��7���*q��:	���L�o�����r�Ub�@�����]��F�.Y����sQmY_N��p�=��^������s�.���c��<�R޲�X����k��n�,R�~-z&捔=Kxw.��=��$-�m���}�Q�gXg��1sàc0 ���}�N��Hy�����{>�~-�	���U��uKg��[O�1++�/�D*PM�]�۟E���d�����O6���B�����u������ϱ����������%���_�σ������%�~6��ca���>�O��Wo�D�m��?�<%:����}@$z�Ѡ��T$��i��a�FD�ZFDZ�rb�H|s�h��(*��[[EQ2�:����(j	<+,=�ZEEQ��г=�Q�����oBU��]
{V�* �8��>x����������Fس��C��lسnxf��;�ꫪ�����ma��g��lo���_E�ѽ� ��Aٯ!]v�K5R"$%�\HK �C���"������(��ZH� m��
��!}	������	�ғ��CrB�i&$%�q�� }m��tR�5A�߫����r!Yp�!]���%� �[��H�`�~��z!��t�HO@��^HM��Bʆd�4R�k Q�����!��H[ �i5�rH�����C�ca~&CRAʇT�H�B���g�� ��\<$��5�<}pp���>�Zi,����Cj�4�x9��3��a~n�/�||I�!� eA*���$���~��$����m �A�	s���E�ŵX��J�CH�!�
>3 ͅTi-$9�O�T�	i}ۏϠ~H������\���S!���=�{�X��xv��z��p�c�.h�[H_B:i/���!M����)�|H`1Po/���>Ի��(�S��
�[xwR-�Ր6@zҡJ�n�/���N��,��S���ln�}�Z�(]^X��Q��Y�p�**�)�G4��Q[X�t����T�(��pT�Q����
n{I�Ǒ�TDQr|�Z]�r�r�����t�O̐H�TWו�ڲ���ʒ�ʻHeT�NsT;�Rae�'�\�P{	���p����Sl3h�Բ�j��**Ta����T8Jݕu�T>E:�UR[V�(�4���Nw:��$�v2��v�(>��r����fԖ�9kJH�!�J�8��Z7;�1�v�o{��lGIC����Tz��������AzT=�ms֕:\�0��	�f@{�� 䠮��J*�u΂��eՎ�K��^j)Y��ʥ��J*ǌER�ʜP�����u%e�{hsVz~nz6?���`�E��eu��u����0�r�	�O��D����t��K\.��v�9���d�'3h�lu.w��ҝ�*Y�4�	�j8U�ꬱ�8Kj`���lU�����'�V��Y�ݙS��Ϗg4e�*���R��H��~��{.<��ǣ�\���P�]N�]�X�,����Q�r�)�A��x��]SRY[�\��Dť��Jx�TTL�TQ�sK�����K꒨��U�ti5���b6�?��Қ��Z�Sx Yk(����Ƶ���:-A������(}������ԕ9PK@~���N�%�K���+���<�S���]\A�ީb��R5��R���-e��aDnG2������0��Z������\t��6�r�ڀBu���ӣ���@T1�dU��
�-s�ֹ+�W����̓�L
֩�MvS���\���(K��.��5unG	L U4#��0��**,�S˃���	���Q�`�_��ð��*��,�-uT���ֲ;S	�C����x�c�'o�A�� ���j%E�+ʯ/e�̩ur=�Q��D��7�x��]]]Nm�'3j���pR�+agST)>�`p<�vE��]������?뮥���䇷�aXO\شn�cEz=ԑoK�/T�#��ō6�| Zj5E0��V�.)�6Q�t�GP��6{v�Դ|;P�BgI��߼�[g`>�GYzS)�qA��QOu��M���/q:�L��m���S���Bm�S˂0V +��k1N]�����)��l'/X��:�C����t9y �@?��8��� ���G��r�7�]\�o�RT{�L}"��T`]����c!��~����NG��@��4��|.�!u�8��~]��A���]Y�S��K�,pԔ�W�9���4��zHQ�q�x:7��<�~X\X���?Ձ�xjM�4V�K+
��:Z�C�E9C��M�G��N_	��U�9 �8�QC���u�{j#�;\�"�}l���{�����p��F: (��}Gc�N�{F��φ]S��QSMS�)�M�~��{	a����L��t�ܖ�axI��J�t՗���hes8��~���Z6��AzB�q��<���z%K����!��z^V�;�j����{���=N�a5�"�+a�T�Aˣ_�sX��sY��:�ɶ�(u�7X���� ��!�]�S[)�o����9����!j�8�]*P�`.:nxO���#���#��g����=8j��g.0�c�(����w���]����g���7pK�k�֓��N��m�J'OrM܃��2��r۝z��5�%�ԫ�o��q��ɻ�ܯ�j$�%���Q�i<!ˍ����!'ԣ~i]���^�hD<tˇ�y:�b��~V�<#��​���!E���S#<� 3��ND���mQ�
la}��
��7��H�(�S*��޽2�c#F��:
}�S_JCIe5a'�GD���je�!p�`���N*��j��������*Bϝ�B��Ҝ%��s+�"p���A����<| �~3PTbr�j��h�7��8�%l��8B���J�Ƴ+!d�e�.Y*���5ܓ"�Q��>�i�V́�\_��E���������m3�z�BT|��S�n�����%��\Og��re����R�p\%��,�W5�������ɿ�1�(���_�~��C&���sklx�s��bJtz1%�i.$	�=�(Q�xH�R���L����-�D� � � ��O��BZ)҉y��DH� �/���VA]�� Q��wS����ArC�I)��.��.H�!-�$Y��{k=��Bu����_*f��?퟈����v"$T�&�g<|΅Ͼ9q�y�~��[x>LLQ{�	>?<����M�FT���FQ�C��vEQ/G�~GS9��z&kSMu"��(L�'(��'$:j�� &�<aNa�݄D�����V:\����M7O���ZW��Y��8��Ĝ�Rg����ϝ�u,MI�2s�v�,�^��պ�<�Z�$`�]Sj�rS@�7��j�6(&$��SY<�=�o�U�(zT�^9rx"����
!+����_�)@
��-u_h�Ф�pj��']�ʲ���XT��f%T15?͆H�+�����ZZ	O�a���Rg%��,�9Ivb>P'+a'���W�4M�	�N����~���8�	��Q�~%��<s:Vx`�e �6 I\�p���̒�`7�A���̅���yB�kFmC�r�sB�,�ʔR�a��j��O�i�=�6x�L�b�&���/8�9�����*
�����S��m5�ʅ�3�o|���e�[U�������G��"�o��D妜T%UK-��*�j�5�R��S��b9H r��s:���lj,<O�<5�J �J�M	�r��s��R���rA*�6In'�ƿ%���J�DB�i�\�l%��`�i���SM�%B+��ra���I�V��jա��R
HZ�&'��]UP�D��̄��ób(�1a.̍������2rh��)	��s�&�����f��7�kD�S!6�[Fr����ሗQPE������T��CM����E~�lb��o�D�.��gs9+���sV;H��³&򼊺��H��(�����%�Ii��4�s|2ju�@�Kh\	oqkH]ө�~m�]�_[S��F(��q ��D,���B���I��%������-���=��F��O���G[4g~~����.�v���[w��\x����3~oC�^ϒP�N�߻���?��R�;K�B��^��<�{��9��m\���E�s����	z+���A�������W%�UI����*��P=W�P��z������������k�_{^ۥ�����hu:�.Y����e�l�B�\�T/�����&}�>M�����������%�2}��Z_�w��[�O藘���js��mn2�2�5��כ7�7�7����0o5o3�0�4�2�6�1WX�-���ɲʲ��bYo�d�l�by²ղͲòӲ˲۲ǲ��n9d9l9f9a9e9m9k9g��ⷜ�tY��6k�u�u�u���z�z�z�z�z�z�z�z����o=o�^�v[{�&RT.�\,��'��r�\'7ɓ�i�,y��^�7�W���[�����{�{���C���c��S���Êc��S�ӊ��s�je�ҭlR�R�U�(�+7(7)7+�()�X-QK�2u�:^��NT'�'�'��j�Z�6���i�,u��_�%�2u��Z]�v�w�v�v������M�L�M�L'L�L�MgM�L_����.�%S���D���i�,s��f.4�5/4�]�Ug5Y��i�,+?W�K�e�
k����6YWY�Z[�H��܈��T)S�)�	�D�\�R�&e�2M���Vڔ�TkU-����M�ͪ-�'T[Uq�xM�&Q�������kT�ƤI֤i�4���P3W�P�DS���Tk�5nM�f�f��E�^�A�I�Y�E�f�f�f�f�f�f�f�f��]sHsXsLsBsJsZsVsN��M�&i'j'k�Z�V'��*�Z]�n�n�n�n�n��	�V�6��N�.�n��^]����������k�_w^ץ������(�X/�'�����r�J���,��үշ���7�7�7�ߪߦߡߩߥ߭��d�8S�)��hJ2M4M6�M*A�_����$��0��P:�N���d�8]�.A��K�M�M��u*]�]�P�DW�����}��� ��0`?���s�H'��ɴ�V�:�D�8nR�R�U��׫7�7�7�� �٪ަ��g�z�z�z��]}H}X}L}B}J}Z}V}N��گ>��R_Rw�{Ԕ�_��:#պz�[\BQ��I�Y�E��|�|�|�|�|�|� ������k�_~^�%�$�� +$
�B��S�+��$�D�d�\�R�&E�"M���V��*�����������'�����g���K,eĂk�t�h�7�_o�BQ��W�M�U����z��&�f�����m����]��ʳ�sʯ�~�ye������-�'�[����v�!�a�1�	�)�i�Y�9��f������-��"��Y�-	�DK�e�e�EnQYd�8k�5��h%��>p�'*̊��R\Tt+z㕷*��qf*K�/)�dj�:E=_ݨ~E}P�������k&i�5�i~�yCs\ӣ�����>�ݠ{G�w�M�iz�~&Ч/���[ߣi�lP���ن��j����{C������s�_��2^1���7}d�`�j�5;`���O�W�7Y�-,��w[���i�����go���m�j�J���
��@qX�oE��J�R���U�[ʿ(�}��~�~�>JLw�Wh�J�����<�����>8�����i��~�����X�(W?��2z��4n1Z�����3?m��s=�2�r��˝�%�R����/Z^��e�o����+�������^k��:պ���Z���~d���7�����ĸ�$�'����|��3�`�#O���_�ኅ�E��E���K�.����ƛ ��Lg�vz}7��d'}�^����]�����U����eL ����T������ru������}�1� ��x�X��0?g��V����kFin�ܩ�h>��E3N����-׶i�>�ݡ=\�7ڋZ��H׬���C���Z��Ka�Q���K��>�0�p�a�a�a�အ�p��O�O��|�v���q����i��j���]�ß��Ib��'�uf�y&`X��Q��?8��,��h�Œmɳ,��`_�Z~�X�C�O,��lo��������	����,��D��!�qr�< �A~7� _ʿ�t�H�Tha�;�
��7�(�
�&V^��I9Y�TZ�����B�be�r���v�A�I�ʠ�Z:��@O��aU�����.X�������t;}�>CK��/\ƨ
T��ǁ��I�O�y�U՛�}���� VN��hi�v� ��=�뽚�@�E���ah�h�Ӿ�m������	����i�˺ׁ���=P[�~,��9��@Q��o���?�_��F�7�dȀ�Yh(1�bx��n��p�p�m�7*�c��n�73>	+������ogtv��5�AS����ss��G�O湖E�M�#��3�K����"�Rk��*�;��K���� �LqFq��'�P��0�z�te&�h9��^I���*�*C�x�wTU�nR���4/h��o�����G�/�gre�JC���C����7|j�����ܨ5Ά��7�4�k<j��@��t�����)�<�|�Yc6�g�盋�u�V�?�~~���EbE8�b={����?�x`0����D�b��\Q��n�O�(>��+�w��J5pt��]�(T�N�M���e@yQyUI�C��t=आvӷ���T*�j�*G�K��{�z��v�]�5@׿W��ib4� MQk��0��i�5�hFhe�#�k��۴/j��Ҟ�^\����X���	�L����b}�ީ_�����bn�fP�2s��`��f����:c��N�4��8���~�G�O�g�w�f�֛ ����Vv��+up��m����є���^zD�{��b C�T�]e��Re���F���וo+?R�R�]����zJ�M���U�7�>o��SU�kf�\�y���5h��k�Цigj�j�ڕڍ��ڗ��k��~R�wZ����xTx������'8 ��_�����Iڠ3d������Eƍ �"S��Z�bS�i������9��4�l�6�3'�o7g� ��i��^�|k	XD����j]am�n�>h}����X�e��0�EQ9\�//�����<�_~U�+�S\���b���K��W=�Q /�-�v?�����^��������d���@��'�J�V�*S=�z^���*Zm���3��M�c�&S�G�K���=��[��������x &Nw�n�.0�CW������ڝeh1��b�q ����y�{�Ǎ�M
S��ʴ�tvѷ��)˜c^d^j~�����-��B�<���'-�Z> �+�:�z�u�u�C�ۭ/�l�c�܊z����C�ǀ�>�/_<���N�k������Yy�Izep��g�I�꫁>��f�:��g�f�h�����*J=��Tu����'4Ok������k�k3���u@՞�n��	a8�[ �:u� G��~ �š�޳��?�_�k�&�,�jc���x�x�jӣ�'LϚn7O1�̥ #4��6w�?1��� p6�X�� y?��_�!-˚c-��h���	T���2Us"���$�{s>-N~D~�F
�r�b�b��^�a+~�xZ�T E�AyI)�`
m*4�.�⤟��U��Q��T7�쪥�Z�]�{U��T� �sPu\��J�N^�)�^)��߫m���<���_����T��l�bm�v�����.�k��kպu_G�-Hz���B�<���ӿ��v�M����J�#��p��e��Fc>���0�s�?ǘ& ?0�d2�0��n������g@*��t�y�y��p���@��bN�L��Mn��r(�G����ZnuZ�l�m= {�Gk���b�#���%�(�c�S�/��+T�&t�0P�"�U�*��	d�?��Vݡ��6��m~�ῪYl �z���Ú 9��|�����
�i��X{?�?h��|V�w� ;�AJޭ{Kw@�3�����ظ�а/�o�`��,�\�"����?�1����!`��3N ��d 
��DD5�G��_
��e�t�i	p�� _~���ኺW=D#���[��i�׾t��I����S{A��v�j�º����?bxZ�h��0��r�kƷ ��My�W�^0}m*4�\-�� ��'��v��Q ��Uܠ���Uy��1�}����<��~�>HD+TU��*��Rūoܾ`��q.��w�_�F�,�y���^�@ʬ��8�t�.��� O����m#�z//���y�ņ�C�#��W=�aF�/��U��{����e.19LN��<c��t	���/o2�@����g�k M�,K-N�S���o��iM��߾����q�kַ���Z��8���$C�R����7�S�V�@�@��2������B��u@�_��w���k
�LLQ7 ���E����0W�#a�Y������k��S���DW�l��M���)]:HZE �>XHe����EÛ���a�Fe@�U@�3�w�֘�L�fA��-�n�8�x��-ˁW�r�a�)�ER�(�M�[���B��P^*�����d����+�nW��8��8�� �4*W��o~��!�/�(�:ZGOη���W�����?���*�*WU�jT�R1��A>yO�89Q�VW�,<
��
�]�G4�k�ji���h��5��ڛt/���o�O�/�;��i��	d���K����^2\%��h��%X�� e�0�xd�i��ƴ�4�<�<٬0�癗��A�{��,�*��0���i���e�5֊P��*�Q�ھ�~�{�^Dͅ�I��L��:��r�¦خxf'h�J����Q���(�e�M��q�xZAk� �4���5�%*�3� ��a&�����«^��P�`B��)�,׬�<�٩yYӡ9��
�̿5F���Z����c������]�K�����t��ͺ���N�>׍Џ�+A6� )�]�Կ��n4L1���n�ß@
�h�Q���Ѹ����F����9�=��/L5�3�7��OM�f����o�����o�5G[nL�bɰTZj--�e��eK����pN�YU���L��e]�>뻰���""���ˑ���+an yx��cy'�e?�)�^��X�(UT �{`��	�0��ʩJZ�S�P���*Wn��\S4-�8�.��%�<��}�����g���_��,6T%�x��VU��NՠjV=Fh�G�OUgU_�P���D��j�5���h���~J�'�9ͷ�K�۵S�Fm-�U� %|���"�P�X�Dsu�tu� ��Lw����^�"Fd0�B	7��r����[�p�� {M7n ��	����5�4ɔi*3Ղt�����G7ǚ���7��Z�����(�P�$�
K��n���@tGA��d56˱VZ��#�y��oQY�?Eh�M>K� ��9�����F�$�\1KQ��N�IqH6�+�??\9J�0~PyB�)�k�E������L����'�i�z�J���t5Ⱥ8�T�����U}'�cf��|���ޗ�EU}?P\L�05GCõ�af`d�7:(�[n��Bn(�Kia@9=�l�V��[���\Z07�T4SJ3+�AZ4�����9��٘A���������y��{�����.�	����;%��~<���n�3�ER��>Nړt�x�%���ﵧ�m!ʽ)y`��%?Nz�#���d�7� .ܨ������ӯ�?�UT���w}���Rz�w�jʛ)�oq9�:C��Eq��S�*UL�J�,��
�ܜ�68mXڤ��ӞN{>�}��� TB�:Q�����<�g�:�*��U���.�]�@�#��n��;<nZ�|��ƽ�����&Z�K3H��y������4g5��g��vW�z��w���L�0>�8���J��_Oؚ�EB�������E�ŉw �V��|/��O�&�&�J���$�(V����A�V��Z� �C����kWj��� ��]�Hn�lZ�L�h�D��dk�%���R�Y�[��S���	�^�/�3`k���Y�E�������ӟ��:�mJ4P7!%'�
��oߥ������>3�35�Hm����vt�T����B��2��3�S�i�r�^N{=mSZD�?c��6H0���3ԃ���ϩ_Q�zoSqC������'b��}<�-��{�"N�����k�h�i�iT�}�� ��/~U�s��o�?�ؤ���	�	C��.^
�iU�	�%|�p"�y���}�'��'��X��'�Hb}��ˉm!��֤��@�'-K�O�����M�v�ɺi ���^�m��ӵѷ�w�������W�m�z�)}��V)z��F��RV@,����@��Ԇ��![���0h�mc�"S�`�oI���ԗR?O�>5"�k�)͜6,���{Ҟ/�wZ�	�����Z�֪G��_�^�~[�U��� 8�:v3Ĥ��"�ڃ�]z�Ÿ����}Ws+�x�F��K�9M������(���(���x"'!��#	N�H[&�K�x~&س�A{�[v6�SR�$5pjQ�B�W&�B��'�´1ڷ@g'�N��|G��A���]����ҍ���
t_���o�~���������c���,���2=eQʝC����L��}�����P��+)R��x>����Ii���צ��&�0�HP_���d�:��ꎱ�k��3b�c߉��clF�b���^��������-V�j�/�g�[%DB��N>�5a#�ew�_	���7WMK|>�e�x�$O���L�V%.I+�1{)P�M��mm?mؖ,�(�v��9�Z����y$�;����|9�z]w��$�+�u� �v�Q���M?G�P�u�� ��Y}TJ�Us�P��J����Y�锎�8Cؘ�k����ʫS3Ro�r��`�M�	�A��Q+՝��!bU�w�
�Т�Q�SOV���]R�|�{�[c?�={>���޴�1x�4�3�P#i�h��#��,�����Ǘ��>�r��'ㅄX�Q1aI��	+���͉�ġ�������s`7�&uH
RY��~�V_��Vd_R���V��Ճ=_��v��J�M��\	�uw��:�n D�stuKt6��ހ���VI#�J�M��`�I`�����V�{��)c ڸ-�ޔ�)O�D�A^S@^ǃ�9��6p��Ӡ�к� �2/uY�=���7S�����Ȓ6b�� �X�v ��%�5�V�2գ��̅��%u�؈�������w���|��bO���3.5nx���Ҭ�{%nw�!�����l�(�8��<�j�Z�	�/�1��]o�r�4��wJ0EoM�eb]bPR��h�%���Lz,飤�I�`?��K�/�>�ސ|Kr<D&�%�I^B+n�@Vk�3t-um�r����I�g!Z�H�EW��^�K/����`�;�47�1|	6�w�2��dS��f��}.uOjpZ'�d9i�=�v�q�Q��荠�
�w���/�%�H}P}X}R}YJk$���ľ�p����c[�E�)�]n�����������2����?ܥ9�w�݊�'��:�Pf'T$�^Mx��$�A�z1�-�+��%N���E�)�oR,��LM*���=��9i;x-_&%i��;/��j��~���7yh��d��H���5�����g�-S�WWb�װ�����s�������j}�0�"�-�5�_�nH�*M�TP�E��H���Wջ�� .⵳��b��r���mk�N���5���f�x�[�f7����a��;���gǏo�n��׀mF�Hؒp6!&�
�{m�W���{��o?h�v�ULӮ���$�H�%�lr�NKr4H��[�{�����a���)�{������B�cSSL��f���,M�'���SN��M��iP,�M"��Q���xd}ꇴ�x|���p���)��W���rQd�z�{�u�Ziv'D��Sb'�N��vk���?cq-��ĵ�Sō�~��4]4�5ɚT��x��f��z∟4����<�!���A���$�>�΄=	q�Id�j�/N'�.�T�t!��6A;Hkͽ��o����'�����ɥ�w'��m������p�u�B�bo��� 1Z;}���~�[�@w�H�fn�S)�����	���S.�$E���N3�>��ڦM�I��y	�2�sO���uO�
��ܴCiG ��5MP+�h�U{��nV�z��/z-�zL���_��H����-��;A�3�+�Vgqm൸q�}�/�8�}�o�_���%>>�Z�)����@��v]BU�%��;����8 �l�:��m����� *�KI�tcR_�}�B�u0IІj�h�k� �M���urr2FY%oMޙ�urW]�.VW�[�{��`}�>�O�~�~�>5�u����2��p��lx��2��o�u�� �lI���L5�}�&�+p	N�(u(ط"�l�2�@\�u���ة_l\�x�v��=F; �q�qE��W�m��w��
�sZӌV�GǇ$�H� >�c�5�'`��%ޙX�<��(�Ɓ7���6໧i�joӖj��>�]K;��I�@�"R��h��L���֠}U:���~g	H�z�6]g�9��	��b�j�i��V�����w
[-��oRZ�$`���֐nJ�IM ����^ڛz4��T�/>-b̑�S��=��b���/P���������IO���������,���ǀ�6�V�~��� 
"zh��ƽ�>�dܯq��R4F���Д���$h���N7Ǐ�Ԡ��	�@OMI���D��	��vK���>��Ĺ��+m�����t���W&�$��t:�r�N����"�����?jÒÓc��N��|;���䗓�I���	�+�N�3�&�C��\��nEEa��������@����~	|�Ȕ^)���)�S���J�I���CO�0�k��cx����i�:	����so�nM���Lj���i��Yi�i7���/�N���<�<	�䟲X����]�L;̯[K8�u��6��Y-��"�)(_JPG5���k2V=A�G�f6�ۻr�OS3}��}�����>�������>�����d�[�GVқ/���.fzڞ��6]7�ֵ��m}�ew���E%�
��y�g��N�={�U5�@5�t��h��4,G�'�o�aX��V��M�7���lA�������żYOׯ�م��o����[O刢��'�ٙ��O�0���8��-A���g�2�����
|�&���ϊ`"ޔσ�q�R�;*�B�W��U�����e�`�|sD0X�<*��pmA�܄9�1��N
����Z��/k��Occ��������A�0��u�{�K�n����;�A�ʖ���W2o*|���\����0?�d4���6�7`���0�OX�_�J;NX^�>��e��u�{\�����|z��[�P��x�@9��?���s|1�/\����%��J����q&&���`6�3�<���<g��,�#���<�~�:��}Ɗ�4��?����r�\Te���i*���u�oY����y�ΰ��^!_����z�O�<D���be�8V�x��?W9X�6�+*CN���,㥨�ex�Ov�	�/{��T����/�SYu�Iv?� �Kͮ��z�4^�a�U��u�-�z�Vv-(9ܶ�����?He�	V���]�Ku�_�!kّ�y��T�ǯ�.e턥l\Ue�z+W'�~�CT�����Þ��x������e�>|��q�ee1W1�K�Z���m��8]�����E��p�j&p���e�v5���������8�y�c��=�_Վ���3�_\��?�Ju���)N�S�|�z1+�Oޛ'�����՚o?���չ�~1��=��5�c��?�����xm���3`��gU�-/�'l�β��|v?��V*׬e�=��~�/Lde�"v����v]�+O�bp����[�~���\^XYq��K9����b��*�]������U����?��g+�u�'Xim�ʊ)��y`�׼�:|���x�7*��d����WVʟc����B%+GֲR��(��w
+��R}#+׵�ϻ���֕Lo-k5�����F�1+�bX�R�2E�A��Y���z��Iv�6������u/'��T�_ˮ+z1x���u����nfe�_���"Y��:�O/�~UL�j�wd�{�ח?�Y'���r����"����ǔ��c�S�R��0�ʵX�̻�=϶ͥ�X����F���W�=De�w�~�q���#�n��5�����r���`j���j_Ŋ��}�������\�������?�ʥg�9b����3?���κ��&}�n�q�j։�O=�����ʖ;
)<9gОչ�Ώ��m{]x���e�K�h��E��8��w�/���2��c�G�<~n�:��I7��+{u�K=l��j���v(TL�c+��ٱ�{jO�������?�|��мݟM�헮E<�g��Ĉ�R.�\�f��ѷ?��������ͽ{g��Z���p�����b�~h�y��UK�[���o�t�?:��������n��uZ�\v?!�|'	n(
z��;�*�:X������<�kE�I��u�v+������_�ڂ��Ek�)^0<��]��x��m�w�Z�-(���y���?�~�����?�����V��g�J�\�d���m35����8�#�kkV�sUMAhz���=����0��p_�?�;���S�.+��x��)�ت���y/>�r�?������/Z���_+玌��vO�6\��R�QE�ԴO�����Z��|����K������>I�3����k^z�tW�y���y79�/�3�ݭ����h���=���u��o�O�����7?[�(����~�n󭯘6�cH���=-���~�����O����}���z���S�ؤ��=�xa���O��:��d�������Ǫ_Vm�x[g_|�KycB��s4��|��륷����_��_��|oKW�sG�s5�O����Vz����>�rfO�꽫>�䦙'f|��?ּ�S���,)*+9�损�ۚ�s>̩��ώW�:��-<7�J��}~��9��xi���w����%�k�^��V�{�`�m�VM����{.o��u�������u}tΥ�G_��z��߽sJ�C��B�߬	�;w�GI����u�g�(W�x.���æ��G_�$4Чׅ���+���X�e�����k�s���~�h���x����n���{�]��y^v����2�!�"+b�8���BZ�����ÄVB �
�^o��^�
w�Vp�5#�o1�
��!�w�W��/�^X�ૄr��C9&8:��w��$
ӄ`�N����Z�y�#o��7^���"]	���@B �y�{���^���<��M��J`�x^�~� �%�0��g�0��H��Nq�/���x��#�%|�Yxa4�� �4���9�^���2��ky��C~��e��w���G��'R̓����:���E?z���O_�G���tU��X$������?+8^2��~�μ���#;2^����SMw@|�z�DlX�b�YLx���4�.�g��l:�Pʂ++�Մ�Qp��f��KxrT�T�+�ܧt���)Px���Y��3A�
�.���A�m��t��Tx�I�Kͦ���.�L1+`S$􇞰=�<�u�+ţ}�[���"� �yTΆ��3<#�;ݙ�s�TP������'M-�S�
 놧PMF��Q�\g^�yS��X�?���8�=���Ӡ^)ܵ�WE�3��Ocur��gx��H�ʡّ��2ӹW�g$��<�+WDx��fz=ˠ��/�e�}��6؇����e�Bv�q~���Ɵ���]G?î�y�+#�������	^p�7=���ڶ�Z�wz�ޚ?o�<�����em����U�:7�$���cr�]o=�%s��a�o�p<��Һ���;���'����]��>a�B����?��%^FX�
_ů��u6/S���,�Jx�W����@��tj��8ME�^Dg�M&��OUt=�s�L�������ózɋ����C=8���+��ͣg�r�Kk��I��U [����|7�C@�!7��RӰ?�S3Húe�
�+�Hs�p+�9�N�Ԁ�2o��3#��P���k$MѴ��WH�Y����4�:�o*ԞF:�s|*���ݛ���eBS@�{Q{BZ�s
U�e��{�G�crt�e�b&?��2� ��c;Xٷ��/lge������6�����[��׭?ee�Ȝ���8�QD�)����65~P|:�a�ĩ"�>�ts�ُ�$�����N���d7Z����!nn����Ȥ��R�R���E�ݢ��ǡ�_�������xi��M���Ɨ�m�"��P+Ѩ�[_�dpb�gH"��Ԣ x���5e�l��$o| n�ী��?�k�����W���i���㞗��iS���/�B#=Z��;���l���?yC��~*Pw��8�c٦���~�q��fu�����$�<���N�{�a�n	�9f�x��"��l�����[z���*���f�o�g�����y���������� �x�?x����"[+O�t��&�t���!D�t��E����w�a}y�^O]�o�����)$����H�7���ќ��S�{Ґ��s]��ײ{��ԛsTt��<�%d:�[#�HwzbՔ���{7S��%�=�����)Pzz՞�=ǋ�pq���iO�޸��;�d�]��<���,{cTc|'�ܩ>���w}�=c��׹�ς��В����4�Q/�j�5F�a��m�a�����T�\R���������)�	�����_wc��^���w�~(ޯ�1�k}0P<�� +�?�rk=��+?�������q����K�\͟ց�e�YՊ��x��-�#��3yY|Ǜ��x�;/�8����u	��=��;���,�Y��n���H1���������Y���&��eݽ���Ɖc��똉�l y�*���x̵���˾���F|V񲖗!�t<�w�߅�<��[��ݼ�ȊM��|�nˣ�Z�\��n�s�r΢�S������>W��x��?&�Zٿ��B�ԇ1W�U��+�ǿ���@��Ӧ���N��1��kύ���Y������v3����=�l��h���ɲ�Xߟ��o���ǮW��ֿ�z��5�����|�Us�s^e�'���,��W/� �Xoo��	�����\�ӯJ����
�'���K�M�@��2>h�G�c6��C򕇆5P
����Vw��l��/�O΢�D��=�����K��S�|a]I��~1��d�������xC������ �>}��^;X��:ZL��3=�{��M�;�n�2���D�R�.��BA�U�تF���T豄���#\�Wf�3!>����>����b8���aش�{Μ��ɴ�1է��x���{�zC��i�W��bٴ�i�Oc��apr��ӟm��Zs�,��ny�}��w+����3��c�+0�֔MM��,�>�"�yM��w������U�Vۗ�]��]���צr?<=�Q�-~�^>��/��������é��]���'�r��x^�^z�#�ռFv��WLg�M��i�����a�άn��U�X���c���uMA�vp�Vf�a��Ȯ/i�u�V��cy������0^:fr�{+k�u~�_��q���2�p�;xy���ΰ��߽���1���e䄦�丆��o�u�7�C��vN��_��3�o�������+$����m�\<��xh��+뇟J����o����;��������/6�<�6�>������4z��~�k����s*M$ �y�sڄ>93�״^�����\�@_��k���a��}\�3J�k����Θ�����[����]po��S_6��,�Sy�i�O�+�VOk_�n
}|c�k}�߆��k�r�����{��d��rV����n���27<����s8ry}޿��]Ը=)��S�d��?\o��*����	�L���������1G�K��@z'��S�r/W�r y*Y #�+�u�,� rAV�����"Z��� ZŝB��eq�����;yZ�9��G�O+����iI1�p�<�1\�����'��Z=����Q$OS)Ŀ$�^� ��FL�e���F���;�[��Z����7��MX;y��ڲ�+�|�Y������������c�Jc�շ���N���9��39����wI�+����h/���Mo�KVK��R�3��qf��G�Q�;��?�d��Y�*���E4�EĹ��4f�e?�w]B.e������7]e�v
�����@�|�Tm��
������y�b1�����I����}�:�������%4����z��Z��R�t�5��)=^}&*���ᠣ2���y��o�/�h�,�hnur]���at�=ɹƑ���\-e����k�=ǋ+��ja&K�8���GA��qhJ����F����˨�%O�<b�C5�?)����o裦��o����>�'��'�Q |�)}�����|_���kj�޿�5u~�
��L6��W�Hf�)����ϸ�J����<���lɮ^���J��?��2熓~��8B�Z����[��[��}�@���z�\�e�v�����>�PU���]��߶����P����y�ܰ�yp�0�vSJ|r��C�@q&�=�F�hW"��aS��SG���1V�k�/���^?�vz�;�8��L���ׄ��'x�r��xֽ�,�����*����n/Q�{ӳ�;�4J�����o�i�
����Ρ�8��Y���=����Lڡ�`ky��rN�?���tK���s��J�I�oY?U�v�~����u�|�dP��i5S�_?�}y���W�oM�U���	��(�ޘ�k�9���Jo~�UO���C����?���_��&?7&yW�k5����o�� �K���?�����}|�o��z��X�;���X�ܫ�&|?M��4o����>�����#��w {"����:��>E&��7lϼ�C~���ڳ6rT�#2�Ȍ�1��.�`���6��3���H��EP|��|z�w�V6}鞙��ס|n�����2P����=>�Ѱ��f�t�����h�Ԁ[3��L��w%���{=�x�M�M^-<wd���6U��	xW�����k��^S�a��H�9M�?�0�v,gK~���&�?�x�$���28��M���>��=���y������u{�,���m�>����`�Y�Q@�aٵx���e�<s]��~�������vRex���)�����W�^L�3��{=�a�4�-P�M]�������@=^��k]u�Vz^������_�w8�f<���@���O��S��{<ٴ��9��'���1z���q�؝��1��A&�J��x[�t���=����+�%X�۾S��0	����v��k�0�!P�����;�u{��9�A/�w����?
����̍[/�����8�p���<���i�.qq�|
�q������<�줩��p%�����q�Y��Wf�YW�5�����du�L�{��?�x�g��d���O<��A�O3���=̥��h>��ᦙ��Ｌ��y����{��@����ɭ�|1�>�����<cy��L^��iZ�
��^�ob�j��/�ߛ�.R^�⥶��D^N�eqە��^��m"��8��Ԟk��煮��?��|�`�2r;1l� �kȚ�� �R�7�Όi�������an�?�̰L�<uQ�̢�Q��c
�ɳ�g48���s�5���O�,$�����ZH.Q+,r��)�"i�|�v5ﻖp�K\x�O�cC���r(e|<�8j�+YF�E�J#]��#��b��`��C�Zd�(�Y4y�̂+�������tw
�ʫ�#���1xRU~�@>'�?E��3z�'����<)�}z*������2g���s�͚l��Xf��Q0k����UX�,��)���B����O��P��;�6/?��:��Ҁ���9/SR��U+��kK2+�xY���#�߿�F���~����e�����f��¡Mߑ����A�������kk�w�����s\������7~�dg<O��/d�����F6�=�l��S=�gQ��.k՘?���JoW4��F�p|k5ֿgTՔqzֿ�qz���8��7}<���E��&_�Y'ٷ6q\2��r������/W�>��Г��a�ʐK�y�켭��F6����{�20DOxł�v�4E�ߪ�T<����C��j�z�����G��x���v��+�+�~���iv�zk��Q	_|���-?~��W�4e��w~���(W��pm1v�����}^)����#!����=���,���:�|1�{��i^�?3߁ߗjl~џ�o�[	j�~����ت̕��|���W�O�`+�!���|���A�!g5<���K���=e�\���]�����ο��{b�e�J��>��,a�!�k�G���@��f`~�2�+��]	���#�O�'�����'�{͐�)����Ȫ���`9Z��l�{�M�'����t�1��4@Y�\�^:~<��2�7C�}:õ���G����w��j�%0&������א.���h�%�'���Ә��?���/c^��OڇMҗc��s��x_�|���חՒ��>x�r��Y9�^��~�ݏ�i�T;��9��ge/᥷&|B���|�#��e��[<���#�e#EJ���c�]"���G�ur)�׏�*/>x�E\�X�.<�򘋅����^�B��	5�o�sI���s��~�H�X��ϧ�)꿾�WC)~FS��@r��_}���"�������qb��u<ϻ���� ���n�r+K0�_<��NL��p�]���b�����ܮ�잚��㭙��_���^���_xǻ^��\n7�r=���������ݫkח����i�WkO�~'�������z���{M�;��J�H������v�����;rLq5�,>)xhw�ܾ+��ؙ"$�ۛ��m:ԸZ(�����{X���������s�������볼<c>� ~�8��1���f��SN�+�Kw�a�Ƣ^��+��n^~�ԙE�����>�mBt�h�FG����B�9t/��f�h��.�;���*�2m�ӹ�#k[�Ys����\6!:~�w�N�����P�f��R�
m��l�;K�a�֎�r��P���lK�2��.�(U�/~<Ÿ����M����n&�-��N尻�N������g����j�>zW�&	��CO�p:7� zج�as��i�������=�<<w*w#��\��� �Ǿ��P�LM�f?TnE�?\J��L�v頴ǩ<B7��oA��,��"4�jv:�� �6(R:j�*m�Wh�Di9#��3ǡ�
�b_�d6K��R��,}�������)O�q�q�q�'�XK���\S��='Ju0�p:��Q�~�_�%S��,�ChZ�t������N��qՁ�t*[�;�LR�%9�'�+m�~U� 4/��5F�R��} |iGQ
�F���tZl	�A'��z��F�����$4J���AE�qP?MS32:]�vgJ�:����2x�a,r��l�tʬ�nU�l�qq�F�l�Q��Y,�E�����`�Y.�b �����eJ;hJ�?ujv�����Q�=�B����@�����i�-�uf�	�(�PjQ
rf�н���;�Gp���݈�/D��ƒV��.�Z����1������6+J�#-t������8����f�V�+���AiCgq?x�E� ���h���hm�F6ݬ?jM�f�kW�������7ZZl%Z�ɾ�bW�9��D��u���;�����V�y���G��%S����R�D7S��5�q{�ג��>�ߏ
!�^,���N猝C�JQ2G�r�o8r��@��X����@8���wep�Qq/*��DkG���ˁ����R`�9����͜���	I���j���h�>,�8V�`�Aa�����5�2��C��@����E�P��@�����GO��N8-�tf� ���YL�h�2P�� �%����IƉ�	�b�O��p��ˬ�h��"����73nCR�k�ȟ�7^�G�>�-}6��!יAWE#�	�f����lA��b�ɠ�o�EiK��Na�p; �f�u4J��}Z@��,6K�*g��1b�O1��E�����F�&�B��⾢�v'�U!Ԑ9�+`���W��BJ[Շn��l}��[cr'M���,m� c2��S�Jd���q7L:׏�0��= w�Nks�fұ j�W�W�{�1��t
T���Π�@u.�+�ڠN�Ң������.J��ǂ�/�Dʂ�}�9g���؊����S��>%]\�TNV�o/-._�2�u� vk�(uY�.j���D~�}L�(U ����d5�F,�ְЩT.Dօk�(���	x�[��?�y٩<x;|�a:�Z*[���cA��oMwq��B0Vŀ�B3W0h`8���p�tJ�N���K�����#�:,�ucrnTiǍ�R4飡k�f����AQ����i��T�[���.������ ��j�p*S�+*���E)Q�/�.�Q,��D�k�oo��i�t܀Q�G�t�+�JC�c��o�b�E�&J/^B�i�#s3�m��l[F=���<\��d�P�G�UQ��	��<0�Z2���a
��(&m��gĀD�dߡE�&�����v*Q���;��oH�P��c�'��c�r�EUc�RI���q'�H�!@��Ne�;�*`:���@����3�N�v�6�j@�c���p*w�	��f�eG��s�r���KF�O�H�F^��卬%o���+��@D�w0�Y��_���u/�S���f���VN�pU�=Wn��T;�����l�c�)�&��,0E�<�X~���9饑�1����>�_�`p�E!J���}�EC�����t#<�F�f*�g_�r��O0
�5Z��٭�n7�*te� � � �+�sK}��'�Q}��1Tc9 ��V�bZ������'��E:b��C����4K�fې��ʪ����rDn\��q��Q@��`�(�[��/7B7�;6�eNe��;�*�^L1�Zk��<����N�R1 E*����m��O��� ��,a�K������fW&N�?�{H�1��w�-ݭ�����}�@6�����y�wa���+,�8��0ґ���l�3����F:�J����7u��%��� �]al��" ���6���+8	ӱ�3�F+5ϸA!��A�� �8R:lZ���bk"jݱ��e���~0�S�G_[�{�vL����8D!��̫D���c*;]��E���N�x�3�ͪ��x�t+R�E��7O���^���1$b8>��4�m���4cE6sby�<���0Շ�)�����m"�X8�u0
d���f���>��1����B��C���ˏ�����:DS徆1���a�c�T"��mA�>	��:�"@�:T2@�>\Ř5my��>L�|*b�"x�~sĠjO_m��nTY���� ����1b�\]��><�l7��"��G���F��4b�>TF.����l��+7�G���@�2�1t�g4@�A|3����=4$�cm���kFqΚ�0,�[D{�W��8"��G2`0p�I��X)®,')	E�Q�`c����	�V��BDb�h[]F�o)a*;o��@���uѫ���TVD/�&���R�5���u*+�������4'ҁ�x&
��F��dR\�tލr,�`�~C��l�#B0�G�H[P#�@C�3�7�n���˂�"8�K/.�8�,u+[;C���މr�)�%��HI=q�` =���z�E�̒>3��;�G�2:GDշ�H�����!jrx.69��y7��;��cP[v��ڞ]�T��;-�#��5h:r-�XQڎ=8H���w��pq�݌��C����x)3f��=3�؀1���vA^0�Ou��c���+��� ���d�j�q5�ʈ��*���gU��Jf���N�K�tm>�&|�����)��T��tF�_�t'�V�&Z]�s��BӅ�z���؞�����6�>A}��M.8x^6���9r�q�4q#v�G�~���;�ۓ�@��Oբ���Rf<pL0\!��;�"D�py\��P�E6|ދ�g�A�p�5Ƀk�C��,�y]�]�<W���`G�v����	Ƴ�x��܋�Fk�OW�z����9��V�+)8Q����|�Q��q���@�"s�1b�Y��T�Cl\G�\��j�o$��*����� ʅ��2������)���9l�~:�Z�Y���ܹ�vv��~u�JMɹZk7bl�Z�WP����'8�� ���dX_e��t*� .�Ð���t#�'���k���.��݊��4�5���#E��X��V�K';a@3ע�yVQ��X�X'���V����Bt*�W��L�>��t�v�2�kXA�!%0Z�t*kfњb����W2ރ'���i3<���j�Kf/i `/�^���]^V��>��;.��}��z�R
{�Z���D�9���"�jB ��ΐt�^���V�����C��-�|����0qH?�=�
ܿ�q4�Ί���9D�j���^� w�����a^�4h�E���W�")p��(�q���#L,�%����qK���FF��i�Q|(���-o����G�YDT�d�����ⷉ�m�bFY_�CG������hID&��/���΀��紆�t�w��M�Ezy�KGG���2��z��hѸ�� �62:�b�2b@����l�j.,��Z��ڭD����J�B�����  ����e.}�i�L�_� �w����3�b��]�Ў���Y�u�?��"Ͷq1���b�⺎r&D�̽�IEý��-}j��i�پ���y���n�ʈx?D1���f��%�R���J�X�{J[�������?O��W�J	�U���T����vk�hkhg\���h���S%����gK��ͽ2XT���?Z�W��l��5��`��v���کf駤��G��oݫ������*��Z�~�D����!8h����G�ں��ՆV���H��v���N'�����}c��4-Ӷ�n;�K��>h!~�f?���'�թ�ܗG 0-�jg	n�c�Q�#+�N1�ס���8r�� �������h�I�7!~5����ўCb���ʨ�!�_�A~&�'�s.Kج%��u���1Mϲ����7���q�-v[$�� 9����X��;���:��_n��`��A���il(#�a�6 j�i���t\
�[�0�$J�;��p��\�C���=��q&�E�V�fk��N�)�,e�*w۠F���3qA͌�q��^��<Q��<H�|8pDM��h�b_��ݻ����p���섫Z���������,���=��E���@��O�����0�>��Z$:7���1�~i���iZ��,U����W�x��?�l&\��F��c_cK��%M\�iI��Z�G��<(_���KkGQ2��N�nM_���
���ud61�O�F�+�A�^���J�ʵ���(�Q�� �5 �FZh�+'�"��� cF��GmV��F�-7}
c0��&��Ӫu�#"k�H�ɥ�]�t�?RF/�=�H��<��<
���sU����FiD9=�.� ^9��E[����7�?T�>�Nk{���$U��!�s��>tifx��/ۗ0�a��]OM<<%w�,�Fq����O��>�^�~`��ʧ��a��9���A�*"�O7��� |��he `2m@��DK�3TXۼ#��Q+k�YK��z!���~�B؄��h7D�w��m���(ÛÍ��h�@��iM]�(�yh+�'Å-��� .��-��V��b��:�v-��]��w���B[��tnl��$���q�	B}�X�#d-���}��B/����n���<7�?�]V�����殆����Ëz`��{�O���5�%�s��tOF�i2��D��tPX[P�6�n�>aJÝʍ�Ngy͓8��X�����IZ:�b��zBQ�%-h:�� ��H�h��CX6/�3�� ��@�wB��������7�(�.ě�=��v��8]_+!��+�����8#6�u�L��r3ky;���[V����Z�Z��ky��Lǖ�r���%NV�� ��0�f��p�:�_k����]�cqI���$�9p���
|	��Uڒ6O�l��1��>8ʩ;�V�J�q&̡M�Qs�v�7�%��t�=�Hǳ u�Ы�7���d���t���QF[�1#d��HZo��s���{}�S9l���T�9��I���\��0���/��A����������
���ߐ�&ܜ5��(��)}�)9��,�RO9��:�.����ø~o��QE�At-��h7�g"*���&��V���h�wd�BH^]�������,��&`�G-v=�1�[�E�3}ƁN��6��qPD����ֵ�U,�ztF����ѹͽ���$Z�\^�urce�����ʟ�	kH8`�f�p�$��*����3b�U�V鿶�c�*��¸��n�����Qq���#*�c���Έ�A��i��a�4귗d�����GqS�{3Q-�{�n�
8La���2SHa��2���U!���r�x��ė�y�Mؠ=6�v��Ռ�p����yƥ�;����`��R�63�3�l�7M���P���[غn��w�b7ފt$v��n&A7Ę�,�9oU�zZ��Z��c'M�]K��"V^O�ܝXٸS#�����?j;U�Q�#�a�O��,>e];��[iw�gJ��VpbBsf ��-X�7[��aIN�[�:�3���ʄ�$UoD��X�kp�l�-]$U�� ��ڻ0J��a S�0%�</��Wp�$�~�.���Y�?GT�����ߢ�e��T�"th��%)��s�fh�L��Q��!�"��0�-Ʃ���[*���F�A����T��Ne�X6��������8�O���V����B�Ѕ͡Wi/��aԔ��K�}�l��.ДF�*�J���6J�B�� *�b���9jU
�)"w��^jxm�)�1�ZB�-��i4����L�b*�q�ǖ0�f4�W>�k"�#�����[5��k�xO�YNe�1����of�UE>��:�(VD��u�����s��>�N�G�gB��7 +Ah�O
F��; Nr�_�߷��^ܬJ�(T��fi/D��9��2N�ө\8�j��kQ0��I������iLQ����綱���u�c�Y�s�#���S�Jh��ͼu�l֏7���"Y ��alsQ:m�6k�o�H��k��|��@f��N2�r:��D�Y5إQ4e�i��y�؟0�C^G�'�^@&�E0~�;��;3:��2�@DWTx�����Uy<��11=;�%�zS@��4�Vy��OA}$WD��$X�z�(Z� _��w�֝h��cC���0�5��:�>|c,�K�P:�-��@�9���RA�2��H�sX�B޶��y�-�{���`���`b΢6n�j6��W6#O_	$_��hA��ۅ �-�P��4wG
�����:�Cs����N9�-Cq(C)g�ː�	�|	�:����k ���8��&��YL�h��N�Q�*fUj��z� l�GԖ�ƽ���^Z`/̩�	�Ts�rq�y�}���h���4Aw��qb������i6��H�#���4;
�p��1ݚR�d�c�'�]��H֓H&�م����QqO�q�q�!�+e�����]+��
溩q}3C}z?�-D���چ�.�?I��� �F�]4�p��p���\r��%��x����!�E�{�+��ƩLI�5ө�2�T+���v�>�N�>�⏅T�I'�N�9'�<O#�&�w�V4��z+�P}.D��#�r+�Y[K5��}3��̽���]<vZ�{!4>�E�b�jB���DBB�)EiLg�8���~�T׏�'��![D��A\����3�@�N�3q�5�b��ŭ������� �=��4�y�sd��p��2��ПtA�=Ϧi4�O��7���'x\�sXR�;AGD�M���p���J'D�aV��N����G���c�S�"6v���:Q:�Ė3�ü���r�V�\�2�\#W��j6ge�\sFH��7�"|��$o��ĵ��������A7�7K�f�V9 ��)Luat��[��[8^U2ݶ�r�����&}�g�o���u6�M�����Қ &+&�\���������B�P��:��#	��<�霦��T������ $��si��r�5�v]��g��9Վ?��"}æh����l�ֲ)Z�9E^z�؄F�VI����^z��bC~~kqѫ��[֩4/�Ao�.�K�od��꩷�&���e`}&N�
�����^���[���-�\UK/�/Pa�WY#��N��F��o�T7��N�/�/ì�@獉��K���s_"t�9)���A�*r�l�~:o߃�w��mؾ��$f<8C�܋�>����E��b��{2�zdI�Y���ADX��"��\3,��ԇv�*��XH�DL��\�5 j����o��5�:�'���Z�zUZ�z��Ko��`;��)�N�(�m�i��s��ygZ%��E�>�#`hW�>���a����[�c���X%;�6VWa���E�
�l����=�L��jq����0٤�h�ਣ���x��=��M��ybo���p�W���=�=$�_u���'�e$˸�ѩa*�k�WW��X�.����\�ā	I� �N���1�ZO��w;��~5��F��=,ny�l��=��:Z>�|�,��-?&K�	������W���,�R�:n_�A>��bi��>$R�[�m���Vo��S�3��O���f���;5\~�h�	��%:4Ȋ��I|��cW�9�N��LQZ� ߳�$}/J��?q�|���D��tj��OvVoc�o+ma������+��Dt�)���ާ��� ��.���/�}�Ⱥ�}������97j����I�Ԏ�ܷEr�����I{�;x澅�s�N}{��Է�n��&��q�WƔO-H썾�l�:�}��sQ��pʈ���i��BVG?�f6~,�:Ϻ�n��X������i0�o�Q�4mǻ�`uJ�ʟK{����C�N�al2��d�}T+ �)����xͅ��Y���k�*oܛG�^S���r�8ZṚS7a��w+�8_�\ߔ�
��s�F����v���Y�9_ڢp���D��э�W�t�|)���
=�`�R���~���W�� ���(�<K����_�|Y�#Y��0�ئK8�wmeJ���2=�w|ܿe��y���b��}���B���P`��y�nx�{7�)���W�<gr/˟/#>��U �������e,��/�t�j;K���?F�=��|Dk�t׳cL��S����e��"�e�M�br����4*b�Nu��3���=�y;<���G�ޟz{�5~|�?�5X�￹Z��ٗmp�EZ��8���,�[sy��nfo"ڳk3�� Ǘ9��hU�N��4�m��h;�������b�7��h��CT�\I,�ئ.�	�ث�r�m�o��~Ƅ�L��'SR,W+vU+)�Œ�� ��e��C^0�#Vs�h&�p�a�*��jz�#���wt.D:��<}�=f��D�&e��>t}!��A���u}����;����5�}����˾!�*�9�1:����) �}��!O�sU\�tyG���<��ҫ�:"Q'��g�ƾe�����˿?�ӿ?ؿ����g��g��a�WA�3/҅�t7����
���߇=��^����<���_����/ Xk(flo��Q��I������&ɨ�����	LN��ʤo�H�����g�Q_3��o�>���x�z�7�C�p���?5�=�@e����a�`�L	B�+xnvF��3���gq��&��~�NlgkߖPSīE�q~#��2	0n��%/�TҭY���M&9���W�AK�tl �k���e^s��U�2_��Y�ς���z�.5��NK���u䴌��}z�=Ss�"�˂Z5-3�#��iSߑ�1j�.��������P�bͶX�&�a��o�ֈ�������a"�ԱQ�t��0�{LѸA��Qz#�z�K$���D�����7��(�uT;Eo_v�X-�-�Qg��=�莄/i�^�/U��k�g�km�Z}��])�ѱ7�5��]���_�f���q��0O���K`�
&�^ �+T����l�\{���2^\*� �aR7�!#یb��"7Y6��n��^[A1oߩ|'�����A&�kcģ[@����J�������/P�rV�X��m{�e����������ֳ�������@�׾��e�XȊ��X͊�Y��լ�aE-�h�7�dO�h-T"����22�ob���WŌg6Y[��~�7��t)dr�E@�o�����Z.��Ҍ1��<\��8B�i4LnkfQ��xR�����I�ד���u�d-=)��rӤ�=�����j���<]��t%��,�[b���<�m6!+�^��5J�t��Źj�T�&��ߡ�嗅ң�T�����C�;�Kyyx�N斃_���43��`z���b��|�6$����`���^��ڱj%�KB���A���|ߵ�ڵ0�7��n7�&9�
N9��è��e��aA^�e;^{�i�+��M``�v��� � ��� _��C�V�?��D�;N�̗�� د	�c ��y������[�c���?�������q@�Ћ�3�ua5�r*@��  Ol@�����`Ѕ \��ÿA _\�2��B�l����d[��MM	�<G\Z���+|XT��fU�س-gi�x�mL4�;\���ҾX�S��A�ܴ�i+Y���0����b-Zz���6M�b�D�(���H겾$�ضʆ}H�ㅇ���Wx� ���D����s]I�]�%��s�I��_pZ�8�c���½b�OZA �������Y��!gق��rF�ô�U�$i~�o�N-���Ml�?��V���:�،jb3K���{��!�>���6���Abs����A��%�R`�Cȩ��z�B
9U�G�O���0�K�ſP�������?��\PG��m�a�Q�O��(��1���ᚽc���ķqKS`��30�G�|{�3�
Y3����QT.E&���L]n|N~
!�_A/?�|�����s� �{K Y'�R��A-� �a��T�%(�v��;}�	>�+�f�Ž���仮7�χ�N��G<���L�ω�7�'����_��=ɾK&�n��1��BL����|��1�#����و���+8� �������8<��+�Qq3|�&u7�Igp���D?�N�=��ەf��Iʒ�ws�0�(�ʉ{�\YjG�Z�R����MD�.�b�YG��ѿ�$`��2��Z���S��-��]E��w�M���c��x�CE5%S�Y�Lv���f�I��Tv�ENÎMgi���J�Gܛ��g���k���W�s�;�:%�R�;���gAN�n	Oʝ��ʙ���EAr�4�S�W��눊R���a���r)��jcי�h+�u']W�vT+�"��R�(��/gDE�]��Oi�Xɨ�V"��8�4,�:-���7�X�IZ]�V%�)�/}F�#��G�y}�rg*k�Z`L�3���v�����U�ym�(�oY��#�,��Q�q؋ �$�%ʊ��.��B?��~e w�eD��'�J�V��cOorǖ�^�>�m�g���8.] ���x������a�	fp��9���FU7�
Ƿd�0�[(�_ �4���k�jD$;#�N�(�LN��ܕzLx�5_᷹"Aή:�)(c�߽df���9H���M64{���F��]v�����s�՞�������%��G�����L[I�ٖ�~W8� ��N1�b7���"*������gS��)�m{��h�;�����]P�?;��$f��X�V*)���jy����z��Rm��.儧s��u����kx��cΏ��7�/����2��e���x&i`6��w�	tX:�	�Q�N��`����ȉ
��+i�C4zr�FĠ+M�nGO6��
Ri*�~����1PA��?ǌt<;Y���� #*4
��p���8�ۄ��[��Z��[O���c���z�Y�W�������*a�q �%�"R(�]T8�[{�h����@6����i����B�XV~!hA�t����7�1�W��Q~&�:���i�i�Ɋ��D��:��^}k9'x<�2�.�G��tEM�#S�s��0u?���\z���6疵�byڑ�j�(*؈�Py�;�"*�Ge�.���Y�BzB9�%v�s� �c$���?�}y|Uh��R�H�U��_���M$�	M�Ȯ(U��H�H+��JP�wq�T�O����eG��}B@
��;��;�I����{@����ܳ/i�G�#��/��%��i*��T6��h��/��Wr��&�|y�3B]�7�7w�x�Ay�&��Gl�w8�����)]�X0&e��&��� �xpwj���Wь��#��ݠ�=Yl��Z����N�K��W��-n�̋����x�W��SB��P͉�[i!�}n�}ɵ.@~n�-����D���*̡�)����z�}|�N֗VUQ��W�~3T=���o"�����9/r��(�w��;�ݺG��rs���+Q�1+q�X��!e8�S9�
G�n�(f-(�g��k=�)�宼	Y�o�������Sw���$oډ�R-֕����Fb�咆b�	�`XwX�U���77k� ���6]Ca7��ug�q|� �I0��-�;M�֘ٙ�S��o�l(�?̵��+ob���K�n���\�����l�B�+����Vײ?2�s�T�1���DG������	o�O�¶�;lI�ߒ�4dS�*�L�p�m�c~	����6u3ӡ�GjK���Fl��Ad41!�٫qf�^���ҧ�l��4rG�p ��`�a��6y�.��q6)Ĥ�Y��]�6❀��m��3?�	�Tɜ�v�].��K�P6���
Ѱ"��d��|�'��ՏP��Ƿ�D~�.��@��:�����-=�/�O�R����]a�x�m��6ι�Rw���)��]� ��1 gM�JS.:�җ7�P�;h�n໴����KO&���Ȫ�%u�C򸵪��!�����_���W1kFL����V?�����4�x�G�/��~���mb+���c/��h�ɝ�|�?�m
^�cڃ����m
\�)p�>c�3v�>c�c���s$'{
�w���n�Aԇ�o �Yr���� ^�����5}�7����|�n�̓{]M��/���Y��j�%Z����^�ߗo(y[wڬgԀ���Z�|=o}�ֺ'����^���6�����`�жA�K�km��m+ّ֑c����)��dЏ��Mf�:�eu2���#b�ښ5 �7���av��S�<�g@��nX��r6���+�-�b�JC�Au�k�NS�����,����IO�K�%��_��/W^D�ؑRF~�<c�q���q�X��m7�<�V������a�,&?[�'��T5y}Tzds�>�r\�PL��?8�^2��#E�a�P�]8�l�Z�/H)H��F�ŵ�5Ea�n�Cn�HO�#��౯$�4/��6�Km[4͐�S��++˯}�脻X{��S�@A��/�2a��i�4ڈ��n���7�g	X��`�#�ё�C�w���Zj�ӻ���MWq?��>�+J&=L�Og��!��Ey����/ʤ؂+�D�X\�7Y���xQL���G���n?��]�1�F[|�N�����^©�U�������#v���TY2���W}��|��p$�$��f��L�Gv^����Z����4Ј�d�-��[h��J���.�}xr&�(� �3�/�׎H ��#ؠ�v���O~��b]�O�U�(�N�ǤR|K!Q����vЃ���*��@��RA܃��^D�͵`�(nN�����V(����
t����ͤW��3���k	4>�6�;%��[:�go�K ��9�ņ�suɳXӯ�(E"�}�+��7�z*�Cnh��Z��y�&�/ޢ��ғ^�S�)n�!��ON�_m&5�5�4gz?+��^D0#Dl���G�.�p�ovO�S��P��][8�Z<�'i�0<`�� >�^�nA�o ��#Na�CeK���Цa�
�;���CW��غ#��=f+_�]���,Y	[yǽ)X�4��aM��r����6��>�>�O����NE��P�@��w�dqK�L�6'�+]ɓ�pW��|}& �c�R5>Ȇ� 짥�F��ɻ����\��}�@��抉H����\q���5m �U��$Hɡ�$e�|d�imx"���#�sw�XT�D�B��ުd���ｹ_Wh�s�Yr�)�����K-�:�
�H��ER���x���
eZ	
�k�>Ub�ID�pze�4��m�G��. �42M �Jqؒ]�%�-a�N��6��[�o�g���6�&vS��6e���#�ڔ]lS&eh�2.#ަl���.�m�##�)�)j��(d�n�lJ`u�?��F�������ek�|� ���]}�؍���ݸ\f�z��N~+BoB�s"���ҋ=�VH(턈	���~���H��NB}6�W&w�'������5��TQ��P��_�s�m���N
��l�Ӽ`c�W~�W*NbL;�5�s48�A�xUi攆����3	��Ƚ�\���g�A�J�o�a��g�1d\��8�Sn���g�����2��l��7�۝�E�1m��W��䷉8A��ƽ�0�+��3|j|���ԃ~�k��&�1epz���z��KL��O�0BM;���fa#z��8H@�w���q<lA�N�^��[�v�����ki+�\�Ɠ�~��6A}	�@��h��P|��{��x,y�'�9�ڗ�g���iYt��R��Sxp=�Lgq��[§s�z��S��8�{��[�һՅY�ꉀn10Rnq;M{��2=�L�����sN���wǡ�p
�(�q4�D����o�Պ��`�}�v7Y$y�5�ۇ
�|��/���L�
½�*��(��p���*�E��R<�\|I'��Ws�?�и�+�%˺r.�G�K�y>�	V�� 1�+���.��Gs�
r{�`��?������.s�1�w��H��Ʌx�sx���}�����^9jA!-����p Hm0 )�ua��]cՍαs��M|�4z2�rEq��4��@��_���L��%.j�e�Wr�s�G��
�S):�paR�_2U����Y��A�N�2��þn�*����i�'����Q���3���_��M�iTW��&&�e
Ұ������L���Nk|�1�δG�:�=�V`��`��9�#&�!�ñl �z�]��O*Ç��;�
g8��^Y��9�O���F��� �ڐ�7�J<-�A��$4t�I�nK�����T�t.ޗ��YЂ��th�}�=���v"�R����l��C��%O@�/ި+5����Fy*\2�]�J��O�:�����0�
ҿ�ƺ�6٫���.�&6U�\~�F�{iV���{ڛ�&�_��2�A��&�BjXe��9�F�:�%?��Y�m� _wf�L7W��8)�:����8� ܝd�S�r�p�2v��fo2�ߊ��N��O����A瘚@����TW|��A�?=݀٪z���ה�K�_apy�������J?����܊@�K�!66$*���)�#�[E��^�;&�;�jjgV�X�R�L9�^42c$� ����"7��7��̔�4�Z�����J���'�?un��҈���V�:�L�8
��0���9��Bqk�;��Y�Q��)����|9g�t�d��|{�����T�^�
FۃCV���ާ7g��,�+��M����V�!��=j��
�!#���kN�!_���Ψ���x�4�����V�;���a1���Ǘ��3e�Q�̳���3��	�f�`��{���ߚ_�]-������
z�"VҁV��7��/4��ϭ����[ջ@=g�]Xo1�c��	d�N^�M����+�,��/���9��������i%V�6߸�ȁ7�����%C�^�2�T�?Ģ��zE�~���� C�T�e*N`_�c�8W�vIN��"[4S��S�>� �t�|��6�?ы	�z�'�ԣ}<m�+�`-XrK~�X���|�6SҜ�U�PPcp1�C���,�=�QC�f�h�?fD�<���x�r���a��}��Cj�
*ܹ�\vx��,���(^C�e�����`��=�T��~:G6_�1�z��%�Ӥ�r��60��,�ai�~g�}9��k%�?;�e��=�Y2�d�,V�Ϗ��L�S�1Wc4�����bs��Q4h �d�I�)�ע�hpz��?G�<�/��c��8?��^v���UV.eP7��r`+�Ҷ���@��[�w������o�|@��g�>O���������a(���T��˩�ۄc߭�}%z��,7%�K�a�C7h�-��17��_���o�W<���C&1�m$B��
҂��� ���T�|2��"�w	f�>�]a����AlE�������7��(�EXJ]����h
�l��b��x1���5����c�C�HV�Tf��CH�R�J�<�Ix�F�x����w�8i#�gX3�i� ֖����6�T�)�^��\�!�u)?A���W�Ù]ϛj�|�e��jPրAJ1��ˬÅ��S�_I``���U�N���Oj	ذ��[8���u�9}��;�r�	w���e�~�����$�p�-�*�c����b\��V��\���q����j�Tf�`�-�o�ŗ�C�(��G_�����'���#��.��,T���S�s�T��qQ�Y��K��D,��
Zr`���5&��X��G!FI�:�G����#Ș��U�J��	b`%L�%?�!��g�>f�7��|<ԆG�,րI�4� �����r���Si;'V�g`���H��:,�\js�ڏ���bfmM�-�쪼�b��o�Y�Kk�\M�=:�C�)���K�O��&'�[�=���c\�q���idH&����#�(�*&4�To7	�u��@OC���%���f�EA<��җl`�1<T������ϡ �}�w/u��� U1��23�����x�0����f����!GL(~T�㇧Ɯ��9�A�y�A2�=��s ��E%ꏭ������
�Q]� �W9�'�X%2Y���W���Du�m��je�bWk,�W�.u&��F�aXa��k�����2��+r.PZ�}¹��-�k_E��H�<O׵����q�rg2I,S���NV����I��\�ki�kԒ��i��z?�u$_��i��&X��Z�=�)W�Z���g��0[���:��Ab  _tPďd'̣���}L�!��"t0���1�;V!�؋������5��TǛ��|��99c��L5����i�yn����v�S\�d��|E�l�$�\�)�^T}=��C�U���w�Y���W�4/{:��u?a!.�e�3nN���r�X��7l��K��q��Q��L;�^��/ ��
��83��%�*%$����� }��hAC��"�nۑ�,��g�6�G���ԁ�x4xa���F�?�g�xAh�]���k5%�%�J/�����cP�����Ry�ķ���l�W����b4�aEc}?��� ��P]��90U�^R�z��yu*�5�;R����}{M���Bg�R؆{!�m��{w� ���{��2�l�Jˈ~�S=^>�ח������b0���ADi�MvJD%i�T��'���Il�Zk���#Ъ)k����a��Ɠ_ �JD�����S�ͣ��r[����'t@�9L�-����������Y�����s*6��ϫ��-|F�h�.f��0��= �r`1J��z�zJ�x��x��\u�bTZ�V�>�(1ц��Cp�s���Ɂ�hA��f4Л��m�e8У8P��e����:Aȅ�<i���(^�!�K����r����$d���U�LT�e���a���~���µ���c�|�D��Mܢ�-n�+�$��_Ih�&q6z�'�6=0���HG��\ߔ�4����`�E�N���u]��7�o�y�_�椀x0Vde.�D1�X�Kw7���6`/i<��\[$\�뺰"&�(V�G�wEWP�m3�g�<����Ũ�K�}i��Ŋ`Ć���iN)?I^x��{$5�]{�I<�Zg!�t
x�ʉ��g~��N�'�8ֶ�W��"n��eA�wG�zŝ�Ȼ��ƫ_�������	1����.M~�)ޑ�q֓�ȭ(G�A�)�@>0�B�j2�1l�{L�~�a��"��(a���� ��C����G3�L^�x]^\c�|�=R_t����<��w����ZbG�LP:k.?J���J��RA��2��ĕZ
�;l�M�3�͘$�2����L�ilbr��ƴ�g����5�4�"e[[:{+�Ȣ�}��@�>cӢ
c�5 ��5���E1����QA��ul�nl(��tB������W��W�ǳc-������5�nfq��z{#j��Q��ЋdH�Z���Dr�kH?���3o-G��_�]�i��	�g��Tȵb�7X�+��Ld� a��a���D �6U��X�|�ϠbU����2�n�t�I`S���N�v�0����*0`������,�+�|DV%ǋ�ν�J�������&�-`���tKB�U8k�~�k�#��Z&+tx�/��U�*
���X��i��;��Sr<��e�+3�Y9KtKB<肟����j��ٕD�4j�[�%0���u&���<�QD���!�=V�\%j�{V4>�秛@�� ��<`�=Y ������TX�<α��mrSb��}L����ޢ[��� �bC�=Ic�jR�6�z��Wx�I����������+�z[bU4V�ݨX��W��F,�ݵ,7��RzG~:0G:��x)����#K��Ñ�������#�-����Z�#	��b��G�6�_�Ȧl�Ą�q�/Fz�1��t^�#���Ǒ�֯/�#{@'�e�Ǒ�����i�r�5~E�8�!d��2�fOΘқ���.�cD�_]ܝ�w,�S�&��I��X�~:3I䪣̅Q����Ⱦ4����ڰ�~��5��&�h�?ϩp�?	��7��O�W�Y~��B_�8CqpKT�1�Fh4��u� Y'�����ݱ8~�5z���?Jɋ�/O�����[���o�QB�MY���!"��4�s���e�tEl�+��"�Y��^���\���g��4xM��tM���_���k���X���a�۰��kR�^Y�_��&�gu�䪧�_�Y��t�:�5i��A��]�h��!ьz�D1�Cxcr�h��4�߻�&n��]��x��q�������_` �X��0)y6%��vR�5&Ky-X�O��S��o���qO]4bh�������zF�v>\A��/T�H���a�Z��bEi�G��0���Q7 �8�*99" ?G�a�;�/ ȝ�8�q�� ��r@^�2�x+��Č��M2��
2#�s�SjZ�7	p� ���L�|�E��Yo����9@^�0��~փ��*�V4`#�t�ʇ��QeC/P�@�7�@r������SOc0L�������{h�L��@�x�ɛ�R5���}��Y��g�k)�P��*I���o���hO�&�l��"��x��S�`��CIdϤԛCu�4���4�����6��G�a^m)�����0���16��60����	�~��k���zù����ߏ�~�{�߇}��Ϙ���E}4��=�F��W��MK�j����xM�Vl��JϠ���l����e��5�q��I���h
���~���1��}�6̳.}hDcT���v����ILd��tip�P1�<bR�Ud�?�h�?��3E�A��]�Y>�ｚ�ll�$�fU#�̾��+��[�����(��{�i1��|��L��ɻbs�R��8�ғ��L@��o���c���n���B���E^�Đz1�;�JnH0t�N�n����Po'�ki����7]���/ɝ���|�n�W�5O�w�������u�������i���q��Ѯ�[ y������Ġ�[����%r{Dd�\�	E�B$.��x��[��!c[`V��Wb��K�Y��o��g�>)�y5��K���ط[x{�9e���/n�>�c��I��8m �4�37˃��~�h�?z��Ɓ3��ں�oN�Y�&���+J��>a�����̪��j�b�C���<o?_��r��3��(�"aޝ���+(Z��x���\����Ś�#�|�����9g�g����?h�#��u��Ґ�?�5��G�,ԯW�eG) ��-Pc�G�O�u^♈_���p�?��_/wsT������7s������XA
���V����hI;��1�3e6�%�#ʰ��ї��+�c?�2���Iۅ� �|A<@�>�����4�ۿ�A>�}���;�ì"�|z&l�b����fk3����zt(#���8k_��C�4x79���h���������%,g0���+�O�f��{�X������|E���fj��0���FC���P/����v&�p��f1I{ކ�*��Ѓ=���\�^�O���M��F\ٹbNx�-�;�V�,�����?�XrOf��*j.ϟA���աm�� W�3�d�B�-ֹ���{?тᜀΞ3),�k�<�V`�Gcɽ���R��U��GE-�Ф)CIj�[� ~�ಢ٨�E'˷��`h���o�)��lZ_&��4&��~��d䯝L{K^�A����_x�#�q�S�Љ{�Dqw=�K%��A!���P�
-֍��/@�~0'ss�xL<��ZA�O�G��9���zM�?�|H�g�˘Xx��,n���h��k\b_�0�g�wf����X�A;�^y�x4`<�`��Pq#w��*��l�6h�^$�f����$\q#e��A��Qv�E]��/c}���T6as#����a?׷�`�O^t�����z�ֈ�Ф[(�]K-Nc��d��*��gx�OAl��K�~𣿡��dQ�n��z���Ǘ�q�؄[T��aXK�O%f��1�C3���J���5�M�)� ��0�#����#��m�(�wS%9�(+����$<m\�{�ۂL���f/��fj~`j�@��7�O���>�� �ɲv���}���5FѸ|�q��f& Z��Y����W.~��4�9� ;�Y�79�Ń<r��5� �Q2=�S��m� ��/�/���X(@K�Y#%�J��y�)�8����w,����}�QE�J��2�z
tA��R�y�J���@q��9��&;b��
�[���t!6QD�,��l�^���{%�NR"Y�I�ߍ�I$�[�e3����rߛ�O�Wב��q�oW�m��ܡ�ސ��D�!�K�zfZ����l�����K��;N��8~]�F �C@�)��|%�*�$�}�l��믋��^I&mn��,�dJn�( ��L�p��13� �P���(q�\wm��O�οȑ�_D��OC�%�9�c��}&	��>�%d��|sQ;0Y9�|�z��!��y����y�csLN�����"���YL��.����-?ʭNwN�ix���ph;T˩�Ê���m�' �F	�z 9̨�K��+xz��bd���Rot=7�֋�3�4�v�tz��l>��2Z���C�Og�檏�}��2~N��}�R�L��g�%�����1{���Ty��E��&���f56�D�@~�[r�T-����ǈ��-	��[�=h�֬ǭKT�qw���ꁯ���1��X:�ꁫ���x����s��FY�{���Y�o���^�z��?���1����êƶ��_Z�o����l�\k�7vc�޿����\��O?�A�}~�!�{�|������\�@$��r-�ɸ
�����	�;��E�Jy���w������Fx�����J)�P�O\�:��v$F���a0�5?�����itz��S���È����<��Cc"�+�'�&�������#�;uy%G�7���C\UHbɈ0���(�.����c�Q��F�B�4��Y~�+ܣ��W)���p�k1���g��hԗ����	��aJ�{)�~{H%0B�Z���~���?��ܐE�+���IN�|�D�C}��>k�C!߂	/S��� 8��^v����<������q)�ݴ�4\J�H��=*�e�W�E�\
���=?>�V�p���"�����!s��L��2�ɃzR"�@7v!�9H��\"���4���[�~Cr��Jl�i�-�ú�/d���f �A�p�Y3�<B17M�N�n��i��G �6́II���B1f�ӻ���ӗ��n������]O>'�(A\�m����1˭b}�u2P�6��7��w���Y3�{ �jc�����d �M�W'l\���0>���O�㆓GS9�H���xD�7����-tf����SQh';�;��X�E;iS�;�$wNU�%l���x?KĲ��k�-+��TĲ8���|��/8f����B����A4N�Qy�h�Ya������\�T�D��YiX��.���a�;��/�
��!'��%�NT[oӴ ���8��e�Q�R��ix�Ֆ�j-њI*Rh�-Cc����WA���J�: `K9{�'�С ?h8�X^q/�����uU�o�^/�V�~�k.������\�*c�[�W�u�a����Q�����覸E�Z������X4ݐR:�ÜP�շ�{�00�PC|�-�*A���#l�Qģ3,��	�PNyV%�4D<�����h��a��#J�M��uTCT�@�9���$�N}.���|��Q���:������C� ��N��ZXܗ��G�%_oœL9z����d�\WG+X������~)M$����%��pF���Y"�{��-�X����dhYx�ݤ$�͹��NQ��fv��x9�ͬ�^=E���{�+�	\L<2��щ3땡#�|��
�g�u��?U�|\}#y� ӳ@r��X=�%fv�ƹ)����,�idq�)ڛ�.�l"��$�g�K�=~N9gV�?��'���})�/3��r�2����c}����O3�~+�-g� zg��f������K��l��iVp��k c�����v�f2���뮡����d��E��X����a6��j���v��x�դϹ�2�Lt�V%�8�F�#G})Z�k�hc��+W�}YL`G��6�&����!�����iFCUp*��k�������9��A|��&7�kp`EF��'��F����
�\l��'��`4�����rjYxW^?�'�{|M�ؓ����7��ꤤ�����qmo"u��7��Lr��F�q�c�f�`
����B�s���b�r��SL���G���T5�L�G����f2]��Q�����dXJS	,�����!��9�IWC��돱S��H1ߧ`e7�Xf���LËO�}���!�i#�F�ȧ� !���ګ�qga$�@�?	-ة�*������o�HbU�>��iB�B���v W�p��w\lT�7J�\kSO`����F��1̣kh�i��;o>��{�ˍ�@I:CT�Fl���្�Q�w��`��~�V;*�U���1b�3 �����d�[���Ct}o�X���y���Gjߡ���țƨ�D1IX�
�!�>o<�&P��YQڶg7��F�}/=�>�O���Ǩs{t�O�^HwJ�CX�%���9�\&>{ǈr�v_�S�3�?Q��8S	�� 2e�׸���|m�r�$i9unڮ}�Q����y�Ų�ĝ�4��X�L��i8|��>�ئzIR�s�BQ����먗�XŪc5��>�7��L��mσ�Ô���6�C���Y�"��{��6� �P��1wɂ�}�T�GjiQ�pQ-U�j��!�I���wy$��d}�|=���8�'�-���G����[���������5�YX�@�5f���F>�J(h��v`��-m��Hۣ�2i����Zݘ����P�G��i�!M��!/Q'����~�	3ObNv7�
�<�'9����5����g�\,`��:��U�e|/�x_ǧ�OST.�e�/��n��4��z�M�I���}�S�(H�����o��q>�dr޼��l�QP�
��F�1�}��$(��<F��k�ե�c���pԜ��
D���4� &��
��~L48{� |@��~�{�x�/��k��B�T0��\����f����`Ok�����`�`���U���o �V�Ƣ�b�-�<��S�(��J�J
�w��;�<w_��n�th�p�vG�#�Ұ�(O���^�����*Tf��1�N����������u3��Ƽ��-Л��5Ȇ��F�΅/w+��p]�֯h���&x��[��7��Q�a����3��a8)�ӳ`��rʣH��t .PsA���:���瘸о*s����լF.Y�Hp���b�1��S��h�_j�/ �O�qD)��r��M��W��j��B�u�x��$ G%5������m�Q���/�:��K�bu��.��"�cL�F�[��I��?�2�Z�ɵF�a�p��t���Be�l���h�tݨ���xR�T`��o��L�Qp?�Y-3b��*���[�����Ɨ�-V�[�@?U�^o�K=�>���Ys��\	@����J�<�O^fJ�����ЇC��N.���5����@&�:y�s��7�d �{[Ը��fŚ���o�j�?Wӈדu��24cL�i����j�qx�Y��S��\�G=��`G:HAAJ|�(�L\��M���T�X������ �`w��.�۸�b9	D�7�I8=�Y��y]\��VAZ�pqZ$�RtR����F��ӝg3D+$Ї<Q�؍T"�]�Do'�F�h���diH��kx�H�$���j�\َ��c�p�e�YP��Xok����"=4ѧhe�� N�\>�p4M�\>K�ZT��FQ��5��Q�ड़�F���l#��1���6�mڲ��V�*�@�"�!xD�����<��XF.f��G��b���Y�@����`��#8�9�����)����ߢ���7�U���ux%"��f�+���T�v,�6wsy��|jԂb<A⌒aT�f��c01���ٽ����x���u+ۚh��J���1���a=���t�PCJ�A�s���eZ&5Ԋ�y�\w�._�[�`���_��7|N�D��Z�F�`8�Q�+���hšb�����F
��\�5(Y�܆�d�bV+�e��-��ժԒy�N��h#�{����uޣ�ۧh`<S�q��Ry4��7�S���U*�h��<J��6�(�F��X5�ԧ��0~�LO��ir�����{7�پ9����_
ީ
��C���)�}!�ԙ�Et�i�|!�'��ӆnt_Q�E�b�L��&��[(/�[܍YtB��0�ҭ�!���ծt^)�)!gr%$����`l��F��v�������&�*�L�L������2�l���C�{��/������sL|E$y�P���]�@�o�|��,�^� �K���)P@�dNe>]A/�*��Fo�5�s����Ϟx�i�
h����4z���	�[�獘X�1	><�P *k�������h�_|��8//�2B���8@�&�$���<v�����y ���ٓ��{2d(���x�O���8;1�@;�_���H��E�ǨnL��Ց���!�v��?�j��EX�� �����"
+���^l���"ҡF�H���u�jc�t�ڍek��Ka����EÍ��n�E�f=��ژ@|�������_0�~'>�\��ְ���P���E��V�{%�����'�1n�|�I!7��q����ª!����N,��Ff��u1�W{A�������CV��P2)_��K�������Go�C|[X��,� S�	���s��j'�O�S3�������#�k`"��w6�Y��\+EqIw�HhSJn��Aek)�N�l�Bl���\A���e[+2�.����ǗP'{��M�8�}� �����>~.&�L����;��t�w-���x���e���^6����L`��O	�S��<��e����O/ї7�����5����&���~�#0��D��
,���tX��(+�?�r�� �B1�/Ε(f�y�[��^�����\�=��qG�����C�c|�e?�~�S�2)�&�m%�v�F	˱�c�r��T,���;�<��>s}	,g%f�ặ���Z���T9@�x�7zK��o�ݬK����={^<����dJ� ��/Ə�/�'�h�I��Ft�x�$��M&�+�ޤ�G�{�e�������6d;.�#݆�s���?��=��?t���C� K� K�������b����Ì؇iF�!%x�(-�[��>�"��bz��=��}(�ʱ��[�4)��>DܱU����I���}��>bMQ	/%?�.`�����y������Jɿ	G|��9V�jo;�!&/��7h1��c|�>��$D��5	:� ���^��Wm _)Y��E��m�IYu#�H-��+��L����!I.�\{ڞ$�qun�����Yi헫��K��a�����?�T����a�S�>��Д�FD��*ў�G��
N��Ϳ�8iː^�Azu;vk�F�Ժ� H�dPV�CL�R�T���oz(�ף<�t�����?U�{GM��6��o=�;囨�������i�����V?�FS^k�6�0��q!�U��2�W�q����o5�-?�*��k߶��!Z���c|_%��c�ͳ7ӹ�������*ҹ�+�O�ǉ��B�¬A���<{1'�*�&��Zh�!Ա�5�h�|�^E^Cd�z~�:stW�7�C�ڳ�O�B���K�<��=V_���C
j�T4��/�6]���,�o�uB�ֱo��S#�o�r��}B����ufd���y�Kt�J�ӜX�Y��G"�W�j^W%r��A��
n�Ա����nh��C��[5 �
Թ�Ƴ�*��>xD�zP���>�*�~�P�@�K#Y�������i|�-�}'R'
m;��[:�Z�w�鯳�˱T����{ܗI0�*;1���w� �jL,�`G�e�ƭ�0^�����$���-����K`,�F�k�,��C�^�X��2�?*�W�Lf�@��I�9��􌱨��,�%m��.̂�BwE�Q2��|F����F�25��w�"�f7)��CI{��5)��-��ߗ'C�g3��}�< C��b;��֭�2+gg�N��R��md��O5�0��(� C-=���#�?�	�&��b����*��eTQ�� bx�Q���T���ޤ��k�UbpfO=�9"~�;!��no#�<���3�x�D�5��KI <�4�?��9ɪ���O���z���������ŉ���xo�$ �~J�f=��Ap���yER��N��28���	v������Ǻ�C)o��M�}� s����b6�S��<ǉ�u�W�M3��w�T�'�'704ja��Z�GK�EK����h��v�[};�?��~�ޏ��:D�ǟ\����I�N��>58��h���DQ��w)9dLVs�	#�����YLQY�����	��&��_�~r� ����p�W �
�_�+Y���E����T�K�b�)9�f����Z��ư�0�r::�Y���؈�P��?�������Q|阐�'������m���'�$��
_��f���~;L;�H�r��b\�>�@�p�R1*/��3lsbXٵ���0S7��=��o[��������on�#��6�BGW��)`R"?��=#�{%�o��-���9P6��88 ?�7�(w�p����ް��h��'�2��CgX|�-�bI����ֆ����w�R򨽺�0����x5���Y��4�j ���Cj�<�6��L�oQpM�u�N�ZC�.tJ�m��8Ͼ��vc(�W����b��r@1~�P��˷3'g�T/�C����p�o��j_����iLE�D�¨X2�B��{�}���ϋ�V{n�ihw=軽�i��?9ɩʧ,#�ɣ���Z�z��UQ�|+Fo����!8��&J,�cͲS`���$�̓�1�Ԓ�H���L�3��<.˹��{����%�u��F�����_�yʩ0E,��r�����A��wk�'�ߝ�}f�IyvwX9m�$�=m���
�\[���8�ϱN�S<k_k���<��zs�Ӝ����o��'���w��z,��e�q]�f�I��}��`r(�Q��=�vk��᳎�څK��F�a�}���_G��BU�Z���Ol�ໃ� �UìNX>�����b4�☰�JL��d���4?������s.��#�!�
�[v:Y�Y��<]҇NqS�}�wͻH��O��ȏ��������
�Ҡ$11��*�^1��	 ݅��)��Q�{���
7�Iߙ�I70�] �q6���#�E��!��$�Ʉ���6�|�0�~��͡Ov �P{;{�2��ڈ)�0?�n}��*���w��a5F}�KԽc���r?7�גcy	qۮt[�	�
	´$����@���?���X�;a#O�a	5��8��gc���*]��4��.=7����k�d,��:ͣJ?����ٗo&�8;&�Q���5p�!���p/8JIȷ�H�S�l��x���N�ׄw�.�,-�nq����Sw`f���`-4��MNe�.Z�%N�	���RC�<R����fc�%%/�1��G<�W�����+��eJ{AB�D�RE	`�h����2)��n��M���|�mDbfUC��b����o���[<�H�m�+ȯG�3��ʙ̣صӜ���g���a��}Yd� �g��mx`<�q,ԟ�0��3<�	��tqr'L��7�D�-��F��^ ,��5^��N�!~�lǢ`�[q�-�;M1A�mM�������@��.�����h���H��J��P�J�����*_/߅�?��(�y��U_�V��˴�ϲ*��3�䘞Q��=ƨD�,5����1���2���0�s�äo�����%�;����xq7R���z�;jDYRR|CQ;Ei.Jw=5t��eԫHˌ����Jä�����TW`��X.
+��t��%q��[�
��@7 �L�ZXA����T����������0���Ɇ������H���'���1� �s� ��]Ǖ�x���7�`�&u9
�(q�R��(
����D����B�1�"�R^�%Ѧ�umQ�.�&:��G�Qa�Lağf�{�P�Rn�|W�^LΊa��������΋aDЈ���pX�K�,�Q���i��q%e"�8�4`s��d�$E�)�}���2WR��#�x�slNv����_� `��Zt�mJ�����P�н�i?\����Mǔ�6�E�ޠz�`�2:�<�>q��^�1���UCp9!���%�R�� ��hH�2��<qNe>��O�Q�����S�N_���# x=�*��ǷhB�ߊ7��ՔpGoPS$c ��ѽq9^�1�{7����Y*V���RM�{��e�ؼ�N��Ǭ�y��c�Y��R�KF�J�|(:�$��ݏ��S�O����UYw��o�Ѽ��C&%� E�9\����b���nJ�����`{7��9�M9=^������A"�c��5]�F�c;�Xe���<g�u�9]�8(X?�Qh�>����Lwʼ!���S� �+#�#�D~?�0-���ؘb�Z�\}P%(�r"��R�'�d����ڧ,�	��g��;DāQ�o�#�v���d�\i/M�W�-�#�80��x����K�ؤ� �и3��؀CG�Q���h1&zKJ~�@��u5;&?[$6E��T��� ���z%��3��J�+���C� �'�3sgw+U
�2���P�[���x��1��x���"52o����a��9��1~�E8�z5T���]�V�#�FN�D�Q�T�L 0M��?��Y[;�h'w����I�`%C^���5�J^]��x��������<�m�Ǟ36ڼm�l��s���$)�n��𺟋�n��;�v,]N�XfL�X��9�tr��;>�<�V�@~��ҷ�ܕ2���+�?���^���S8��NiX�P�G�-/��/��R:������k���4���QϩThĵ�LA��~�l@ʷK���%QO�G�
����rB�OV��Nn?
U���.�^#=��%,�-*n��,�}-��Ȑ^-(���B6�}K��,_���;�c�r�S,�;݁[5T�(A���9ţ���K�Aӝ�4���$��BJ����*��g`r3�h�챬c@����|���+��n���2�k����FC�Ҳ�70֢�)�I�
y�ڒ�"���K��~�"�yL�9�,�fjKb��!,���K�Y{^b����p=*�[ɞ/)B�D �0 D�:�ܪC2��.^�<�?A2t��W7�ʤ��D�	Tëi���q��em�~�*d�9�-k���i�_�:m�US㶼�j�-J�E-q{T��.Օ�F_u��ȣ^�Ŷ�~�hBO�l.�@	йF̰�C�O�_iNd�i!�9�0	��Q�g_w�s"�^��~r2�@��pZ-s���|�������d�>ŋ��vIwY�g�HZ	V��݂0�?5���Y����yj>�{�q��6�|V%q~c� �ݱ�i1���]�vt��`�Q`Ձe4��ü���\�8ސ�s��ǯ�!������t��R!���B؂!
n)ו��׵@�����m%����d~�t�m���mI᪷�_����3OR��݂4 &�#�^�<c�{�@boz�����A�
����9���5A35��<�%,�ò}�u���/Y����L��flX7���䅹s؇F=�����\?V���,�
�WA�v^�]#1?2��G6�=� l��h.'�׈V�"�D�e�ͤ3���o��L����\�Lbδ/F1;�B:�X
������S
-�<���:����&������y��d���wֿZD�^��X��崂6Ni�ej�>	�u~:�(D�? >A-9D�fq�����B�k�B��꫆"C�(7��*�,�b&ޅ5B
��J�`v�	]Mf]M�]u�t�W�)}�4ll{:���t~pJQ��VO$�����%��4/� �Ԫ<�g��,P�C_�+p>9pÍ�e���nq��PAƊ ��c�D��������<	���n�/H�yC8��@91S�G�ŋ�2��0�x�]�[8{^�:���\���W�u4L��u\�]��'�����k�(�d�MZc��QIQ��&W��yc�>�s�� Z@�l�(L�2�Q�7��i]T�W�I��>��%��"��5>@�r��*^���]@Ѿ��r���܀��<���#�l���<�������o�9^������(sH�Gyn֗o�hD��>rJ��MU��ͧ5M�o�W�{XgX�� �oU���� �X����Ū��vO9�Q4X�oVGBs�'Q�XI1���4�ϲѧ�蓹������㶀���d����b�?k��7���fUvU9�W����F��!�O���S�Un�FB�u��Mb{�����9�����_m?q�f�`?�$@E��s�����A�N`)�34��g�2
����U^e I��狼�L�`k��x���_��x55T��c�sh4;�p���0;ǜly^�<�O�l_ D*S�uV��qªV�XK2Z���c�<��F���F���,:�;2�`����#��y�Ѡ%p;8�%pˢ���A��;{��ȍ��� ��,j��x�#PGA��<����0T�N�G�&�a��Mx�T�ߗW�υ�(�C�Y{��*J��Lj��Iz5��㸥a%x��F� �/IXz�֡G�JD�j�6��f%�w���Sl�}�XW��w��kZ����s���$����ޔ���e�k&��h�,t EZ*�=�M^,؀U����KhXt67:��l��?a*|�W �8f6��o����n?BE�U���W]�u���@1��,����Jh��9���)r�s���vHC��>D����QEai"8��7��ns�Z��$oGVT����	��W����E�Ű7��О(��#!�A �����6t��V�c��K����}�=�m�@~�^�D�mW~�'[n)�m�%�R�Hl�ch��V^���� Nn��h�Y�<��z#o�
�q�u����?��w�i.���
����PtE���M�bAϳ8x���=_QBfʭ�3.��8�t����%����o��8��F�~��2P�F��p���т��[�bZꍆ�������"t;PQ��Y`6Kv��&�֙����)�w��ƈ�R>Y��.�=��K��Ø�~i 2u�v(G���)�]��Flu=����J��H���cY��^� ��K�x3��\+�K��8vsvS����	��"��W��	�n��H�s�>J(��-ZhȂd��P�o{E���y��D��G�M |d������&d�g�݈��j�h���k�g��\�9|"ΡoX�`b�q��s�P�./+�%O쐎<h�.�BۜJk�p����Mh�l�CY����IuL5�7ӣ<S�s*���¢1Y��L��[����޳x�n8��oE[��)�9�^�����{v��g���N*�d�_I)@mqe��,� "�fyn"	Y�cy�`/�D�Bf&�2�z$�$�]�x"���t�lb�&�f�� �_7g6�,"ʰ�q �LO�v��P7̝4��s��-�k�9s7"EO��(�G�L�
��w��|� �����r��nB�*��-�у�].���c�=�IZ��I�n��/�u���쩮�bcXw��uӚ�z���zi���ڊ�+�Ba�SP
�r��v�2�.q�#'�d�x
T����Wj�#ݮꕜT*���y�>G� ��@�+��@1��Pq�\�%�m���ɩl���>�nS�B)�R�&�rG�ː��	D`�-ڔ�Dg=�x�q������A����"�g���/����?�a�O��,��腘�N��f�ro$R�+t��W���F�3͉w��t��FD��7M~��gT<3��Ӽ̓��"��m����K��X��ߖ�`1`�u��	�Z��B?�xTX>��� �B�9G���3��Γ�qw��*�{���I��^�8GYl�D���� &~@WmA�`�;�h�:8���~Fr�f���XI���=�ٟ��@)f�Fv_6�c�{���'�c��sp,��Uo���;s�((g3�3X�L~�T�����pZ��xZ����Θ/%��&�z�+Kw&'�r�ތ����@��dty��@��@eq���m���4�@el �� �;*�?+t�չ:Ņ,V��⒲W��P�D"��_��M≷i}q7���H�3	�IB-����t@��^���50���f��#���MH��ڎ��g�O4��e1LĎ �� �y[�_��Qc�yz���NCT(�N����oy+>�q>a�	=#M���#>L'�#�(�a�*�8�w�q�Ŕ�r�w���ŕ� �׽�at��jcиڕ���.��IGc�M5���A��pqA:��*���)�HbJ�2�I�������l���
un�r,�53��o�PUc�4�u����Nzs������0F��;15�eh<�����R;p+x�M�>o5�)��d&H ���d�b�`������ަ��Ç��)��W~�n��-��2Kp-]�蝻�b�bdк
b�����)��GP��)��w8f�Le�s�D%����N4=͐k�6Y���K�͢lb�x,�K�Mt�Z���1h��E�Iȯ'���djlNv;_#���"�N�oV�L�{�#��WB��P��o���7�"}���	5��~�PRz�ɬ$b�y`+iG(+�CT?Xd�Y�~9f�Ǎ���N7U�?̳����]�e(�W�3*���?�2bY?U{j�hl���kO�6��+�f���Q�.y %q�J��6O� ���K��(~,�n�r��嚊�]#�It�h�,��q3�;���[��:y^���Lޢ��8�FX	���%��cu0.��rk}��ڦ��*�ᝬ��,i�(��4%,t�L�(vʘ�����^��^��4Y蹡���`Nx���Vݎ��E�"<�� �l��N�k�����z	�f!�uU��|Pdr�РsK�!=H�4�\N`���k
��&�R2�^������t�܎���b�9��m�k�C��2���!J
ȓ!b^@�� {j3x�S��YG�zk�F�6�׬�дV0
`�C�W�<G���E�tT�3�N2v+0-��♍�S�� �@���v���T���Gu�1W�x�o4�%��=�6���rOg�?��f�L�NiRo��D�GL�{��O�mA����d�t�ī�v�o}�
'��g+�
��(֯�J`�zø_=F�ny̨/,%��3_�a�/�w�w�	��އY�X�L�1��ơ2��c��]���P��̳9?�˗� %u�J�A���ԇ��C��TV�u@¡�;oo՛C���} �߲�Z�F�X#�|�}a�AJ���V���� M��<h���4x�AVlKd�g#�T69��g!Z�<0t�)&��q\!��QH��v3� ��B��f\�# ʩ�b��.BX�f�� �qbr7<O�M�E^=�_�)����ZM��W��vӣB�;��/�	�S/?ǳj$?�z����0gh��}�ڽ_��)�������37ol�2��#Q��l<pB�߾�0��xsq}�?�-�?'�NV1�[D�.0<�A!��w�8�½��И}�����R�Ǧ��}9����χyQZ9Yu��MfB{���S�b�۳S�m��.G��Vy�D�j�4�s���A^�V����*�dk��ۖ��2���H�.�%ubKʀ��7]��ܹ$5�坮 ���́.7L�.��o�v�L��������%�~�p�*��%��^!g��{���r%�FL�]~��+�%����T^�a=E�	��r�r2Ϣ�"H�;W�곲�6���*v���J��;s�Kx�m�<q�S�k&��q	��Ѝv�m��+>~�kiط'2�-�u#ۨ���{��,���h̓�,'1��E<�#\-2��nC?��[�y~��|��d3��_�w��ґ�31���XǏ��H�]���2����Q����'�4��X����a��c����~��4��!LV��H`CLh�
b��DR�N��[�1��L:[�X~��YBd�徾0�1l"���p/�	��Ӂ��qB�Y�d����{��l���\{��,�;�1��d�����!^�xy��}��:ADu ��9tGE�����cԳB-%~�"�Ě.ܩ��.�5��(���ư�,�,I>����Q&�J$��$OG�[��{�����4�Hj>&��[��(}�>_c��:�ǺW�i��I�'&q��L�6��$�?�6c<����~�-͌�5������.��I���p��pK56K��G&����K�;>��t6ŀ[�H���uyͤx�)�vjy�fx6�7������ĸ�����ى��ڡ��~�ۄ��Q85�l�f�K��bkP0�TE5�G>�1��/Q��B�0���T0"�Cw��}{�Ѱ��w�N�&ՙ���s�ß�cy�MFz�zJ�^��K�{6ʔ �⶟3����c]ٷ��퍘��0`�n(3M�Z9E��j-Mu�t4���/��kT(0|6�h�.]QVDZVsy�F��+�p�W2>��Y�~~"59���o�Y�4����r8͢ê}Mװ��B�0�iwfP�PS6z�:����^��_�F�F�\3��$�Mi76��	sPi�'���pp�/�4��r����N~�o>J���(�$G�՚�?��+��Iɑm����2�N��)��b'��W�ȫ���3�N��N�z8�����<+ؿ֝�=<6p})J�����ߏ�I�~L��2P��@ɓ�&��mע�[����-�)
9+ [������Z�����*�ش��+�6�t��Z�$�+���h~2 $C�����r�챁����NX@�����^3��i#�nC��G�z�H����O����M�r3mb/+�gJ%��
?�����$�R�S�$�O�pad���Y:��K�
��>��6'07*8��o��u�m��饈f�pX�c1���\:��c{�Ÿ�Çȩ 2)/Hn^-Ű ��}���`�8�5,>�� &�@�J�w����a�n�](L�2W�0F0� 1���d8�μ�d^�&���I�W���<���yO�@Yb�(�(P�h�,�l �H��e�*P��TH�(��.wDQ�XT(�@A��"e��zc@����9��$m��}�����ܜ3sιsf�̙%�������oА�!�V
�XI���I� &)��J8_��ws݁���*�	:�!OJ�q����n08���/�(��;0Y5������Ó��dC�� ķ�U"��(�������=̓�+�T�1B4�I:{�����Å���W�C�x��ZJ�.�i�|I;Z�y�{f�,��5,��k��Q�?��e�9��*J;���T�^�`L�� ��@����蜇��V����VM����bpD�d�_#�;N��p\�����a��P�X��&�?1m"���1��T��E�q&��?�s�
��f�r&+2������-a2N��:�o؊���Q����t��	����9��8X
�����̊������s;�����9!��2&��ɐw8���kAs���c�]>6�[���'��	;�I;�����/�6�j�^ h(�����}��y��.)C���x����g�X�\>�u�$�b�l<h��]���r���>�螁}�����}��_7�����U�bXa`�𳤚z��b7�	Y�
�7��x�T5���9��9�ݮ6p>E���AH97n��\V�����y7�N����'^�-�rg�1�F݋�2�On�=4P'o�<���k��@�y����x��&k�Xc� Tf���(��+ZX���"��7�I�&����N�MT��pk�.�K[c�qp)L�j�q��8[f�*�:$޴M�����wt2�ǒ�Y���gAzWt#5� (���%t�z��Z| [��rm���D��o�$���R�mJCQ-QV8{��/��0Y����̎S��>�A����Ƃbƹ���8��?�E]��3G��0z����@ť�G^����YF{<@�]�s�yP�RvD�6\�uB~XY�-m�l8�c�=n�|�!c��>'�y��y�x�����W��W�2n��n3wn'[��ɬ{���&�-���A�J�?q�t����tV)Ǩ�FF�.���W�����e$u=�kX�Ǳ�S���P>�g݈M��s��0��S?�n��_&jh{�z�OX���3�������^�V���pm	7{ϊD�YN��~��n�o�k�+"����g'�+Y0I�EK6��f��)6%��򪎯ڍ��dZ���v�% ����}����ݨ���zc��pw����X��!�&7s�ms�5��꽅�d2,�Hw��O��NcA</��Xp��n��&0�g�7)'ʁv�>׍�/ӳK(7�]pPM�tubHg`�Xg��´ה��|z<�g�TS
�ӈ?H9�������5Hr(���r���� :�'���2�oeq[)�q�`�#�ee��&�B�n�����z��q7�x*C�)�6�A��94�x��}�}{������0�k��>{IW�s��!���J��^0���@�6&��MJ�?H�,�-Ԭ�#�Kh�ha�T�^�
oOm�;X	{j��had��1s�c)�e�yH��%v�Qgz��$����bD~�����@�-���I��Q��X��D�#brw&����{���T�`$#�\����J���H���oy�N���	ؗ�X�I��QB��c�:plv�EKPh�D��"p�-�˥�"-�&{W����F.����U-���W���k_���̔AI���A��O���^Nu6;L��[�X�7򪣰�3����d��+���0�J�7�e�CNP2WC:4��AXN�����f}�B̳-����'�~�I��G<6��j�v�4�8����L`��2�`���m&�?� k��N��v@c�q�!�������l4n]2�c��'�,̒w��t�3~=�����<�UuS���_��5��,7nD���{��L��3�1 ʺ#���Ocf�ѽ�
�Hȅf�	�������}Dq�ˤ�~P6�=&��D���@y��;
w���"M=9����?�jP�o���]P�F��T��"f&^��L��xׄ��&���yZ<(`���&�՘����4R���u<�������m8�[Db�0~�g���{��{iN���]�렇�)gJ���ܷ���[�r?��}����'Sx~�ԗ�]���-�R]J�H�����/ɳe��R0�[�h��=���G��Q��([<��e�GYڣL�(S{$�G���t�(=(/�����Լ�-_fG��svT�.Q��@��p�P�c�w@2�՟�QH�#�Ǽ�X�1Bh����+`�Asa	·$���b]��0P�ԣ��W͞CP��ҋ߬	��@�'@��@5EPM�/��J*~�&��c�c8��c�}�2n�Z �Y��&�u�����Z��­DP����߮	*��#@�k�z����.P��E��`P&��f=����-BP�u����CA��|_�ڙ�A}���)�&�V (��N^�P8"������8s��d��?������ūC�cEƾ����\�Nֿe���̹�7e���*��:�܄8vF���)�1x��M�e(>�'�C���{���W�kG��a\[�ץ����2��G�S�pLP�A���r�{�"�,`�N��x}��.,�E��S��2�5X}.�����p�;�@b�^��O�3�Ö�¾�������	v�K��g��}qd8؏qEV���`����ixvx�χ��n�[1�5�	}�v�����f��8��!������F����"-)�=���!,�����熅�;�N�]���!����fJ�\T�(L"�r��]C�\�iÂ�>��a,� EʙlM*5��?<$>\�0�̉��|z��Q����6͂�9���gǿ�4�&L�6�}��zy�Ml3��C��=�	=}��|:l8��w�.��B�7cxI�ݑ�iG�5�cm^`i���ٹO���y�!rS1�0��ܪ9�l�O䊏���Υ����G���\)�	��9�)��9�zD���LG�i�{@Ҿ���gj8�I��Q
��p8a1�ׇr��k:��!z2��Q.�aM�%���s� ��4`8���� -8�pb!
.�����f83���8��Ty���e���YŬ�w��k��T%��n���5�)�p����pNډ�L�s1�z&����3q�p�� �������p8���_�%���p6a�:��4��`M��X��y��}�B8��6��1ۊ����]��!狚B�!"j�����b����"~�X�<	?���gglM����� ���� �/��DW|�V�[�N6�)WBc�~�e�@:��ې/=��r)2���}����2���z	q4-��+��v���m���}��͠�o��BWK5�" wG]���uhx�qP�*|�!�p�;$O'ɛ'y�x̶��5sK��*�*���C�_2�xp.�_3����~E������٢T��)2�}���I���US#����
�2�}BaF���z��6��: +��}�A�v��N�ەG��!���*����iTcfț}y�O"�M��?ۑF��^�ɲ���l������jz�������}d3NWM���1��F�G/��#0�K�SUd��{�ئ�1�f�47�ю��M���S_q���I�~zv,��գ1{L
W���������܊x�{����h<S���Ad9=H�<Զik����ѯXD���0�����Vyl�1<{��YR���S���:)�%R�^G�ތ�R������INZs�!'ml���eO]�w@ߣ�~�g�6w�O�����_�,��1�����L�ʪT�U�\��cnp߰��J*��l��������b�A~��06�a|6�#8��(�#<A85�{��گ��j���!�����N��m�D�ȹ�)1��/��4gB���xE�3ĩ��1��y� �{Qj�3��H;s�wD��O���T�>��;�(rm/UM�z��@��w�������͸��_�"G%��Բ�OQx��?
Y)�Ld�`o]�ǫ��S����Ş5!��iv��${�w��~��w��U<�7�����d�j�2��,�I7����oK�[�����ժ��Պ�]B�gXiaH7�ĢSdv{�w�&�ߖӗx�t���vC����]{�sȻ�X#����)ǔ����X�eTe�wٽn���Ր���i���_����uU��b�S䠰+�~�&�^7W� �k�����d��h��J#���J)]ݜ��b$הgz�݅ה��ܠz�w?CV8̫������K�2_��d
e���3̖�7�R��J־������wf,-:z�W���)(-����H�vN��U/X��y�R��'K��������$.]=M�6�_�.c��t�KI�\
empn!rcݭ���C�V�,�R�Iϱq��6A�[\�OG��(Sd~�yQ(��Fm�������'U$��Y�Yn��T����TwF>�W� ���٩o�uUD��{��Y�u��Y�}����ށ1��{���(�dG�|�"`��8[�X�ڢ�ͅ�W45��[��i�����������!)�8��}£b�1�bx�Qž��
}�br��I	��<[�!L���H�g��d�pZY��s,��Ѝio�'֮�����|����ГT��K@ o1��DU�Xihk�|h�kz��A��saD3�y.��b=H���21��}"jh�_Hj��R�/'d�_�qJVRfR�@���3��x����i��@�zAf�%�����^{�Qɻ��Բz�u�������d�[�����I��~b��΀�؄�<o����ҸLL�v
�i��U�H��z���F��0X���%�_�C��K�mQA]u�Ќ�cъ:z��Id�e�5�ݮG$s���c��%��i��np�c���=�=#ܺ�҂��V��9ڏ��@��g�RK�7�UN��U:���ag"}���HP%�QјXt�ق��	a���A|.?�?;�B=3�r*5��:���������,�0�Z��ߝ���^�!
R��O�m�o.�����Ch�����7�>�]��ԭ�]D���B:i6�әf�Mx��� �1n6�aMe{����q��ދ�V�)�ֶ�o��V:�������A��]u�sm5��F�%貕%D��dV����\�ˀ~�=3I���v�VN�\���o��zMK��Oz�%h��SU�r�@�!/e��\�(�t��:��r7�\������D�<�՜����ؿ��F���Ϙ(V��3f��S:�U��,
||�},WM���T���Qa'n�D��l��j�d.o�O�wj�T2�t�}�8��d��71�9�6��;'�HȵC�q9'��{�������O�>n��G5����<] s�V��-�}����]��h��ǁ䏷/��bŵ��RUSXk@v�2?��^'�8 a���ѕmH%e�
=trD`Sg|�����gF�>����>gT�t�S��U���^dekՋ�B\\p}>�4�i{��m~�丛��f�����jO2Xd!�}�Vy�2b/���ǌ1y��3
�9G��V��.g�����AV>�{9�� ��׸�����]4��7��}���CW��>�Q)�")��T��Ī0F�[�̄�),����&VQ� �����Ѳ�2y�rF������Xԡq�
�ͩ,�Ҵ�>~;���-X�N8Y�q2W�h���|�`�T�a�����G�����n�X�.a;m�G�������Buv��Yk��a��G� X��;j�F �YSٰ����_�?�C�T������!�Ή#�U���/���ˣ8�2���aw��������Z��d��� �2����Bf��w�h���">�z`=��-\!;!jF�0�';�9�v`����
"�X�ԉz���c.I��t*���Ԑ�~q9�&p�w��	�܄���b��������?ھ���I0�w�Wi��q�@�k ��t��*���L��r�/a
���Kr�C�y��B�������~Bg^7S������Tz��O�
����Բ_��W9�U:�AzיL�z��<���l��%�N�����t����EP���q��Lj牝��ک�\	Nrר�>4��
ʠE���1�L��y������x��}�{��r`�NIBԂ��>��O��b��CE��������6�/����<����@S���ʀ>sx�j'_̗�t�wDoMHϐRő�T��c=�ӕsNT�Cs�L��J:5!��su����d�ҳ��Vw�!���Ӎ��h�pkԯ�p�l��ͷd`UM-��
n[]ն�m�3ڗ��iy[l����95Z��:0��
H]���?�eS'Q��P���D��j���� �W6�ĥB;�XVA;�(���	TѦ�4Mk[œ��P�vȓB�t�pky��z�?�e��{D��ϺU����oמ��O������^��+m�������D������/n��W3�+�����D�������z��{�v��ە�N�p�3����#���^Gɸ�^�1���}G�TI@�Ǘ�{�=�g�Ƿ^�{�v���T�=^t��{<��Ƃw��6��T&Ӌ���m,IV���nű�K�xIJ`H%qp?��-�k��,�)��gxl��_� ]p1��7���x�J��,�%(U�͆J�u,����l���x3i�ł&à۵��`���(�uj4ɀ.s5A$P��*J�LC���TN��c��WR*U��x��m_�;5om��=L��a���k�6�ߦ0�6��W�������f}���zv
�6L��a�����%���a��~��p�>8�U���Ũ��y`��,Ÿ0� ��vwrl����v�;^�)"=�hx .c�v��X��u��W��_��;<�.��2�&Q(�2�,��7�Õ��A�����x���<��J^�ք,w~T�L$��������B��(R߹b~���#���&�I^��B�b[���'����	e����WY��}��'�Y�z�*5��.8n �*��x����5�{f�W_�t�j�o�j��EJ�����o��j+�fʧU{$l�cB��cX��p�$m�&1h�
w����U�`�X��d�f��a�j����setѳ]�VIK��_Ŋa��j��;�d�r��(8��t�$��97�;(���E�M���5������DѕH�8i�r�ه$ܼU|/���O�D�0�-[�:c>ö�uvE��o��Ũo�Q{��G��wx�l肻︳.v�0Z��M��Ӄ�𴓳E�y;�-��kY�������A��.��<�S�S��)�(M�E�R�3���2%7�y�R.N�wQ<�8DԚ�����sҋq�S�5��s6�K�UɽG��Zc\�Q5��T�NgIݭ@ժ��{�?@5�5�5.���Sç��Ћ�w���ڍZn�Y��5�Yx�$Z�˘Wn
7����D��s'�hB��|�(m<ӝ�	����I; s�yl�=�(���fLG��r���&hF��nLqlLZ�����S�=&Ƴ@ǘ|��9�+�by��14�?]~�B'�RgO"�{q(�WۭƯ����l�,/9x��}�%W��~�"���tVn,���A�S�oVax����Ѯ$i�4����NO�7�w�.�����%����4�6����!#���_�7�5���T��S����
�|@�U���l�GG2��ӑ��G�{W��Jg"��p�ZsCKn�]�FU}f=�����%��n��]���Rg�CϞO����7�|��j��H��[�y:����u�p���p�".LO2�kz��-�Us�l����]�+[d��I2��'!�n�`=$ѹ@D��u�{��#D��?ս&�"���_��s�C��,�M>����9�!7L�p6l25U0�R�%`Q.�d�5�2iϘHHy��0�46�a͹W�U����n=
S����n�a�h�6����$˴��K�hOH�u癌֮T�Y	�S	�T��k�wN��vrSò� _��x�qS.,��y�`���=�n��r���g �ڎ�վ�����GT{ �������9N/�P�u�]�a_�� \��q�rr�x��/rj�����/rV��Y��㗴uH�N48�i��8�%�	s�����l|��Z�#j�3��#&�A<�����u&�a��LJK��?���; ��!����2�i A/oK�܋m�&����L�Oޑ&�폧T���xi|����0�)�!���d���!2"s�q���!UÑ�8�
���6��@�����
�;>�;�z��ceX��\�æ�@-��~DMn7���L�`A�5��04z����bmI����Tw��=�Ѽ_:D�Oh^�gLt�3�������@�*�����C�D���)�;@����Co����/%��(�ކ(\�:�����l�N6���}_k����m���Hh���8u��%�@ΦT�r���Γa�|0��	8Q!p����=a������W��D�
8��΍)<xO�q�q#��X�aAݙ�c��N+�#7�^C54��T�>w�Nד�%Ԅx#�}½�.kc��h��k&��ِ��a�4�����cʱ���i^�*���T݃���1n5r^; ���^��L5�G)���Ncn,t�mЂ�����h���LC��M��>�XI����T�"Y5=Kν/�＠tuXl5/�����+�3�|�;��jr�fzc��zn��]O��7SM��5l�c���Jnr)���30_���K�\�TӺ�a��$��������}��9'�[�ԀU���p#LDIn�Eѿ��i��)��ݴ���E���S���Ɇ/�c�^�	t�O0\¤�]���~�l\'��߁���D}�Cow�TM��	3�-h�GZ�SLC������7���~	0�6մ%�W��@��pA,���y���J�N�RW�NL�#n'��@Pxz��]��X�]S�M!^�S6�Ӝ�/�5g.��;�W#O�X��:���s�t������2|͂=cOLk�Ԇ���b�H���f����wLlNg����j8�]� (j;��S[:�[��QL;��Uv��!&A��QQ3[AS�����`.����}�U����c~ ��^H���d�w�zbnϴήQ��o};>A�U�s���g�w�EW�D���)��d���;�I>)�G�3(��{V�S�J�f��7�yP�<b��?�j.�[���͘J7�&��*/����^Ù����ZxKIkY&Zv�-?a-��wR�8hyF�L�-�����8jǳD� �@Ք^w��C@��ja��-��-/Q�_)��]0�R�A��׳{�!M�{��#�BaYD�2�����^�oZ��ʐ�z��g��B1�"gZ�D8����h�Шh�#b���j��G�ix�w͐�(�V������K�n����5% {�r m4 M�����ާ�"E�9eL��V%:-���f@g�����ڃ}����+Է�iOF������)�����qz�i�r�(n�(|H�zCU	���b��M8���D�¾yl
x�����"˯~G|*=Q^�$�D���J��u$0c��b��AyY��ML&��}��������e�����o1��U%yG���,��|�1�)b&^M�w�׋-_._��sku��eCI����EH�o7������j-Q�WxrFtX*�y��Q��F8���:J�n1�5�g����,��Et�jYIU�����z�GA&.�cM�@-�vʢK��[-�l
L�e��/�eͤ�T$���ޅ�bvo+l�t��w	�v$�UI��`��\y'��||�yEѯ������<�����O�GG#�'�@]L#z5Q,�!�,��{�H�4ھ�0K4^3PR%y?f��LE�H��NOev���tJ�p�2�>��XW�,�S��/1*�$z�@$,�W�*��a4ƪ�d=��[��ߖv	c_�n�|�Lx�J�n����C܆���(��f�i�a^�UGC3�!D�����ai,�c�����`�)��!��و����{��<c��0�7��v��ӈpg9�O�F59����	*��Lx�kU	��&�!G�W+ ��d�2d�'�C�د���������k���qV�d\�k���k�@v�J �����`٣섞�/��2���i�i1�V���f&R���PP��=�W��?QU�Q(l���#r��?����j����������3�d�q�C�O EĲ;�����գ:
�@Qf�ǥ��R�j �y�$y9�c]��:^>�!�����-�K��� �]^��bA�����wu�w�W�^#j5E�^�Z�_-�͎��ޝۧw6v�"���z�=��z��f����v��[�M)��N��U�r�y\��H��<Rӹ��&��Fm�l�ճ��˚����ڎ�m���b��_��� 4�9�s,Őa&��(���D�h;�;��F����$Ŧ�vo��yw�W�x��`���zg��y_�@@P. �\)�G"w���G`���c�Ƃ8�q`���b�c�_}~>�i��&9��Z����X5��&��A��#FJ64��}�/�Yw�g,��ތ'l����c*�q��g|�e�IԊص6�
f,��q��kع�2�U=�����)By�~�5��q�wE?��j&FWU�x8��4��g��?M;nݏ�pL��J:nuI��VQt�4<k��p�iÛ�{�Zڣx ��v0�K9u���QSjԠxP�¹�,t�u������x�m�����X��(�AW�-H��q�Y�� ��l ��iR�gY��K��2���*��Pl	�#
�c<��]/�Ʃнt�wBL�Rj�D�k�Պ̨�A��Bˈh�#��r6�!<;ݒ��\��ңҝ�z�C��!��_Y�pφ�M4�����GcI[�(�q���l|�a��*�~��1�����L��l�z��.�gA���y��%|���G�}n4,�����ċɌ�P=	d2c����dH2��4�#����hb2=��U�&��`2�j��e8d��nY�6�m�J|f��w�3��tb��K4�����\����.�R���|�׌F�'��#]ˀ��Kd(��Z����H�b�gLCax�ú?ĝ�K�˒�
 2u��T�  [�Tĝ��=E��v�=����/n�={�?�q���=�awm���{���l��Н�Q�k��b�����\�U�5�Tw��X�A�mr6��mH [b [�X�6�c3rl��3�5���M��C7��֌C�ՍA;ލ�E��R�j��2�T6����up��V�'>T��L�SM�`&�$�Lb(�
UgGd*Q^ۢ�V�G�;�
մ�:[�%�C>��h��1.�,�l��d�<H��M+�e��n+���K�jo�.�qގi}�J鷋UU��ڮ��x1L�h2i��5�px&��h�q�`Z���FD��@�?�47kBz
�7y2��Z�Z�NTV��#u̓aث@�
�"�0����K���8Є@�#e{�j��_�n�F��0�эpE�au�
�yGF��q@5�]�$��" b�_�tt{+�ldX9�"a-Q%�L_c��\25�d�a�eJ��ڕ�jW6��r�$tImr'��O�*䃡�ؓ�$ʻ�*�YS��CU�M��Kn\r������MCG�n�Q��vF��c�-L�:*茽�X#y`��*������	9�����/��F�)�<��|T�\�� �í�"v;��D)FN�"fN؞�CD�Cn�9� �*�
���~�2ĨH�ϑ���ˊ�W��#�rnH����c��=�!��W���Dv��X��Z��oY}�cy����jsK"���2���A�m3��?�u��9��Hh�9���	hCL���-���+��a�������Z�
H.�ߊd'+>tQ�\��)��GNy�(��T*t�RW�������o��mh���L 7Vi�ki���0^4ټK.��k���w���Р�.�$�WO('䱵PU��[]����{���NQ������e��	L�;���/�g5_s��e܌,�77Ʋ�-�M�����+ҙ�m�Fk���*ȅ�	Hac^�bC���Z���r�Z��"����p��a*x��o%�~��5M+X�W0��|�y7�Y
��t���Qvy`�7s��0��[�y �_����E�h,y-Q��ĸ��Z��o�䮈2.FF�%	x��^��!7@�V��j�\G�՛�Mj|�^s	�A�M�H~n�,]��v#����U�*���T����s�Ev�ٽK�%��'ʁ��0��̶v� !��jT9��42�g�C�ފ\$н/t/�>��G��Ԙ�+(,��=�b��	�����:�6Z.�������A���ޅ����(k1D���5v+~�o�ɹ��s���ji���2�$X��(�ķ���S��vp�T�u�mmr �]N�.Zr�^��c�<7ޡ��m,���f��F|��	$���\P9�EP�O{eUp�G܇T�H�-�H��z���W����z���6��,���3aN�Gw|��=�m>^G���G�#\N��b��, ����Q4���KHv�8���� ��E�� �U#�,E�oD���_���sD�v�`(��,�Ÿ�TWS��:9�S�v�Q9��d,h���h%��r�[�f��pB�Q��x�=�0�T�^4cKy����c9vQ������ù(�ң�p��h=���(�����h5��F"�\��O��<�Lǝ�1&H &r���yͱ�T���'=6cB�NB1�w��5���
=���-�W�����0��e�I.�E�S[��2�le}�Bܞ���'�Q����Y����b�Qm��$�G���w���W�Y�*t생��@���ßnXs�'�&t�����5�����}�WΎ�����͆��{�~����Qj;����#��金[�ð�.��[���O �?��A�;�4dc�S�c<�mѾ�h?ۗ�"x�S����sfh㙬q$o��5n����$�K�Q�Nh��l*�W<��X�Ԕ�}�K[S��05[*��y����x][�ʫ�9?�~�����>��b�>U<�Q��`_�'}���O��#��/y,��1Kc����S�m>Y{wqkoO>ta�y�A�� �3߰��sY�oV��T�
u�g��3��Cq�$1�3-���b�3��dx�muk�hL�q����ro�\1�^<���������A-���'&�#�����
�m��n�^�mt>���:��,�ajU�\X&�!O�%{7��a��3Ԛ��l�8�l�Օs6��d����â[�1�K5����̋bW.G�����q�N�>�Ӊ䥟�s����H�\��&����l$+h$�?�F�� �� |�i�ު[�L��\�����P�g���8��1�)7�
��K�{��bC���W��;(Cy*� �_n�s78�jI��r��%�7l`=>f=����B����,Z�x�����{��e6�[��J7]c�¤��P}ccD�n_1��5e	9Q��lp�v�˗ɯ�|T�v�:8�gp4�hB���՗{GL��9P�@��^P�ڨ�4&:����2?�hH�|3��*Bit��ƶ����iT����yu���+]�ϣ �Z�F|��Ѹg��y�ʬ%����J��ל��]�T�JGj�砰��++|,el�9$[?��*��?uh  y��������� s�xe�i߱Y�kqH�k�0M�����"���+Y�^G3|���5�Uu�<�}���B�^zc֥�U�y�ÌŘ��Q:Ƭ�~��Б>V�G#��Fл�~]ǬU�i��^�"(�t�;
ܠ�P��O�j6��x>E��cNĲ��1v�.��-/Da�����g�Y55e&B_D�t�B���U(O5���R�U"J���g=E�i-r�<y)~�HhE���s����\T؊�����y4"4�-��}�
��U��r�$v�4����~M�H��o y1�]�U�e�w,�l+�F#|�C����z(��%����f���6�P��b@�_<ހQ�(Ұ�٥�����rl�	����kZ)[����rlX�/ZwH^�T�fQj��{���'��[f���X�` *��*����o`������'.]�w6�D"�%<�0�ɻ0�@����փ�S�������?�K�n�]6,+)Z*cv&��&$�Й�jZ�S%w�k��ܙ� �B�����v� []��0)��(0�%�U���X�#�VJ+(�O�lh��ь������e���c�U�a���jtk�Ԋ�V8;,�	�Ϥ�N��,�u^��W���Ss��;p�J9��|��E�YX9VO�&���q����<���ȵ���3�Tƴ"4�U�N�¤t�bZ��u���� �C sq���vs浐3/������'��r�37!(���Gk�A���}�#�&��a5����6,���#s[KZ��0�! J��U'�e�R:-����Y䆿^&�=����7�p�S-�M��R����̀�q��:X�T+������e��r��>ȳ��+)��F�ѿB��@�T�x��?��9�q�;t��T["�9�.�lY|\�K�4�_���|�;`�C�%��/-�MX�}Η�p6f�y#g���Cͻ����N��̋G�M+'_�I�:2ꆪ,� {1ֻV��C/X�
��Y�)^��_D��B����A�4z�(��n�"�"�v��I2�*��$��9_���să�$�p��sО�(�~o���P �k�Lr"�W3�1^��x��?��^�W�'��͈��0_Dwq:�`5$��ċxK�V���cuՖ���2Ͱ�w:p_�]�hEh4� �,~U����/6B�g�KuC��4�����CΣi<"�#�hE�`��F{��_�U̦c�!��}Eð*��Gs�!iE���_Qn�z 2����R.�Y�ޡ���g|u�f��'���Θ�K��G�r�D�sn�D����A�}}���'/��2M�G�_�:S���)yZ���c	]�4f�W^z�Ð�����{C�Ȭ��ʏ\�ȏ��۬g ��pG���Eܚ,��$�Tʘ,�A*��8L��n��7S�a7����C�2�?�w��b7�v��8k���>�P���3h����b4v������"�[�ܦ�|չm6>�t��혇F͌A�RIny����{��E��Y�V�u�B��&�9��^[m�\e��Wɘ^���.�C��<Z[Z���½�M�^�ϧ����
���#�T3
/0�-e�5�����f@�5r�$׏��OnVs��l�aRukR��[� �y�3$�!1�t��c��4?5�����3 
!9<w�g^r�r����b�3[�_�2&`�~��(3��k�n)�	�Y��Cn����S�b"����7����!��/
~��w�,�\׼ӕb7ˬ�$�ӄ\�4��ቱ�z���o�{��p��+��{�z�8�מh���b�Ԯ��щۉ-5rV�l_p3&R�3��]#
|f�U�gl�52ʺ�EF���Ue���G���6�	J/K���C�Q��k�V�ȧ�k��6t�Ӌ0��Kf_��q7\No4�eZ�Ձ}�D����DL>_K[�`��x�WI���;���� ����|*m*LN�U^K�ȥV��Y=$yy�1�[�\挶�u�r]�y���E-��wDG�̥3���7�Y ؚy���}e-��u�YP̢��������+Wja�!
:<�+]��?5�vMc��g*����E+E���D®���Ľ��,W%��F?rgUP��J�( ��>G-�VJu�F���J�+�9�>�ۂ�)�U�6L&�k��(O��e�\dLς���1���=�P��LN�?��鶚��e|�i�S��@[��ă��+��@����8$���k*�7v��g��;�:S@7�Q�1pp±���b���AQ���f�&n��HA��^������D���X��=n\$�-��[|�E"%�]�eiQ��~��>�3n(A�؃`�J�}�� 19��]��v��J����V�_��`��l��i�q�J�A��UN��<.k�R���0��7�����bgХh櫮��:�6�7����r�*u��N-�5uo����b��D�y��͝� v"�x�Sn��:������|�ci��u.�[�i�iտ+��9x��^�D���u�UM�#�A�bD�Q:��X��q���Ey.@x�ɤ��
\W�QW#G���oC�8(�Z���E�b���k�qu4*^���k�!z��6a�O��[�{h5:��h�Vc��J�k�V�`"l����H������1�����L�a��Hv�^g�����׶Ȏ�1��u!v�ײ���E.��{�!v�����-l�Ƃ���<	��"�zJ�� ���c����XP�x6���沙�;�M�������碟$?��Q�sTc)k�6��Bj��I(s���.J�� kB�� .a����F�=�K����U���������ʋߏ����u#xw����hZ| %��!x}���J@�y�2�k���v�چ�8I
9�����N���zp��zB��2o�$rk���a�㏒���j�q_�t�y�����X����w��[Q����?��J�\a\������a>7�����S.�ܻ�T�|�(�7qԪi?�>F5�B�!��\��i$NuՖv�w���H��7�������;��[7�Q��;e�?M5M:�{��e�qСr*���������[�V�����ׁ�uҁ�~ׁ��\���\�<���F~��p:���D�ˀ1r0�|���ĉ���)��hO�U�&��)B�Z��)_��(Q�M�J��s5��5j!�<�4�O1\��x����gk*S#[�7 +QR�U�[I�Ej�#!S�R������b��,��J�4-�X���L���*i�N���<�+�Q�t�\�}}��Q�⅗�"�����0Q�@=C��8�&�8M6��Ӂ��I9;а�,� <��䙠VĮ�|�@�:N{aa���TTĂk�Ć�˲X ����0�$�>536�XՔ�6r��`Lqg���{h~?�ƤlD��Ǎ|������
O�'�����n=M6�fB���u!A�@�>���I��s�	%3�4e/�L�	_���4�1lB_�7W�3�a�)��ٸ-��'��ߞ"����pz�[�+Yj%.���U����w��tx:(��/V��3E����J�X'}�J�B㋾�T��y.���/�����˱�R�������$!�r2��t�!\����:���S������Ka(��\+������Ļ�	u�C�Fs�;FU}vKK�������]:�R��C#���_���~
o��h������%ͷg�As��G�%	�(b9G�)H3�ie���l={�du���e� ��S��!J>)��k�j���\ Um�J�Q�E�:P>N�TRڑ�&WUә
O����dݺ�A�w	|����څ,9�F�l��L�� �2�D8��d"�B2��G�}4	�vwK��eL�_�M��~e�2���o|�y����X�~Ƽ�����[��$a^@��:o�L|c��:wOLԱ��TD�'-�6���1a���J!��":���]L\
9��V���E��Â�`E�YU'�� a�K��f(g'/��"���k��aJ���yHE:����� g��L?ηU!�V�g��z㈺�X�����('��D��j���p��Zw��
?��ϰ_����2�e�%��ݏ�1.^���)R���p�~^pώG)쌖��'��D}��<;�}N����h��G;��j�����:ԃ����j߯�y�z^��z;�}~�"1��]t��-�齥}�Q<��ǃP
_y������x`B�M���G�:�l/Y̻����a�|�՝e��	uݾ����\���T: ��{B��wz
���9b�M��C.#��H:k?���|�YGZp�GΊ�+,�ʹ���z�rE�Փ����r%��!�t�I;I��ިX�y�3�b�U'�T8Ur��w�����6^ұ���U�N�dƂ��OB�I`	m�V��H�]�`�@��;S2��\�G�.t}U ���+䏙h}��?������@�~�� e��gIp�i��#84�0c¶w�.�S4|Jk�����őV|�*�ԕ�:<�Vz�(��K��{�Qβ��X*���d;��1vw)�C.E�׎I����;~�����NU��Tn���V�jXXArq�_�'VH4��e��;E[��T�̐,z.�z.Ğ�fU�Ȧ���*�7�24���{�{�jA������.L��9���L��R)����e�K�;puwf�LH:+�;���+^��G����Y=X%�\�O���VuDO�ʵ�,YE���l$Ƃњ"�����R�ca�(�n�>��"-�����k�p���*ǚv/Va-Ѫ��v�[J:�U����$��hx�*�w�@��}���đT����SJR2 FK��Ɖ��QN��C����{ɀc��<x���H�ؘ�9?��-W$r2˦d���N���z�όU��7N�(ԣy�6Ԧ�I����e�xv!z��_�"����t��F?d�Xܑ�#d;��(��Ks�(��է.�H}�p(���ښԧ=�R��V��S5P�OF^�)�y�x�j�X��:�u��g=f
�'
X���ï�@�_o_7//L]؈�����}OW��F�,X��p��v ���T�_b\�����f��L	PE���vǚ�g�f$��J�,����RFV#(�D�Y�0A�����B�d�v߈$�.��q���:n#஋�7�	��
4ܻXJ���y����H����wA$�6�
w�k�	���	����7\U,���(߃a�~T2�3�� 69#�SZ[Ow6�����dj��<TĤ`<�q<F�6�6x�L������N��t���gi:uM'�4md��� F�2����[*UO�
t���!�
c��z� �s4���\�i����@�qA�/ ��39D{�NĔ ��A��C�	�?r��������������_�=�[aC�Xy}4���,�̔�	ů��u)p�w��	��q�D�"]���h+g�c8��.Z}��k!��aHc����r��y�$n��w�^5��H��U��Q���� ���~�2�=�m�n	([���q5��'7���骶�ۯ��d�j3��GWi-�E������n�@ݽ���|=p����ͪT[�u ˋ�����T����TiA>`��R������NP�M>�[v�ǣ��ly)��b�2H֠�"^����nGokWU���2+_j�3�V�������#y�恒��qQ���p����b� @&��q�wE�l�{p�z��? -[Z�YAl�9���r���9Ȗ	���}�tyZ\*=�8�����m�gG.���3g��$�2�YA諂У=�O�5�{#��w��,��f���~-Cޏ�!��N~
�A荄��nBrw �� �wz�O�У�+G�w�@?��q7G����aD�Ч ��A�.�r���R���� W�ޛ�P�T��\�F������Ȱ�����|�s�E� HW9�ĕ6A���+�� �7��;F[}RB�f����jJڀ��ey����[���t�a	��}v[�\�ִr��; ����lu<T�o(���rMF�w ��@WVuU��/�S�Ӕ\5�&�w��U�����A�+��Ц_T?��N�E���
�m+���
���V����_��X���I���&>�_0�����o�l;�l)\���mI��fn��0�+�OQR*�$��T���W�t��!������ڴ���8C9jUՀ�̡Z;	A9�ɖ�r��/}L��am1���;�sg��$V+ћy^�Je�r�R��Pp�/��X����ڑe2Y��{[_��K�[t+ھ���t���d�V���N��a�g��#,Orìu�tJ�
�����Ϛ�t��.���o����1K�>����١�~9f�p�i�ɴ46<�<1�?�x�����
����@�<&|��-� �,8�p��J���;B	!�*o�®�8!��E�&bG)&�A�� ���E���a?�ۭ�z��%��}�&�j�F�C�qg��P$�2���R�M.���6٧Luav>��\�Vc����^�A]@���Wx�k���{�mY���r����k^��8�?8V3e������]&f��%wQ���\+C>蠂�t}���}�]����j:�_M����\=_bLp^�dۭ��"�y/�Z��f��0 |��inC��a�>��G����UV�;gY�[���Ĝ���L�"C��Wi�&$�����(}F�\��LHV�X̕3J0��Mx�Ӷ�� ���wߤGk>�+[��������m����\�C�{���nW�h���WU�qf���V_5�8�4�CkDN|Wi�O�Պ�b�IL5��[ut��c�NL���G��F]�6\�.�����g ���<�[�Om;<��<��Y���jV�����ۿ���Ë��x�'�X����|
+5l+[��$���Ϲ���T.��2Z%�;%o���w�S��f��im7�c,���%�v|���7����j���}-x����ѻ����U�d���,�f�@3f����K��r�-��8{y����l�g�;<�q�9�0�/�ܥ6��6�G���bBo��ֳ���B�8c��g���ɩȇ))?C> �I���HQ=
i��k�ꗿ�����u�`��;�,s�g��*YA"4�J4�&���g̇�5M*��������s�n(G��,�u�������Bm�.���Vx��=�ab���:�gѕUG'�vSso�|Cu(��� *���D���A��ʂ�:�HUX*����]����ǣZ��8ʽ�y��q|����|�D���/OhB8>��ӎ�A�U�R��RU��6�;>!B��UM�?�&*��� ����`�A���b6��lj�0�"���V,�gA��1��c����qi=��5���ƥP����6��q�IgI�:a>]��K��->�v�Z!o�� ���H�}0�h��.������:�3K�83P-��K����!�#��M$�Uf��Q�ֱ�?���f�$�k��mR�GkU�dC�f�Σ��"���'p�>��9�'��ܰ���a�&��,9O`��йhh2N]�?�v;pߝl�H���u�抱���U����|3e4�"��㴁T��5!��&>�|m��'o��7DO%M"q���~~P�@��o
�?�}�m3�?NOcY��l�!�����K�����MoDK����chi�JU� �D�!jI�����ՕX��,quu2C2b��L�3#��&${�����5�=�#.e�����觜i��[0a�� � ���V����6VcGM���_ �`e�#�uP�z����åcq�b�"O��u�j�_琰곪���, �xmP�X���_7h����c��#�"S���+�i	��.�g�U�o$�ag��E�q�|�Rf�����S4b��)%�u6_�mf䠒�v
Q���	�(��T��Q`�|�rwC��~�xx{�A��6��9�5a�n�|�4�_��Ǥ�NI���鈄t�4�}�����������,$����v�<G%+c&�L�3�g_�X?����Bc5�Iw�^u{rK1���of+����\Y���s�}�Pu&2����=���q���UMC�㚉8�4ƶ�~}�{xT����`�G�H���3\��M�v�o��G(eD@0�EB��=Fh�I07�o�|��w�ԥ9���G}s�s�}��v{�"�8�{���X�b������ӻ���Y;Ѭ9k�Ȓ�cW�S�+��MWy�y��)"ʊ��Ӯ�y ������5+�RQ���k�I�n��g�o�*��N:�F��p�$�'^_ï�g:����su��5u����h&e 6�JVMS�F�6'��	��d,R�pS*���:2+��`�*���䞘��c���O�^J������}�qÕ0��'wcsm�+��O>G�B}��:�=1['Fr��Й�N�@�#r6:?�85���sr������NGT�=���V��ZOS�� �j�ҥ�3�u��J�����e��۸��!�s,���Qܛ �i �ߢ�:�EG5e�cy�7�腫��f|���N���-40�6��/cȀj�������c9�#e)�}Co,|��Ή��d�:Ir=NF�B����US��z���'�a������z���X��q���|���yp�2�7,]m���$�Cdc�ptU�N�e�Y}fIm�����	Vˈ��� ������X�@U���J�`��
���9�����8⩟�>��l��l�N�=����U��k_�}�V3f�
�`��&���y�Z����4�Y�3^�M���|�F�'\�Q����&�4���+�; ?���<����FC���q�`Z�c*ra�/[�2t<�e�ua�ґlt�����[�C��GIy�,���y�U��DT�Vc��l���k)���;�7)*s��z|B�V�●	ݹ���y�&�n��j�7�'�C�ݠ�,$�aP"�I��U�n*�D��o������;G�l2��l(�����`�p�C��Rgd�:�㝹?&���&Ag�4v�td&6n].U|����ﰯ�m�yմ����V�Y�7~DCZ��s�-Q��.i|q�ʉ���I�A������~xF�`�����)0�A�|�VcD�S,mU���-�T���귪=�,y�b�RX�jzy9��qY@�x�y`��]똈!��Ma�) %��i0I��~�%m&(1�E�e��C�3��iEp�r8q ǿ�-�*���Yt�1�p|>�sJ�Q8g�#x�Hf0;q�!����>@*O"<�����,4_���C����i9�3������~Rf?�C1��F{��?�>h��vt�J�ԥ�b�2hF8AI��C%bc�<n�| h��%���A7��=B�:�oj��7u�����#&ܨ�!��A�X�}�xK+����e�63���4�_#�\Az�|�j�݇B���U�#���&��;�7��S�˿)�S�zÂߪ�8��/��� ���K�M�V>r.����OƇ!����&<�ُ���]���ϜT�MJ��9�3->K�V��H�V��H�K�����u��Y�TN�F@}ji�������1����9�.��� �0��1DZ�ŭ� �7w	8���}m��MY�c�K��"piW+�]-�L�@�-�6Y�bP�gz��	J�Gְ=5��2ћ��?Xr���\xw�`�l�����;cG�l�d+�;O��XÖk&U��H��x��+��;�®�������}��~8�+�=Ysv+C1JM�%�l�,��C�ε��9*A͌�*�������m�/������Q �>b�GXS��N/B���D{�B[�x�6Ԭ�lˤV�:n��M���^U��q ]Ɩ*��GJ�vڅ�R�:����V�gj&,�E1"0�Ǣ8�r<S;��o��s��!k֙�FW�i�rX;���U^�4�e:``�@3��L� ��aM���c�ʥ�A���j���*��]�b@�OI�ZG�U!�`�J�)���CY�}l�0�Xm�u��1o����0�QU�Ӊ�c����y�t�vՋ�����,a�+�T�<--��B��y�䞍":�W�ɭ��%��s�[������f�ާ-��}]����${�3�Z�J��U*3�0�ɽWM���i�7�QR�<s?��z�)rx��^c�L�hG�<����z9��nJH���eyff+W�?����"����Ғ�R�h���Vm-ņ�4�J)��Mi���܁VP!�誫.*V�gY�UwE<D�BAPDԮ������̝��}~��{���}/���{�k����kοB՝�����3��Ŝ�j{(xj�x�;_���^�PŞ�b��ks���VE�ޝ�(s�����\�)k�3η�g�2bQa�"{�����{��4�afQ!ݫTd�`d�ʭ�!�,G=�O��	���J�.�6I[�-�Z����|y�cO�5=P'���5k+M�)c��x-�����az��S�<c�]4=����HR[�FU�iIs�qJ:[����/,u�I���OS��L)kZ�̔+,]�3]
g�5R8���I��)�Q<~bT�N��~C�~��cm;y���l3.;O��̱z�#��u�G.4]�\��e��嵖������y�i�Hƥ��'8���9���LQ� �Xy�&l�A�8��#�yHt�z�}�'�J=ғ?���Gj�S�H�M�`��ːG��7i{}W���B*n�V�ӡ���D�S}#z" |~�"9�qEK�.3>qb�=8����yϹ�׈��=��g AG�����§��M;�YG\we��Ǻ����w|��J���,.���*����Pu������)
�ysp��R��s5�L�[�w%��e�FT�$��R�<}/e8ݤ�ʦ�'9�uOv�����/p�ᔪw�Ա���z��59�K���Q�7��4I�5�|�	��:�E�����O���ҩ�uM�pfB�[<y�h����ԹRI?<�	�?!��3|m��܏:T�l����PH��%���*�-�S/"�����V�Ӈ�qq��Zw&�v�U[�P�[|IƬ�
]{�����(���<��{��em���<|���tF�q3�[�/ljJA�n����7�=5�=5���
��r��Yx�rI����,z�Sw[��8p�K��m;JR�8��E6ؓ��G�i�"�;{}'�����3���@\�ϖ�j�|:�5-�&�F�D���;`�1n�q��Lj*CTV̌��sf�3Mnc����4c��܌�D��΢��I���ءah�-q��,��h*��(�d�(�����q������OoD[�c������|�0�2F�;E���I�Ӳ��CZXhZt�����]Ψ�C�����AE�;=d�Xâ�J���ԓ�.c���TF��e���3Z��C(NE?�R��g)���^T��8�f)���^�o��6���~�r����\�3�ߡΣ|�(�VZ	�P>�^ue��`y���<ʾ.c	�{�y��<�e�(�I�oofT�c��R:���svy#�[BG*�3�)��g���JV�6��������J+ojh¹��%<�Ot�Y�f���G��D��l��X����m��V�|�"�:~k�c����Gz��p�Q':�������7Yb�b}�=`�m@������h~`,�q�>��?�4�����{�X~xJk&B���`�Ǵ%�����v'X�sY˄��z�C�,��Ɗy��+(�)U!C�}���/���K-?<���_v�t-U��d�Cu�����cv��o��/�'8&����	N8��ԑS���JɊ��V�y�*
��TQ�w���5�a���0�;�gn�����"��r���ƳM�Cϧ<\d���CD_�o��I,�"7,��,-H^x��
~���}�ܨ {�������~c��(HX~�	��D~az�)�B06��:
fR2ݏ�J���?�����`��X��f�Jd2��s����i��&�T_��-�2^dobOcaI���4�~�r������'����ۍ�C��Ђ��w�D�2Ѱ#|5�?_�s_�F$�I�Tta~4e_0L|�ǘu�ً���k�}�;b7f�v|�ǽD1��LL�ܺ�� &<���%!k�"��x�I^�����
����m���~���I���\��-V��ul{�p���տ'�r9�x��k�*uAY=�~{�:9����~_���U(.sS�L�ԙ=��2k�g^��U
L��m��ZY%Yqf�"������J/)�|�UDI�!:d�-�"B&odF��iJb�K��1u�y�2=p������j}(XI˓��δ����gƯ�oH/�@/J�N�b�ynN��.�,�C�ߢ�ة��������)�]�,��;vR���K��s��3t�Z��f\��k_tQp��F���b�j��qym_D����T�y@���ؼ7��O��3�SS���t���8=~�4�_)��5y�,���~=�w�����m_+{�O{:�\��7�@C�R����Zu�3�Zm�
b���2��z�w�@���h�;4��犏Ǯ�i������C�{'���y,����ﻏG��>�x�X�(�}���q&sQ��yl�}�:Z|nK���������^�%�}�"xh��T��Y������SSȡ��#��7-Y�W���S=%�555p,�`A� i��1���
j~���?��_�Ż�O-��\�'����8<s���z��7Ѱ�{갟��h1�7����=�+"�T�c�!����1�Ӹ;�´�����77��Kݤvx��I-v�&��~�g0h��-�
��&��
�3P�ꀬ��T�L���4q���tί_��4Ae<y'�l�"�}^q)CȰ ߻�d囎� ]fj8�p��3!�3}v����,ۙ4�+(�W,�_@;��^�o���=%�n����\&�X߻"T��e��m��q̸#<��j�_��^���j�y�H�L�$��ۆs�<f���k΂�[�,��K�D�t���7�6��0��ӝ�#&��Ӊ��7�Q��w-B�g0E1{�C�����f\C*��X#9�*��j�+��$�WH�ٶk�V��2�΃�;�����i��b�j������md=~��L[��X>�z��!/��A��ob�O���Y��$�?&�[� �<>17e8T��l�z1W��e�ޏ�����i6,���W�f������D.���t��$~���>���&��LE�hSQ42����SQ'��SQ#Y����� �SQ�d\��!SQ��.Ș:5ZjG
|f�zm�K��Y��ٔ�K����\#�x���;�J�����H�Щ2���Q��u�A�Z*_�<��Z"���K0z���o1fmQfW6�s���(�Mg�\}����Un2z���B�(�ʗ�@D0�
>��t6N��	� <�/W3���~������b�xA��%�C�zW�՛��
�L��1��r�nA5d���]��շ��8���'�"/	����z��j�������DR�gM�ҿ�#���^����vҚ�u� �����{��Y��Q���ЉŨ�4����3���$�d��տ:�23N�3{r�3�Dd('�"zI�I"�AD�ʉ�1�ŝ�����|��u7�-�oi*�w�M���9h���)1���*���W��9S��X�$��s��i)�I9��9f��o���[�fZWE�ϑt��"��vc{��9l�?��4'%l��R��R"�9E�Ӏ�P��z/jV� ��5����1ݨ.�J�D}E�����B���dyU7�o%�4Ѧ�S&��_4ʍM�h���{�}⺧�1��Dne+_�����I���Èf~Î�V��g'��!&K��je��m<�K�.Mlp�����L���&d$��!=����QO��Ҿ�l��=�"�R]�!��fw��8���3i>˧���\���*Qt���!����f�-�qb�m �,>W�/����v�-����7�T�Z�]^���������	����E��L�~�yD�,��;~Ĺ;}�~�pum0�g������#1j�Å:�a3|_cI��b����(�:AF�v��|��+�Ou�aQ|y
�h~4O�,��;7���'6���r;\iߴC9i�0�x�P�Y���sG"Jer�zL�����b��$��r.&C����ʈY�q��{���?���D���ʛԞ�8�X��\�E���{Y|!���m�^�ж@/�����n
֛��թ%w_��*׬}z_����Y����Q��c�{ؓ��ڴ1����wM�ڵUn�֭SE|݂7b�kjW�@S��g�n��}������sO��d���B�'��C����������*U�������t�J�E}��i?|��t�2Nl�21�|��������_�{첮߻��4:��B��R���?Xk�u����El��Lnc�y��r��T=_��!�~��K�WK�OZO�C
�|���M���']m5�6g�������)��e�|������S1-I27mO�à?�͡�����H?BS�A�Y�Sf��M�$�|޵��x�UP�J���i�wf�<�����Ӵ�`�6���|/N�a�xO~�q�����̏w�P�k�#ҚCn�y� �=�x�7\k�2�9"�G� �������YZsH��'��Tw���	"܆����0��C\Z�W+L_�f�9�2+�;.�VX}���SP��'���������~�1$H��x�".L [A�W��n�ɻ;�wF>�9�&����W8�s�D��v��Јp��]z��n�����tR��؉�B0��\�G�V����<
�.�����t���hZ�^pO~���D����΍WOv�р�ÔOP�1bߣZ	k�YS���%����3)�g8��޳�"�a��s��ڶ*�3�/H�x=�:�V�'��1��������=����mnfo̽�-�Zߡ\����ʦlr��Y��t�M����</?����_�<]9��1�7}��|���_����.�ϧECtv�!:g� :|�Ɵ�f�����X���F~�y��^�:��)��
�,sv�]q�o�R�}�-v����Q�� �{,EE�8=�,7֚Ğ�w���r'��J�&���m�t�������L��!Ğ�7Ď��!ߝĬh"@�ݎ�,Z�ӭ,b=}�p�z�A���]�mYj��(5N���s�U"��QD�F
��bt�HD��1hr'׫���u����]�.w�x#�>�[���e	��,����cLn����]���[��eQ�$�"R�E�t���l�?���m�˃�yb#���o��z��N�6����3�y^����)�Y�2��& �I������L�%"�͞-����h�����k���Q�s�K����ojQ�^��J/��?�}?���ݔ�ݕ?>�_�E7�{�:�D���ߊ��w��Y�����>�AU
[�9S�T���(��g�e�9��胧g�����Sra}���B�iI�7��Y[��; ��'x��� ��8S�E�=?'�}1\��q�CC�h�a�l��"%��|����̙q.ڥ� �m�T�|�W��dk��Нt��E֜t������ϻ�"���N{WL��Gӟ�V�4LB�WQ�=|`z�N�.��qO��m¬s�WS��,�bk�J���*@���(j%��O	�o=%(RI��
R�7@� Ew��;���y��]R���!)�M��h����.	��N�t��Q!	.�e�] %��VΊ��ʝ\��K�EР�������	VA@��g�'��m��G�@W�@��@	|�P�_n���=v����W&Py'u>sj#�񢓩�\�s�{B=��kZ�ZD��r�P�+�s�}�������bD�<k/�&Z��u���M��ɴ���j��Zu��-���'�k|�2�D��kC�k���O�e�_-��x񏟠F��QYY'�+\$ph��y�}�3���<��`��� �-���,�Z[���/Nα���/�����B���}��3����rM���}Wd�m�d�Ba�����x�}�G�ӅS����
+&{k����I�Id}��n#9�ȸ^���8eR����V�B�xz����k�0��2z�w�0����)Jg�s,��aT5�a%:���mO�нͼAd�����{�,~$V����z���_��m��@��9'|�������q5��7ƿ�_Zw���1/;��؂^;�X*�j*���%�S�|g�j�� ���Sϱ}��C���a��33��[��`'���Mn's�s��ݫy�&rW��_*�69���'�TJ��Рйqd�����1�ۨ�A�=�"�T��2|[��Rb�n��x�ʃu���eۨ^�k��c��k�T'䥝)�q�OX��կ��eޑ�_ᥪaIm�#,I���4�����t 2��3���*:Mѓ�����5���e4���O�L�c��V0K��]�_���S6󥼴��䝘�74�����sBN$�gi������)�M�p���굂����@tϏ�X n�4f}�x�����c����U#�XG�x�ut2��o%�R[�֚���צ	�O���uy>�~j{o*AX��O4b�+����d������һ`�}@Ͽ�����)�b ��ns�g�@;�ܵv���sA�"�
�ް�::�t	B�I�ϖ����P��9��2���������՟NU�d�Q�-MZG8�r�o��<G�����'LQ��\��(��|�7��qY����Vd7����
a���D]WUO�>P�ό�3,��0�hL�rRgU;}e�t��a\��iq�^����G�>VyΚ��pk���4Z^n%��p�{l���A�G(�U�{�����+ÍM߆�Q���k���4�0�XW&�?�\ �K=���&��:��+��eA|0W�@���ٛ�S�����z���G�ȢBqdQzM����>��Gh�9:������\������dr_��n�,h�$�Uȸ��d�o��6���h�����W�p�s�i�3P�wqr��mST�&�t^���r���=��\#����hu���-�[�,������>��Mv������/i+0M*��DEi���*�mI��hLa<r�QL�i����6���k�|z�_ө1��C���nU۲����0��Fd�o؏�c�h �8�M���&�҃��0�]����C��Z�y�>�Y��`"90�F��F�X]��YY���Y9��L��� U+�(�'��(�E0c$o-�!�yb��q⢻O�L�q�)�T�l��[~�熋��B�P��F7����X�׵�!R�戮\��5����8C�tP���U����+L���@ ��[Ň��F��4�)��zղFܦG1PCg�X=���xo��[�	ޒ+(�%giI7�\6�����>����b/�7�����h� ��O�}�Q����A��ۻ�9E��_?w�/6�0�����{j������|�����f6&�W�v���Dj��3�����׿,N�=R���<:#��&���O�y+�͞�3`o*Q�e�;5����\O�|g^�����7�&w��|>���3�x�e�y�w��������ա������Lj+�������]|i8��	�;a��3r�5�S�#���2x�0o��321'OJk5�������3-�Y��$�6���s�����T��A5��U^8��<٤y#���hSUO������V��hM"#��<�%�;������󬧢�~��G��rI^��`�4�c-f��pOM���y�\$m�LM��]�WTb=xj*}Ҙ_���i�o�5����@�#��F1����YMaw��^����$��<�]�����n~�h�~���u�k~B���hkE�H�zh��BZ o��QSGC�|o=�A������R���z�L�.O[G��{�����\���tue߯k��>�'�+�����v���s���]�)�'Ӻ#v��
�.��fhǪ�f
�!N��@���h����3�Ee�h�����[3���ZZ�E�ڞъa�� �y^���z�5{�?����ΐ�^�몈�����wni��ʟB��Ip��r�+0+�6���Zm?�5������*�O��v_*:d�[n���L�ܖ��m�}��[�{��t��������S!9�8�8��bm�!&�;ŰU���n���IX,�b�byϗw�s�Y����>��6ˎ��B
<�f��DER��ơ�`�����ra�^E+C��-�A@�25A�����=&q�UP�FO�A�e�墿�I�`Gx�^/c��5𻁵th�_���k�<m���h���<.����?@�#�/r�~uG��OL�#��x���*�eUrM�c���)�[����È�����������|.qbO�z#�xT�9�y��<a�]�M�F��|�Q��5�O�����,����=�i�7Qm|ş_躿�+��#�����%���������|�y����d��i]����bs�|L����Ɣ1됒S�V�V�l/��ۥr4wD�_&�+�	��^AE􅁟�^����{^�1�be�e���~��t	��4?0�C�gu��+��j���6ǵ�Y(�)�5����ą�hL�e�{�@Z����=��x����8�t�C�Q4�Y%\��T豈w�v�잓b͜�ؽ1���?��d7�:M�I�|�!K��Q����g��ժ��w�������^pq�Y'��9�U�i۩.@��]��ү_A�|�5��N���$�S��|�6���d$[�����9�`�.�5]3sf�)?:��C�(�+]R�޼pn��*�R^((�Uʝ�V�۳e�p�z�ڎ�i�l�������E�ơ���|��L+ q�<3b��=:��v+�[4�~�V��[%k{�����S��x3P�ߙ*�Q����q��Â�}���6P�4�.X�w�<Z�w�kZ��^����G�n픶л�J��9|�W��ᘑ����!WN�}w|2�o�WΡ~�S�Cw�"Ty���i«g��n�6I�LM
L�r礤ξ��d���q��lM�kpϭ���V�4���T��6Ƹ�qtQq"ߵ�5��4�{��oF�1^y�����-�&�pKO�`/NQG���dƷ���L��J�Ϝ��u�N�D��y߷(�Ϧ�_RT(i�]Ēv�9�CwϽ�W�5�I�%I��fJ��0brG��HIi�t3ߙD�4n�z%Iyt��~_?��JK���%>����������,��Y_�'w�񣅂�f:�[����ġ�Pv����u��Y=�w�du����d�h���Srf��L��N������*?��)��,k����N�-���ռ�,�@�X=�x.i��T�A��	:Ϩt��C��ӛ�v���G�kK<�:� o�6k��w�nG/�)u�|� o�B�%�	�ɋk��㳃D���{ʰ�@y�!
����s��EgqϏ���|ܞ֜���s��Ղ�v���=�_+~>����IKܲ�ƽ.�fr�̔�us@�OQ�=L��Σ�Bӽ����W8��8�m�Y�k�i����y� ݚ�˩��U�|��7�343=��4��/���~j9M��{f�|�U��7}�U��2�=hxg�0%�$��RZ����q˻���K8�H��J����}�;���0IG����J�N�c���)����2��~���6w}�d�9	�.*�Dͽ0��	/�fIOE�5I���V�@���h3av@�����ٴ���%�♟`�8�,��A:]=���"���q�X�0W���������s��`�%��ӜP�#݆�9C�﬛ɗ��yDy�'��ğ$�]L���G.�i�~�'B�E�Ɛ8��wr�y�w�3�M���u:�lu�p֤�W����MtBW�^A������{��.y|�319��.5�[,����`'X%A�N��܃��@&Й��	��,9�:o:O`����錖	�K����s�񁴛�=:�`�	%�N�2��˧K�!��C��g��0/;��O����N��#��s���N���T��[=�ʦ��T�Yҟ��]�s1|���pr�U�x#*���/U^#��~�-�����M� c����a|1�w��,s�92�w����%�]�Q���W���iu�����9/�:9R03\e�D�*Hff\f.'f`FN~��c�z�,d��1��!dP2s菙�=�WE(w�;V��4�q��S(�[᝗�)]�8�/A���>���C(w���k�c�{�bG��dM��+A8�)�s�Jh���Q��F��]�(���B�����wI��"�抆�*�v�}�|�]!d�}&Hvm'�o��ł���A�٨U�.<�F]	�逛��L�C��\���#��3��<���(�D��2QFI�m����|�F���U����D�����1��51Y����O��ē͈1�<�������3R���J��"�=�v�}���h����T���2�#U�/��O-�l�C���P|�B��x~+�1�'���]4��+_H0[~&,G�7��J�J�΅XUps��h^�?��H�ss��q���~�_-7h������rBs������(^I�T�������AҊf"�m
��s�O�h8f�r��\a�������i���.�~��Q
|	'�	�px�Y�?d!����������m0�U���7��oL����7�${~�a�����.9�򯃆��)��gJO����r�ϧ�D5����ݙ�2�6���G]�Y��%��2�x�i��U)}�?�'��-I����%�-yz�9��n@N_���\Ns��E�%z~�ѻ���u�����=��_�̛��|#��8ԵB,�2n
���K�E+����)��\��'U�V��$R=��7;&����]����c�]Fy�ᮏO�X\o3�g"�j�]l�FN���KԳfVT�h�H5�C���q~*���ۂ�L�SF$�v��n�X�k�f.Ϗ��� 3ZQ��d��X5����n7�����Z��F�X�"�ՉY2��5f��ț�/k���st���ݡ��h��ʏ�;�)}i9�����?�D�ę@�&�8n�|�7칑����_���=%��um�Q������*�9�� ���#g��!�͏d������q�mz���H�XH������ǳ.h/�Ǿ�^�{��P!M'gZ��}̲#���lY��)���C`x��̻�%���"��nh�z@�'�RYl�yѵD�{ɓ`���5��aKi����{a�T���2�g�8I4���|�$q$�e<7I�6_�EGHm��jӈ���S�o�Ğ�(����p���CU"A;���� ��o�H�h�r\k�v�ۆqr��J\��<���Q����H~op!��7<��oL���d�aaF��n, �����g����@`#S���bЈ��h8�X�܇<����U����t[kx>[��0�CU���5�d}C�w�aV�0꠺>��;I�｡��ᮾ��6�G!�TL��=�J�|�o�UL;��i+@}�l����\�s�z���_H�0�t]��y .�u�q �[�zѕ����K�|����R�~n�D?6K�����r��f��:s�G���h�U�_�]tҞ�������zp��%�D�kd&�?O3b�Y�3n�ءh����{��GK��+b?"����Ub�s�m��������Jw����{�q��o(���O&�����T�PMijN��I9�/��t�[�;Y����*�#���F�x�'&Y�_:]`��|�F����X�q��yR�(��u���&8g�&$b(g<6�3�E��9*�*B�~v�u�f�4�䄟R`�R�6���X�/O�0�QßD�o���}|�7��d��KW�w��@L��u[��[��~Ó<�~䵱�g�j��4������7|���bCc��@�����Ke��;-F���BT2y��t��WJ�'�x�b<���I�}p�{�t �߰8�3��o�N祯r$&�QRxrm��`0O����~�Gi�>�"��y��� ���nR��A� �@���Ρ�H�ִ���W������Z#��ϣ��G̗݈�=THLP��6������,��Zu ��� �m�K;�2��U���U��ߐ�WA���y����A�M���"�DřG6�N���$aI
��6X�|h�;�j�aט�-��z��	���o0�	���}�'��˓�������8w>%9�\�w�z�b�1Ꝋ׆���qv ��k��-���˥�p�~���]�hF�EGo4�v�Cnl$�����h1�3��<�Th��\ng����,�`0q�E ��;��Nvz.�B2�6�Br�89���������g���H�Z��><�f�.�LZ�)�����kS�Y;\���L{�k�0���������k�0m��|�ol�v�'�TKS��;"�����
ԯHy�wеi� Òu�9!��j�H��N�ig7��S��u��ph�ߎ���'��d�|N;�
��F���[:W{�WTZ�yU�&Z[ܔM�`Gxc���n~����:2z�|�L:;˕U����JZzS�B�қ����CO^�f����S�b��Uy��kt��I���/�B|����3��Yg�ٍt@�KG�ބȚ�Ws����Tb�<��-�i�+6�y���͞ST���Q��ѩѫ�V�F�q#�a 'E1D!�ަ��jQ<��F�l�$��q��\�������}2eS�,ؓ�+�t���<�\����;A��e��y�|\��1!�7JH�$�7
�u ���5��Y��������W��gAT�2�8=�L�s��*�i4o����?��b��: ml�!�Nc�C� �vϷy��s��}�d�q:V��L����'�"?�4�s�|ia����=r���WY�J��Ҍ}$]��[��U����w���e޲+�mH����k�U�_��tW\r� ?_�,��Y���Ԑ������DŐ}A��a��YΣW/��D�S8o�_���/��@����`��R;:�����(R�������<e��,K1f3]e��ݏ�����Zn���s��Ũ5'>O���ȉ^+K�C��R��k�AG�Ǩ�j�jq��-t�l^���c`'����B��h��.�m~��+���i!�5����''y�o��-M�4�J�?|rH����9��N?[%e����~�ح�Q?�w9
r--	�D̗����4/}�/�<BSP�
����pz��@���I��Sb~>2���#���d2�"k�2�:��XY�4��3��]<|Y#�k�lF�ö�a!-ˠ"3��=-��	nڧC� $��E>x>"�f�h�R�m^%3w�����ٮpϖ�>�M�����a�����E���5 o�y��Q���
�C�1�~"��}���z����dW���#�����m#��f
����W#�^���a����4��3��G̛�dt֬Ϭz�h�2�'~~�S�b$����V���N�s[���RkF����F6����3i�J\�lM�雪RPHw�2�h�����+������0b�X� [=�Viن|��������hsg�a����?�#�ݤ���O�=�b>���R� �Q�yG�=K4���-�Ȉ��N���ռy|h4���p5�����D��Zi`�6�!X���
֧_F�/�����/q�qOq�
�9!�}��Awd��(�= ���������!���se�|V���sD��E���ֆ�/���eDO�&�h�'��9j��26?k<�­�J�'GWP^��k�s�N��,��L�ģ��1��a�tg�az%F�OcXS�)�#ְ�ִ�Р���]w.��#]T�1B�!��2�*q�H��)[?X���(��|�6P0�A��Y<�,��[��;��~��d��3=��y���U��o5.��҄�JME�ճ��VZ|�o��eL�u?��k����遳�`��|�stc�[{��kYFc���x�_���֎��LE�7��������fwD�\�Z��I����`���7a��SQ�{��J"�_���k��fƆ���[ܪeI�kYX�@M�����.P�>0�-�.P	�-�+0U7���ڮ���3,H��~)�c�,FӗiD��1l@zo6`L�ָ�>�1�ޥ�-�H�0Mb4KT�,��K,�e��1,�C�&Zˢ��s~��50 {?��K�z-��|���=�Ǆ�Јy@g��`����ǖ��F?D38�F<��`�\�pj@k|K��8;磢7x ��X�é�-}�5�:_я��e��q,� �&D����Pܛ%��]��ip�z��ӝ>��_q/Љd�c��Q�p�O���cz��|,�hY�G�9���C��� G0���A�"
�t�����N-{�)܄�W�fӋ�@��ŝ���ݬ��*�,DW�k-��M?�<�2�W$ˇ���_�������t,y�R��#�i�#M���g��7�,�qx�+��'�ԲK4�"n�G�!1lȶX6D"?� ?�%��jhIL�b��w�SQ-��#��a������Y4�FE���F��<)B�t̠D3��3�m����&&rқ���e�O���/�tT��s��3ťH���z�i2Z�M4�X�I��v�
�<JDA�����B~bT�2�_��ï?���c�1���:6�00=�t@"�q��n�@�x2�ڷE��]����������hϣ��CQ����,�`������(M�&���U�"��-���,��H{������[5����f�FH�x�1Z��җ��C9�Q�}ؐ[� ?HF��qH7d�.�B&*:�+db0���]&hLY�;��.
�顮�����A6P�	c��0ȩ��B�m2��z�>�B�5^�\��D�.)p
��%�:�0&U���`�=xL�>���G��_����z��A�k�i��G��
E�����w�u��y�Z�e:�?��w�OŶ@>C�uP�'��A��S$�Gu���/5�?ގ E�>�:�3hֲв��3�á���DđXdh库x�����-Qv��г��D�=׵E��Ivc���7����~�C��Y"�B^'�5' �3 ��y]���=��Q��1R�Libr/֯b�O������k�o��k�ZQ�V���2m�����q@��G!oJ�nOf]u2���6������T��d���N����u�e��z��멞�Ԇ���To����鏤<.��_�:��4�!�h+C�;���j;Om�C�H���������utNE���쒊9���Ж�`�O�mշ�6���>����9$-v͠h6���r<�9"�hy�'d�gz�������#�� M�{��@�D���5��4��4��G"\������[�}�	�ĝ��y�ۛ�6��G[��
��z�u���=�4�0��@{қ��C��1l(�š����l�!e��E<1L� ��:��TTk�>U��_h>� ��]#ҍ6�?�U���4C��j��/��4h�\�6��ھG��}`Xq	��D�v��m��*@�����n�Z���vT�Q�l@Q�Ee¿�u6�C�@�<]�ƞ8�l�V��g,Qs��;�ک͋o�-)�֖pۅˍr�r�@n�G��8�����vEtg�v	�P������$D��m���6��S��!+�ک�>�it�IOl��m�f��h�[?�[_6�� ��[.����@Z��:�l �H��@�*�MT��"�����#�v��V�ֲ�?�����R=Ce��#6hg�!6(ϻ8䝾���K��.��G���G�y���<zZ���I�K�(�x��?�RH�jPo6��
�6	�m"����� �A������El�S<�y�ƈ�QH�^�����-��8�>�9,�5ï�B�omx��gl&�=�t�և��~���+$���0�1����{���BM��S���e��K��|�.��k�1��������R�k���R@ocHzGǆ��8v��4awK<&�[�$^��,1]�U�,����:�+�O���$��&q�D��b�$�Nߙ��0�����+$Z%�(q��~/H�}�J�+�OH�J|N����cO��T�n��$� q�Ļ%VI�%�w��X�|0Z�v��%n��N�
�UgH� q��T���%�%�!���ߐ���$��X'�Tb��qS%�Kdj|RnJ|C��w���(�c���,�T���"��^��#;��&�'H#�ķ$>'�w$&��L�5B</�r�`����ų]"�X*�	)�;�|I���*1Yb��3R����9��J��_��N�R�5gI�(1C�rI�[��Q���x
%���|R��K�'ߧ�������|�+��Х/��,�qiz{��+�h�῔�5]�������[>�%q��}���H 1Y�h��K̑�,����B�"�;�ʅ,��%*7I99+�N�}��Y7H:V�����a�����Q�.�)�m������$_�Uy�R.�5S춺�*�����~���ej�l�r��&��J��|L��b�QV㲕��oS�#ZTcMM}9>1�UXꪕ겚�;mӪ+�N3�a��2����t���*[�|m��v��ᬪ����9��w�nz�&�Ϙ�4�XhI3���5�	f\��ޞ��u�U^V3�V�T�ױH-���9�<��ށVUk���A�RWY�-�X㑛��*jl���o���(s4�����jeB�cZuݼ۔���4Zi��u9�:E�%c�ì�e�;�56�j+[Ѝ%6�x*tԗ+*6���X^�bst��0
� �4 |-�i�́��1d�����e���W49Ϫ��:|[YR]WQ�����-�G�X���*�V'c�T(���������QV��N�R�1�^���SS�t���|�#�!�GɧK�i(����O7j�JX.�G�ş���U?XD~��@�������4�M7���l�Y�g��3&�M7��3=Ι�6ga�������6g��n�t�Jv�3g�M�-��+s�s�ixΝ��ʫ+���Tqq��̙YnW&T� �������Z3��Y;wn���ٜr�͒�>�攕�V�Ա�����Z����y�[��6�崑�V��m(����W��ri�T
�RrN��>Gi�çֹ�ܡ�\He7u�C��Pn̜�R���Pq�Z|�`�u<�Ú9�w�v��Y¦�s��y���Jue#�s�U���7M��g���h�O%l\�[�S
n���^��!kX�e�b��r+)�6�N��	Q��r
�!�>DC|^��̨v(����u!fз�g����Op����J�
�i�&�̮���zT���) ĉŰ��޲�r[�։�5�ߠw�.(,��]��\^P�jjƠE��c$Nwh����OM��2���	�O�s���|c%�:6�|�#����;�.�*��Zh�?�;K�ճ��@�`(� }�_q��ȳ�P?o�lx��Ω�dE��E��"g�MYHu�j�݌�2�d*S�J�ZF
_z��u�)�Ѧ�h��Ŏ�r�Z�ٖ�i56��U�N�Ġ��B��-4�NԷ���r��rXַ�����U#�6b�s��B���"
,����|�BW����pݴ7i�%��Ԋ�kmF'ⲑ��/V+�T�����Vv<���k�j�u���y�f����«� �,�����(�/p�(���Ojeb��U��׫��&�mC��6�V[f��w �����iUX�"�]*i���|�lhVx���'**�Km!y�v��D�4ȯ&	Դ����]�������O[X��W׫>ա�1��<('�]tOm3��K$	.$�a�5���r	/�x&j�����"J�f�dٔ�)��S[��ac�j��<ۢl�	.���i��z�
D{���f���]��o� ��輩D��h��Bb�j�ء���5h��:V�:*FĔN�Pz����J��vC߰����*AR� ̵zxTj��؂������U}�klRG��I+G�5}Jm~M�\U��ɧ�ab��g. �
P*T>F-�\�|�3߫�!���Fi��t�d�H�$��.j�M�yB��)=��k[���'Ø�߇ҢA�I)5U#�zn��\Z9�{��4�+��Hs���Ʃ��}JWk����s���0˫�+�A��,��3�Y��C��xN��Eh�
�4g�p�e�5�9�E�ߍ��N~3�mI�y;q��c�R��c5Z���o6�q�ۅ	'k������.��@s�W9�w�"����N��dC��Q6��,��Qȉ�tHS�5���2��d�)uw��Iڗ>/����;��X�(��Q�W�3���\�R"�ٗR�2��[lJ�`x�����Q}fH/�����4���/$��WS�t	uI���*D��[�u��]�Q�e^����U�~2ʉb-�u���*�[^k�E��D�r{#������O����s��q}5�e��ݚt���_�Q��
L���x�w�%� �A�L��$��[$n��Z�L��N���z=����Tw�|�;~����/������S6IOb��8���;�I[�%}���$���^b�����d���$��J����j�z��.�Lҽ<���������_�Z����e� w<���-3=��_�;tR����]���A�o���m�]\.��7#��ҲR�c����^�����
|�������u��D�ۀQO�7����/���K�D���e���q=|O�^��i	���ZNkY��i�8��N�ղd��Y����e:`�?�. |��..A����B|N�9��9�'�[����/�R`埑6�P|��@��|`c5��W�/����w�(xk ���g�����8h����]�Kw!�F��?߷Z�	؎_3��4��w�^���%ƚ^fl0d`��
�Z����k����p������ԫ���Wl���_c�J/0o��WJ���u��b�'���� �z:���o��k���<�+��x�-!�G�s�����|���Yĵ�ڊ"%`�6Ǝ���������g���
���.����4�!�[�W�� �S��g���e��'�;��q�A���@�=�^��{��� ޶OЩ ��c���˸���o[��[ެ�;��4 3���������f ;$���>L>,�F~ Ҟ���z� ��o��O���>B�~��D�o �>y2x�(;�	����S��>����>C{����c�Pc�W}	م*pl;���|�]��������	?�}�;	vZ|,�	���	,��aJ�K΢^�5�u�6��.9�����o_@�����F�|� '��G�s�5l/����4����zk��{�(�Q�(OZ�3b5,�����������X��
�2N��� ~/��u�e}A��X�O������0�f��w'�[�>4�����4l6�{�5�\�����7�[4���H�p=� <��X���\"xN����/Fx�7��K5,�� ��e�	��2�p�0��c��?̹Rì���v���hN�B�^�V�Ұ��ְ�9	�z�H�)`�H����#ex���"�^ॣ�;�z���-�:�K�E�n���}��J�o�^+�び�hx�Uܘ�aGP������� ��}p��_�2]��I��׉�_l�N�8��O2p���l`b�p'�K�j�?3d��35�Y�w��(��>'���H7�ҰscE9�fk���4\�oV�w��A���9�[��-5�t�/�G��P.(�@�� �V�1_�1��Bg�L�08�*܃�o����t�ȷd`�)"�8��i6�G�t���~:p�L�1��G�,xH�{��� p���۝��Y���ΐ���u�}��-B6�fk�Y�L��~����M���nz�pZ��g6�S&��rQ��C*��wڄ�h����Ο��:���W%�7_�a6���S��nװj�o�.�v'�W���	��a%�E�R`y������?��u�������׉0��6�^�3�n�^|�^�u�k�V�"���xX����Z���x�C�O^�hX<�M�.o�2��I�}���^ F7�|NNo4g��G�;���ŷ�_5��F.Ұpj��U��G��w=��n)�@��BG���#���h�=��j���-�v���v0�O�D��O-�p���M� ��c%� ���q��;|��}��!�O�]=�`��2|�˃4����W�6�M\v���xt-�e�
|�~!/ '>��%]����탁W�a@'����j`�c��3�u��6W^�G��X�?
���1��ǡ��>|��
�1��gQɶ��Y)�����^#.;������������B�������A�W�4,�O���¼\�v ���tL�wdkX�뢼� /�.��h����K�e]��,����[��s[�̷ �[e�􎆭|G�\�l���>��w�@��q�ȷ��?l2����s��S���{�	��9�;�rH�Vl?$d�4p���+�K�!G��^y<Ý
|�c������N�:&ڑS��V�Bxxٿd]�H����o�|� ��؁O��_ �B�L�R�0� ~�a�=|�K���'�p0��M��|-��C�e����RW?=) �:a����G��}J�i��������j��7��N�Ξ�z�'�:����q?k�1�M������ ~|q���9!�ۀE��3�_J�I�s�
����U�]+�L��!���(��wá���\��y�0,R+l`�<"L�1�(����6k=𱾈�����rY]|߀���v�k��L�1��� �x�����k�������܁N:0�t
�ߎm�9���1�g����r���Oi�ߞ��tV^/�5����ܭ7�]���o�'d����Q�]ҽ�~v�K+P�%�$�?��{�9�Z^f࿲E\>�u�D����Ɖ<?\y���~����r�3p�x�� �/�Y<�+�:�o�{�	~�L�������+��f&x�,�9��"�3�/Zdx`�$-�����p�k
�
�l��
��ɂϳ��"��#�U��m>Y,¿ |t��k=���[���McA��s��g6��g�/��r��7�R
|�&���
eB6m���֠��C<�Q��>|�^��|�.�x�C��X��
�	�+~&\Ѳ'Q��\�z�<I����'�'��6��o .Y$��j঻!ˠ�4/����ˑ���y�<o_��e$p�=�,�g�i�[-�)���E��@�[�0P�;�H�p�G��܊�~v�Y#�d�6�Sr��	�@Ͻ"��w�������}"�7�����
p��E�e���As&��1�x��-��G-��u"?+�k��'E�.��I�+���?f`�S"?O_|Z����g����	y�0v`�s"?����3��������ZV�gY7���"�-f�U�e�7BO����Zfy���f��^�{*w����<F�M�ٯ�ޏ4֧e�6����ͲN��������Nnh�� �U�U
p�;"�����"߬@�v����[�ue��C�3;En ��-ܳ���B�(��>� /�l:���ࡃ��1����t`�a�9x��a|��
�(>�����|Q���X��6��P��<��ȟV�U�Zn;��?�w�/5���3����?�:qB��c� �k����C\����a� G}�x��l�R�q)0�+-���Y�>Bx�Z���Me_:����kQFt��P�t'�y��΄�I�������h>�S�-N9�_�ў-�ŷSH>wv���_߃T8�1ܝ��y:'2uaX��/8���%��a���cl:���75��$-�9h�i��kG�K�Օ�Ӫ��aӋ'����T��*�hQm��F�s�M�b��^6jTRn���Q=�JIJ)�*����QאָT��׋�*I�FQ�2��V;��1	��9���u7:˫l�e�Q��w���ko,s֎^p�ڲ��J�S��[()K��N�Vc���/���F# �
o�X�X�0:ʫ�[9-��VV[q}�RWV� ����h�8��֓V���"S!-������a���������,wT����8��%�*��*ʋ���j��1��А�Pq��|���=i���X����@&�g����B��*
��kl�lΐם��5� �a�-��tE�j����-��os��Um,�<�VYV�u	qM(g�\���ׄ$e�5��Oj��!6����0:X~�c��<V��Ma��l��	pӿ7ÿ� �[$����!*�$�A8����K��
z
s�jV��Z5�a6P�c��a��0�,�L���ie���0��e�n��d�@�t��Jđ�C;������:�������	?'��a��h;�r:5�]b�w�E4韃]Bk~PҸ��f��w\��u-���o:襰�<'n�7���޻�5ue��'�"F-V��M[��-�v���_񭭦�Q������!S��f��i�:��A��(}LAۙby�ւvj��cl+�����>'�����}�����&k���^{��^k��	�-���	������w��F3����6Xy+�v�����w�kT�� �=�0�]������p�@��v���O�p��J�ޠRʞ�5��U���p(�����o��V� �� n�/���V��R�<
����'�YIK!f5�c�L��,T�?3H����J��+��^�g}���ɇrJn#����g1NV��7I'�������G�[U[�C�1���4��ǎ�:T�ؔ:�����8v�/WZ�`�t���{����9S��]y�Jy<Z�oۢ>ש��?��5�X�h��o��a����[��B ���l�ܾy{�����v7�v�n�ݾ��6��c�cݳyOힺ={\{Z���1��k��7~o�^��½�{���������3���+�W�o˾�}��|�8�j��A�%~�eK�떂-��nٸ�r��-[�tn�[LU�U�ت��̪��-U5�k
k�k�Ԕ�l����\���������U�Z�^�YS�m��m���l+۶q[��۶l��V��a�k[��m�ۺ��m�mݵ��W��v�w�vF�4���3i�eg�N�΂��w�,޹fg�΍;+w�b�{�U��5��W��鷙�Eo3o���-i�e[�6����}��۸��������c��oO�nٞ�ݺ�`���۱Wʶod=�e{�����]�[Y/uo��}��۹���;�;bw��H�aّ�ú�`���;�w��Q�c���wl�Q��nG�׎��;:wt�;|;�;�Z}��6��\[_�Tk�ͬ���.�-�-�]S[VKw�v�wq���M��w�w��N�mٝ�ۺ�`��݅��w��]�{���ݛwo��_z:ww��v�ws{�{I���ǲ'$�`��=�{����Ôk����UuUU��֪��Ϊ�*Z��Wq[�[M[�����n�ߚ�ղ5s�uk���[�n�Z��nk�V��֭�[;�vo�[}[�[�j}��:��\[_�Tm�ά�VT/�.�.�^S]V����zs������jWuku{uguw5��U���}��&��\[_�Tc�ɬ���^.o��������X[Y��vKmmm]mC�������������������������6�9���N�3��U�5Aٯܹy疝�;�v6�t�l�پ�sg�N�ӷӿ�ۥ�e��˼+vW���]�]����
v-�U��$�}O��=t�~��-PWX�f��(ػtF��5{��nݱ�G-��}�Ag���׀:c1�E1�Z#	��&1 '�3�(޺fk�֍[+�n��$#�^O�{�&���N��
�����u[�����۽���e��sh/����������=�T�5�r�=Q$ŷ'	lG&X��}���+޷���}��µ�����h/��bX�fX�
�WVW������
�ɿ�K��2�m�C�������������s�l����
_�\��p#�uf�}����5��4�>���rV᳥��Lɒ��R���2s�}�پr��l\>����u�w�����40������q�ܯ�j�#��2i����2�2�Ϣ�����<Aȹ4�F*���LJNeeVY��^�_L��pq�n�`������ky�F�������s��s�!t��q�P�q�*��-�R)z���!��u�6�	셛�,�:��[��:3���Ǟkܳ
A�6�Fl�{��L�cmY���knų�+Y��/���6e��=��q%�%Osj�ԩ�0��MV����x���&��H{��˖��1��M��M~V�}Y�rM\�ף���O\Y�,^Kg���:Z�iᬐ��xr���e%(Ke�,o�r������� >*"tMc+_A\}������F^}b�u������J�u!}i��G��4���24��"���2�a��7(r֬狗��[��ʻw-��8Q��7s��MV뒧��e���,u>|6ͺ%-��8���P+a &�k�Z.��HV��a�Yd��g��,lP(�x+�T�ԽS�wڳO)�&����C�"g��G����'CTnx�d�6���\��!O/S����.�9��b���㙞����Ft
��H�E�b4��w��Z�T�x��U:�A�
��0S��ThQa�
�T��
�U��XƨЬ�Q*�V�+%
�R�+�g��lP�^��
9T|�
{T�S�ER�Sa�
O��?Tة�OTخ�
��p�
?Ta�
�p�
�Х�w���nA��1h
g���b�4B��~~L<q�'�s���6�y�Ra��@� ��'/)�O7�=W�|�ʥ挥ϲ�"�N{$>�Q�XIf��JJ���/3�<�t�2��fk�s6�1K��s��	�� �$ܮy�x{�D�2��)^���l�y{��X�3s�R�sO?�Wŗ�3������KW,Y�������(5�	�"^�/,������׭�X��KJ�Y��Pr�r�O��+U�y+���+9TV��8�6��#��=y7�Q��`��q��X7ۙ�H���^��4}�8� ��'�b1IY)���H2�D2��%Zʊ�Ң�+��P�Uh�*�&�f)���Bt����]nI�*4��X)+�녛�*o��*�%��RV|��b~��vƓ�$)+�����>m��*L"�)�����sA9�Ǡi��;��]q���}��!���!b�i͗�2�L��IC�
>��+Ib�~ͷ��H�w%��i|�4ZTк+�={~<��5ztƷ�5\q?꺏5b���Yꀘ�X�pW��x�l/��/�:��vߡ�&9GJ$�H�KV^�JyA箼�4OG�(e�'(�{�R����c�*3{-��A13�'�0it�3K'e�YZ�Ud�(>\���%�d(5�3#L!�	h�~we.�d��U����|W��/��ߚN���B�-�j|���Z���	Q�!h��P���y�#?�(i��R� W��K#�]՘���,K}�uR���R���5C�(w������%�hX�
�0�(�.�)a/K������#��X�b3_~�V�����qJ�'פ���a^Zm��U�r-u�-ݍai
/E7�a)��6��E�Ac����'~e�鐓4�C��g���j�m��G��]�O����e��ǲw9C.�_��Q�I1���р���ҍ�������ժ�1_i.{?v��;�$(#*F2>�@y W*��E<Ø�Tx�&�?�R�p�S��'z����Ϡ���Z���c�xr��%_������ӵC]gz+�/J��r�ژ(t(���KcLب���Sr{�|��1G˛0=��,K<��.ՒNlyP���I�_a-1V�.5�R�����b=i��5�襹��]Mާ/ ��iE���E��*=X*��$G�ǿ��s[��0��Otx�/�D�.�k��Z�}�4�G�t�/���	�y������
�_��f֘N���.5�y�A(�Ɨ2A�+ڌo�� Ȫs��&��$�'i��~���'��b�A� �,�!�Y�A�TV�\��~�VӘ�nX�
���zH$%,��(i*�f`����O��|���7=���r�28x> Q�>B�ƊE8�#�#�ݓ?;8��Q�Q���ߏ��0 h|�4Z�+�<��(���n���B��Č�9�;S>bp5O�yi6/M�>� S�M�E1L{��M���ci}�\^��J�KW��/�}��?~C��_����AF��\�yučt�����%Z����G3��z�3֧��Z��c��v+Vh���l��>��piF ���{�������KM��f�4g�F��k�F,�h�>+��vsM���뽵����;E��� @pn���埣�%��+��۝�i�A��xaP�G�~��h����g��w]�ANT��� kNa���v� �m���� �JU�(���N��E�Y*x#�Nz	�es�R�?�_WN�ؕ�Ʒ؇�b�+���J���½N>�VUb�� ��J�O�B۫�I>l�y�Qݝ�rk��)Bj��t7�\�8EFڗ�E�:!�႑�h��!"��Q�B����(�����\Q	hn*A��AҢp��'51*�5>�d�I醍:����r<�тc��z!;z�蚹s���ސI?`)^�7w}�ͲQ�s�l���=�l�6�� &ĳ��S��|�پ�oRb ŒLK���z'�vK�54��ՙ��&���~�'��s�B}��By�.?�i>(��z����4�SIf�GE�.��L�-g#	i����p��ШTC��� �~�VJe�󏘇���[����)Iw����V��&���Q려�If��1"�mt������%�;G������Y:*�ә���S:!5In�_�x�; ����������]��U�NG(�b�eft��ZPi�|r�(��i��x�m�~y�#} ��C������/q$��Q�^����]��-V~�C�d��A�� F��Xuʹ���/ب?^l�G{��y����p?���Y��,ϹŐ4�A��1�x���2���>@<��f��+%?���:,��W�m�Q�&��_cёN~���oCb$�Xդ����j���哮�_��6�n�D�iJ�Vc��%���ӌ�`|�ו�zλ����#��K�G��4���%,��^���,a}���B*��@ɟ�C�l\J��T�iM�G�������
-v���\��<~t��b̸>�}�{Oe�4k\���NZ��W�*B���2ps�TV�o)H���q��1ڬCuht��j�{/���_5_��y��00�U��+�Y ����>e��9�t>(���J���:�էQw�n�����D����t��M�B��:Hs�ٓ�]��b�$e�!�$�pp&�����}2�)�E��}C̈x�����g���HbJN3��d�>y�a��#gD/O�'Tw�X���)�@�H�gJ�WØ]�K}g�=RG�Y\�k����OM��*��o����+�Kn��X�q@#�w��	h���XZ�m�F�4�m�F�4�mӢYw۴ᘶ��iwb��O�i��K&D)S4��v�DN��z�>?�S]�2!'A����V���[�Q�<�sWM��z��_�&G��z�R�G.�B�^�=�U��p�O�<=�9GZ�;V��=����@%w����6)�W4
Bbӹ+}�Kp�3��_r����?o
�^��W�W4�g�#�4��l�X����U�Y.�OƯ[�V�]�t)�7�w9��v��F=�I<CL�����+���5ӱ*��윭!���J�K�c?
�h��/<�K�]R�//�q�B[�x���/���^�i�����B���7%��2S]8/�G��8C2�jLR���1s�
��]���Iן�&�`7�4�<��9�f�aX.�hذ��0)��'<A�P�	� �,Ǒ��%��1Y(����p2�Iԯ�Q�UΓ�r�/oɲ�R$ne�����.e���)NwiXc�d��V�y]vN�t����S
��d���g/�1:
�G:��dtd�g}s�<�c�"p&��!���)_�N8�w*�q�,��z�Vʸ(���"�[kt\fYz,}+.�.t����3��4��10���3�GD6g|������%栐��Z���Iٺ�9AO2hY���H[�٘�A���?�dcE9#(��y���yK���)�b��`<���7�3�i�XCHR8����7�� ��rF0�)g�@z�5�lYQ�¤�3����Ig�P�4�D��3:��,����Ci���6�=��<���L{/�(?��z����Kl;�O�	�.��J�Wt,��hq�����]��+?�_`���+�J	��y���^���׌���<d�ߡC�^�W$�ca���y��/��"� F�wlИ�28�
$�b��
�HV����D����\Ƶ(��Wb��q�&�U��
R,5(E��HIo��;�/���?���k�R�W���x:�������B��QT��P�:_=��wǰ��_��8�=����\Hr:3�\�i,���9h4�q�5o/�{�(8>������i|)ZU�)g�%����2N��U%a��(Uѳ�ì}f5eeD��ͺA�ͺ�t�xGS����tf���,�>ǒ�,H��.�8{��J�j��f]���E����La�w�bp���o~�XF浪L�F�4�4JI����O������� �y��k���!��>��)~��%p4�*a5Qz���&�x���Ͳ;��X�����7��*��M�U)��k#U��ӳ���_0�Go��ɉ�2r��u��Q:�F�d�{u��)"K�g�WY��c�RؓJ)4�9�j<Z� �2+ؐ�~����Nt%�@+K�d.\X��h��X?��k9�kӵ%�WܸW�,���ߒ��b�Y�����E�uͿ���# 1�����.�i���t?�� �龖�8�����u.���[¾��=3w�4�AX;��F:H�G�
k��I���|����/����ڤ����������4<Yވ��?c��a2Z��#�t[� i��X�J<�w�����6`_Wt��t�I��0T�i	3���������$q����3�[�P�%�-5�����ˊ��E�;�<ǫ3�ٴ�t�w���`k6��$�Rf~�-=�xT��eβ����������F��F}��2Y��_�Ck�ˑxW���'�*�M��V4���*�V�
x���j|(K}7���a�z��s#�4���j�I7�����!$h/��4\�Kp]v��I�<,���1M��	in�w�	�8��V�Uf�9�=�4��K\G3a��{�(ޝ�&�Ԯ�9�9�i�#��(���7����b��9f��q����}���8lF{�5�]�:������f+��9F�B͔��7���N��5'���b;03gn�]�Npy:�v@���%Fz�{|�� ^1�^+z�"��	��b�+��C�
����p��Rw��R��t�w�6�g�Ϗ��(|��g|��3>9]��I�sZ��+6��x����-���vM��5��~������owFY�
�d34�g��*>0���|�l�t��6)�m#�M-�6�iݸ����y��m{ �)���]�ʾ��0�y[j��p[��WE�c�v��(!�s8/6����/fr�A�ќ=�%=�2�^������=�i��/�����U��������ǩ���?P���P��d%�0H����z����`�ٍ���p�]�Їjen~6��R���M�bxk~�@�B �F ���H����\�3�>��Wp�m-�|�q���̭�|w���i�K�	.i�A�l�����׏�3�)�3�q�B�r@�� �����Lu���#��(��4b��&�hɖ�1��� l��LpJ��pd��沋��sr��n:��!+P�H�����Ǎ7 ��|'���p,�
<'7=�Rm��HY!m��v�і�]V��xZ*~s3��Z�#Ʒ�����pL,�,ޯ��E��v��X����)�2���_"r�d}�^VH����q\��z��˯�~p"g�z�ڢo�ן�*	��~\�>e+Q&ѯ��l�fJp-tC�zH��L��jx���@����z'���/�CqOĠ��t���PJ`[�[�nU�n����#-��L�����8�4���0�g�r�k|�&z��rR>
��]����S����Tb�����`yw�܌��i]PG�à�U����K�1�z���7��R�8n��7��@�Y0��]0s��y��_K%*D6`It ���-�`���q���jH��J��Q�>K�ȦȲ+#�C�4n+���-�.�Y�c�U�Ə�>a�@�d���
K���ӧܧQ�Ogi�R��Y((�uִ��T��&��\��SǑ�֍Ӵ�x�z�IgT���[8�le%������ϝ����P���3>�����������Y�������vvV��PaܤlJd^��W�(�la����F{�0Sm�QJ��̨M�H!�Fx4M�Bkllu[e�(P)w(�%G�F
��|�H�b���@1����!�Pd1[:,�Qf�Z�<���]�Grd�it�.7�ɵ�6i�R"�{R	Q)#��]36\����c9�x#6iS"�Ycr�@�yG�����M�Q�8'�+u�}��7������K���1�c��~���8)�:���q�B�q��'����g���Rbd{���1t���F\#�KWa���@� ��D��;��I7�u�z�t�Hd�q���H������=y���p+D��N���l��Yk��������6VX�c����^#�������#B9��,�j���#o��l�7b�3޿�GN�L��t�Y`:�}�#a�õ��;b��}����7o����+h�_��k��<�1���L����j0��@(l��&�#��w���%���]��9'���+�EA�T~�)}�5�An��~E���'��9	�qh�c(s�u���2��Hx���ҭ1�~��0����j�a͖:.�(��)𞤇za�_ 
M��r�J��@�p��X�/=k�~ܵ��F�<�!ߋ����������?G���GU�x���N��2�s:ua0����쀻,55������u����0(<��i�0�j͙�&��\(U<�/@���4��/�g�A��ܐ/	��2QS6�#��{���\'zubc����9*y�Ɔ�7Ʂ�ρ��Y54GI?J��l0դ������ o����Ub��n�Ig �X�A	+�tȆ �q�Xq	��V�If�ȴ�|��_gs���Q�J�F�͵��k6]w-4W`�؍�;��i�Ƈ�JVͪ{�Y�Y��IN��Z��(x�b&��M8����\h�#��@
8��(`�����ג�[�i�I[�Q���d�2��M�s�Q�V��P���ldhC�J'�=���2;uK[U��
y��@n���Tz R����6�Q��Vf���������C����ŃQ	��s�,�L8��= �ݖϤ[��&ѫ�
��,�%����2U%Ez,���a�H�_���"�Q���P������b�;E>�A$MO�����.%�9d�4�I�q��6��T�Ls�Ҙ��O_��>��ŵI�{Ц�'x�������0a��0�Ǿ�UJ�fx��\�����'B�7'���9DH���)ܑ)�x'��i��7�����6�Cuy���{<��;�wh]�wp�Iod�	ox�!��N6��"9��K�����n/ۯTD���t�Q&���1@��=AW�t��7�s>�d6�r�Hz�p��!v�:nL+����$ӟ@s�A<b�	Z�]�	l��(	��iah㰽�	G���$r����Л��T�P?G��3?��' ia��o��	�n2@�"�������6[�Y��$�M�s�ݝ����Hy��,(��K%�����S%%M���������6�OT���yځ��_����wl�J����WP>IJ<�Ό ��*)���Q���hg�R^����m8ׯ��XV
�5�zA)k�7�·�˲Π]�N wO�8׹�����^N7��>���h�gQR�^�59������#�#�q0�Lh���]�䩆:��U�&m�c;����2��鱙s`���)�u:9�<��D��N�Lr����b��:
�1샚�b �9��V
�a5'G�.���7E��ɜl$g^ ����A. ԼG�� �n(�S�#�uf�H��1���X��B�[hfiR�Џ�*��&F����J�����W�GN��')�N!�>�ܩ9If`�D<)|R0~H��ra�/���l�i�x�"e�t�;��n�^�G2������0|"���<�a#6��S��R�o|۽1*�E�f�����D�����c<���Ʒ�^a�DG7����*.(���CYM���W��W���-Z��z)��Ჴ5�o�.K}��QͶ�����IX��� �Ɂ���b�[]|(��هI�H��V:��I�¨IL�cR$��Ō:�~���S���1,���ǵ<���+q��J*ϼ�!� H�)��?�S���r= ���b��ՀÆ�����A��b,����DH͉.)B>��K���J��0�LC�t�eѬ�&�MY���Bs��D�d;/D�8ϧ�F���T�h���e��b\�O��#�MY;���0P����n̫���5��<xZ=�[�8��u<�r���a+K&�a�7Y�'ך|r��iu��Ё^�����4���#[t!��S��g/�=~��$Ρ o�M|�W#$��b��_`y&n�ǚC����v&Uj*�!��G(hn����i�����[K(�Z�M�����Ib����x���2I{<	�a�d�X�h�m�p�|�M���Z,��_��gIݯN����<=��ٮH-��P
�h����X%�*���]C$�<��уα��f�Q�i���Mz����ܧ�Ə�Ĳ4b2�3��J=���C/O�0ѱs+JK=�6q�V@L}j�N��5Z��粅�;�	�����/��,��������jO�K���d�^\��6 ��L�7�Y����3����V2=�x$�E5H�GZ��1�0�`J~O)� �4Z��lR�7���j��(��K���6���[r�`�%gi������;\���sb�V�/u�����X����Sd�g�g���Y�&��25	�Za��L�q�^j�X�n��A��=�^h&cE�wlX����M|D�΄#6q}�����{h-v|��XıXa$L�����B@��~v�%����
y>@����s�Nc��=t����g���� JݬOè��J���΄#4�j�:��t��l�F�!<���q�zO�78��zt07VT�d���甬��}��`Y��Q�T��>���-��/*�푺��XEX�0J�W��!P+���Iz@79P���PQ���U�{j�~�x��j������1!�`�����{@�HWA��~��5&n�ǅg�y��)<�.ǼI�����,~�߃�x��=�\�,���c��Q��8��y�������a<��r�䗾y)Y\���@PŦA�1Vh�����d�IŁfp��	�!�����{�|�_�t��"�-��t���Kk��%z�<S5WQa(g��(�&�=*�?%�A[�>�MO|-�sp�S�(PO��h��flt餢�h�&�����z$��-tW�i<w�W��&�%�l�acŹ��A�ϡ��3����޷����������X-�������v��Z�x�� � �T%Y���������>���]���p���8�^�l^@�g�s�&U��u�cL� T�������wX?��*Kh!Љ����\�����5xbYI���{:n�;Ԍ��l��=qe�T[�0V�AȬ�9tO��4��+?"i�U��n��5,�fAop����8���tV&�Y���\��\Z�?h����e�e��S�)�r�u�{>�4I|\�a�T:(�=&��iI3iյ�&��9V�L7�U��=x�h{��+p��GA���<=��b�fF��m�gtܹeoM��c�pg��������lh�j�u�q=�����>����m�m� _��Q�E~�E�h�� ��pT��E���~� �^�	�N 4�wg٨>ܫ����~�ԍ���Jf��˙	6(mPڠ,�AM`���Ҙ�T������+P�ζf�)�ol��ھ�Mc�"OJ�Õf���Ac	�ԃ�=<���;hqw�G*��q��@A�g.*u��F���{h��х��gd@'aL���hhG���15��
X+E�w��_�>�Ws�x��4��!T�{���`[_̅���o%<��v*�FTU��~*�k�g����6�]������#���˿�0�W���7�Z!ā��Mh���zo1�}M�Ai�e��f 3���\&ں��Wz�|�j�������z������������G�6�o7l�F��w���k�(���Ub��!3�5T���k�A��m��1��F갥UU��K�l�g$7�qܛS]�,=��PV��[,���~�b�F����:�I_��|v�U:� �L{�ǓJ��+5�I���:���N��a�w4��������@�W���N��6D�	�F�Ԍ��֣��0:��aa ��t�zx�o��vm��e�0Bj"���a�	�����u�O��)Zx+r����7h@�������I�E����9�Ai�7�0�A�� �JSK�1���/XP A�ۓB��=�]Hq���`<��pL��"���M�r�7���$�b��5���Z1�������,⬬�����Qx���{���'��:G�fj��TN��MWp��W8dVp�b���2��P����l'ZQ�5�:�͍�������]��A#�̵�>��.�p0O��4�X�yy[�Nnd�A��蠿2��c:W]�P��1�*2���D�RVh(�B��а�0e�rEN&�+\�j��R�~g^ 8������k��U��>�y�"M\�;=��q��<tm;���s�i'L@AkY9�X�ao��N����)9Ϧ��}����''3�A�d�1�H�جݱ�N��C� ��mǢ��@��^�r	4�J���SB[�,�3�0$����J�$�yM'��)<+6�gn��ԩ�b��-JD��0�3�P�x�3V��@��bM��5)��ؔ���)���P�2HX�2�X� �b4VT!b�������+�sC$}��_�'����~�Šs<�V�b�J������jH��:�J�St�؞�����򤿓Y�"�N��qZ2m\8JSY"]���J��=~c}�c�O���8$1Jꔾ���z����C�N�9|���w%k@�y6�SM�63�m�Cs�צ��Z}$y.��"3��/��@6�ɏn\�Ƨ9I�@&2����x� R�Pve�0���PaR������ aE�h�
\}���
@��uZ�\xb�NT�����+Yf��_��cq�U�딈�=���N�Հ+�y0�����-|��4��
�bH.�&�t��fKJBj��
�3#�Sf��HJ�.B��M���t��q4C�3*Z��O�T�����dyL�&c�I�a�,�&Y�M��5�o�M�+�$��$�N��'wR�K6o�����<;P�0:�r���`��z�E{עX�����6��&�+��	�;^��d���W�t"ީ�W��t;�f`�t�~��MS4��IZ����n����y{ު��q��3�F�E�.��>]�
h�q���<�	���nꋉ��V�����/�3�IϹ�Z[��󫊼��_�T��S��->��d��-9��v��~)ɣ�?��
hN��v�u��us�����G��c�����}�q�A�1v͔75?��}Qŋ��u��D�Dc��5׍���\�d=#K#Y���lP�Z`|�Uf=�VK��[~�IVZ�c�aM��ѿ(<NW�K�i���do�8͔)���'������$Jt]�@x���<�>m��$~�����pg��^\��J&z�kS�����%��q~L��˒>��c�i��ysǬ^<��2|R^ϔ�S�U��l��`\�uD���p}'$O�R%c�$hk��ҹ,B��������<������u>|܌�0\�H�:�iΚw~��"3x��{��rx,G�f�6��˫3��5!�kA3������	-q�pD0��"H<"�BNA�|�)����<-�SR��u�����濲]��ߣ;R�yM�����3:��d{�7R��,���Ir�F:�uu<��'���'��A���k�플��S�@�a��{A^���d���4�V�;G���e����^�ҷ✔�M2��''g���y����N��XA�\��5�Ǥ���]\w7̅G��=9nܗwN�D�_�10�00��8M�i��p�i�BTG7}�[�ȸ(e��ut�NZG�̏IE�Zbm��zQ+��J�i(^�d:`N?G��|��Q;�֢C��RJ�/r|L�EF/�q_�E�h� M��qb������t�k*9�J��s�"�?F��Ʉ�L�y�����,�_y!��li=QY/��O��?�J��E�5�x0x⸿Ȼ0���~؁�j�.����&ЮQ>y��>ؚ#�����
$�<e���p�u��=8��_4q�1��0�b[c$����߂��ohh�`<{)���nD:/��H����A�6#+��8rw,�*P�9��"�K�BXr)�B⦿�E<�WO��s\�:ia���±�f��w撕@���ұ����%KW.��O��13n�Sq+��gƦ?_�|�,�[���iK��c'��8�΃���c�ψ�o��4���M_��tl:ޥ_��Θ�q?/.[����㖭���-�<�U���R���+/+����Nz.��,-}j줌8 q��O1�XZ���VB%f0����轰By�47�Ǌ�%%*�Soi#(��Ĳ!%w�-|��(BFĕ.ShL�y��J�"�&*��7��uSҖ(����X��4�OM���J�N~�Jo����i+���7�di*���.L�
���^�S�a� ���kސ�qq^��4�d$�m���S��_t�븻�|W�AbaJ(�O,�
S�1e~(��R^G!��MY&�*,Y�d��d�߹�4��iKV>c_��2|Q���_2Y�-��G�q�R��"���/�h߈V�;��Bp�]���G}�'�'����>)c2�gsi���tAq������K���E���Y;��~��W�[��0׆�|4�T�b%>�X��p��s�If��8�U���m��ON�g\b���e�Qx��'�.U�s�d ��}=N��eڿq�����zp:�x����S�D���~�>�
t�Wh1b��{>�@�i;.{�*d�ю�y>�IWyP��9���Zݹk�}	����op�ē ��5�㵬�h���_�Ζ��$'�Ð���7F�����o���$� 蟀�-����O�Jfa`�Dn���,�b�{������=���-��O�4�\��/��*<]Z�������b�:�sa��� #&qF���Hk�o�q�W٘�9JQ�ӑ��1֟ɥ�@�m�M����4"����UDܟ�-Ҏ�����:��ӱ�!`.aC��BCx�
�b���>��6S�{��*��r)ݻ��0_�R�%¹Y�~{�3���]��]��>ږ<�>�Q��3��Ll#�`��u)<�-��-B��%��Pu�}t�ӹ�C�E���?����������a�Dlɝ�$�qd�(�
Xg�r�&~f4ַM$w�;��L(�$���H�p.|"բgm?fkɸ��>_aF�ՙq�Z���P��'���d�l�u���g	:%y>����+�Z��8|�L�?��;J?�;�B�k�=7@Wxo?�l,e�3��!d���K�����&e��X��J�׆}
>w�S|�[�GeG����܍��nT�v3i>P EL�����A)V�ٍ+`-�$V����L������ �b�,��'.�b�u
�x�� �-n�#0�� �	�ol��ܒfz��md����>@��J(�Z�����x�]����PQ���Pz�~:�u{Y���si�.lqc}��������w�=sMY�N�A�
A�v����|%�p-D�?j�ob����B\~s:~��V���;�o���=9���4ߞ�k��d%Zt�t;�a�+���#��Z��/_u�'���̓3c:�=��r�t+G-�N���6$�c�, -c�;�����ܖT���2�,�H�X�
l9��J;QSm�6D������KR�=�1��~��\��I)e�B[K��<�k��1�L��ۿ4�"VJ��y	�]'�cuw$�L��Ԭ�w�qR^�� �`���%B!��x6�1��xIh�ɳ��/�'��2L�g<'���[kA�F�H�U�Ն���Z����g���	c�pg�C�@�ו���l�-�^�S_SR-�SBy�)���O�J]�R�������j�0z ������.P������'Bӗb��U�o�5�CY�����ީ7ƭ�!8�;�������n �+?�o�/�ѳ���~:� �y+��T�ۡ��B�k�+:������ վ媿���2�2n>�u������M����������.O�-���ۖ�&��$�$&��\!��m)��I��'t�.�۽��,M(�υ�NM<���7����p,a���m�2萂�U���d �%��遹��e]Q���(ޝ](�g��5��N`.ť���y��؅���ch�nT���V�:���Q�H�>����)�?_uW�­t�6v�'d��sp� �=�Ў���7g\��H�H{�Trͫ�ZT�"��a���_���8�ކ'e �l�Xk�fAフ�G����v�pg��8aܹR���3X��l�θ��S��ˣ�n�/�ѧkp�e�95jQ_\W��7�gk����m����?�s:��q��S�0(��4��{!��*�3�u�ҥt���E\A�_�l����V�HT�HE��S&.J'��Q���E�\�W�	47�J��kI�qB���a�C�1QpmF�'�Ǵw\�sD5M�Q��7��}���0$�8�����@g�Q#2�*6����`����S�X�w�ߛG2\l6��C,���<v~�=CI�REe�<|��6:_�����(
���Q��ϗV�}6�+������R�i"�`����мເI*>:d�>2�O~�>�
�	ǰ虍����w,�«~$�]����Q�:	�tA4-���%��~M�����ezt<�����d`���ˇ..Dz��C�|�,g3�[TQ'.2,�U�:V���~?^�8�W8�$�}��$,<�~�7��} 93���@����*���gSr^ �� 
܄�\�~��� �ؤ���8���ʝ7��c%�����x�X�&�l@`/��LB����om@����C1�o;��\C������)�u?f��
-��褋8"maGw?�sc�d�8o&�<}���;�-?����^<xz���,�b�ă1�^��H�l�^T�/%ыW��a�_S�U[�bqц��J��ѭU߁_��-*�=����n���*ˊ�2�=݀j'�D/4a$;gM��"}���P�@vc>�ħ箹���R�W�`z%餻.T4�Ѐ�^-�`~,��&����I��ϡ�e�(qL���a��5�����#^��4|�Ti
F�,)�р\� |y�v8��[k��\z?^�8h���|bѫ��N�>9�Q{����;*�x��[��189m��/�3B-�1��h�����N2����&��*�n��E��n��ע+3��$��Hy�����q�;���?Ã���s����:�]���p>��ď+5�y�Bot�� �`g^{N�F�Î������-�4쏊/�zP̀�u��f�A?+ϟúp=v�?�x�� e��`~u7Ĉ��0��ԅ�B�w@.}1�$��wX�6Tٞ+���4q�(NHɥ?eӎ�'�7��q���|��Q��rg�ר��WEA�*U�l���R�͑��ri��7��J���m�ɫ�D��X5{�y=J57`5����HI��O<"���Һ�����Ea*�-�V��z��0��5ќ�cRʓ� ���ϡ�f3���O����Ӡ�-R�I���P��5�t/�,Di��ϧs�-֪J���hڢ�z9�];��^�e�7����NUЕș��|?|[���b��CP��V��b�؀/�s�&�����!��M3 D.�Wr|U�	�x��R��p���>�ս@��y�}���ot��K�\��*\���*�Ϡ�N�z>�Nܓ��c~"�~���Ȇ�hU?����4ˬ	Jd+�`��
1�t+;4�h������(8`��d��Xh�P��;F-L�_ŚɊ�qj��?�8��PG���X��U�i�((�EU��Z
.�m�n:�;�ѡqW1���ND�r7|���7%+`X\g���9�aHXC��AfIx����sK�g�E/�E�w���X���!��� 5f�BxI�ߨ�
{T��
{UاB�
���
��0���Tx]��
�U��
Ϫ�s�S�*<�����У�*���
�T�W*�Z��*�P�U�'*��
���
;UxB�'UxJ��U��
Ϩ�K�.6��I�nT��*lVa�
[Uئ�C*�@���#V��*�S��*|C�o��-�򃼠�ސ
�����G�>^T!e5�t�f�����	S�'Ωx�*<��N~��v~��VT�K�練�T��Z��dԂ����9i�&���|�X��5�^�Q�j W�a��(h9k>��|���Ze&�������v�Q�U����P��=*�Ua�
����*��-��o@��?T�Q�*\��5�����c�4�J��uB�֏�^�9%���!P~QY?��M��bj�4��[��J���8������6�O�Y�!�����e���~)�tW��y³�K���>����nB�cx̬�TB�d��
ޣ�
��Zo[���}1����ݿ~B� M��'Q1x�[y��U��{��z����#�Ml3�$=�mY�#��s���l|�؝H|k�C�6ѯ��4
����~yӉ��.��� ����_?��1,�l�����~5�<�
ej�F��f�vϽi�v�(��)��c��n��-�w#}�;_5�ɗךPRg�����U����)f+��7f"$*ŀ�5�̑�c>���Zy����t�"�|��o������6�����uR|�b�؉36�������#}�f�5ŗ]�P�+k��x� ��͙;���C�L�����Ǽ���#Y���+_:/^4%��$a�Z���^�=p�B�G(+�Q_ ��J����Fň�bx�o~O�y�<v�D�����E���퉔[�!�3����I��4H�G�H����P�������b:��4^mWls�q�	ר��W6�1||ʄ-�1�Dc��׺��X�ى�1Z�J~������O]s���>V���WU�wV]sB{e��ޣ���Xc3��������	.��ϑ�0�|���/G.�O�z�J��-q�Źh���o�D���n�?�5;|��j禇>����z��V��Y�e�&���v*�3�߱S��Z�Qgw�p�\+���x�Ea �;d��:�M��~���S�9�[)c��嘘y�1���?`��08��� ��IZa��k.0w�X(��	�d]�!Z˭h߸q�b����:.K�ǹ�a�Z-Ee�|ۆ�e�f(��U��;ݎ6d¶{f���F�+f����&(k̡�1/���י�ُB�O}�d����Y��\�5�$������,
'�μ@�U}�.�m�
<]�A�<�R�$�C���]����׿�F��I��_��������d�P�B_����ؖl�)�4և��{��d�L9���d��o̶�v{�_�h�w돌i���y���Z�E;�4�|�4�9L�z���|�������`�� ���K0�+�W{9���#w��ԬJZ�t�ʱw@�r�?� fa&��;��4�̱)�*ok̥�
��Ւ���������|��A2L�`W���ʫP7������VǿrO���10���1@_�C�0����`�߫������E�)Z��Y��I�l�3����p[	J�����_	�$e��^�ft*���-x�Y�6ȾW)����/gz�~T����<^Q�3�u�A�(�P�~׌�����c��_�(��ܯH����Ѵ�8��T�tW3����c����5��'�*�/\�!ܛ.�������>'�B$OO�n�h��l:�+b�x)��ҟV�2Oǉ���==��E0�N��ĳdF8Ķ�%E	��G���V��z�EṈcž*��������B܁�����XQL=�{��[�͢�;��JS��|*~�[��Jt~�,��i�~Z��]|���H�O�2�DL��g���Nf�n�3�l����HP�G?Y$WU�%�}E9�6+�Z��@�h��]�+=E�7ƁX����T+_̪d��o �* B�[0����z%�4T��t��s�u�l�a$|��(gN��gG�@�jP��Z��A��I�\��$nw��*4�g>��^P�ͷ*��������s�%��V?�8HS���.�*{�AQ�!â"�6���}�yG��%A��at0f�
Zh��¢]**kٖ��
�jTRJ+*�H����1��X�2�ι�3�H���|���7z����v���{�}���>�ӷ́ak�]o�y1�b.P�j���P̝qw�*x]r�I�F��c���v�ߩ?~� |�i	K���a�1l�><�oۙ7:�TAK1���l��m�>	��wE��,R�A6����uؑC��kN��8 R˼f������א��;�>s�M�#��N��>߃�d}�|���ej���&>L�!v��/���	�8!L���ύ�1@�iY)G�c�-LB��]��q�'���P�ghxj��F��M/�6#+�4�V��g�i24��6gr�ƅ���9�"mΥ9��l��L�3�йd�ͱ��h�tm�)��[R�04D�ϳM��Y�Oۣ}�?|RN��4�317�VR�<�� ����H����H**t:�
��6g�3'�_��l��9���B'ф锔��¢��w�͙R�9
s
X�GL��Ō)���YkK�)	s�͙^T��,r����G�cs..<2]��E���?��Jk��h�7Q� {�>%%� ��$�z����vN874�����oà���6����L���&����L��q��&!��W$��Ki���y<
�ɟ�5�s*nq�(��a=��/�����U�X�:X�u��޻�F�q1�'�;0����>ԅG/�����ߞ�Tח�-���H[���ؼ~�;[zY�hg`��g�dt$�L̨'������M�ҙ0 }:�B��#@q�hg%�w,�/����tő�H��<П�k�UK�����z�,r�;:n���f�D�}��1�����F����}��˧C����u��=�U��$�@�"����E�B'ŀ����%$o��	x���ӂ�[q��l�yX�fZ�Fr���K:��h�o�$ַF"9o�B|�+
��,�h��&kG<��ˊ��Q�Y�x��_4;7"~1j�֟`�8�Mg��Z��:f�	#�:{���C�����Iz�e6����O_���xV�H'��g�L��L?��I�zſߊ���p��k?w��_Ǝ��'GT��.���#*�� �Z�{K��_,~!Y3E��J�ԋ{g%U�x�/ x��<9��=y�Տz��țgP��ɚ��}�����./�f~�ܟ$����I��� �QhM�ZV�[?��<�&S�������W��-ܫ�����0b-�n��uMٗ43��AJP��S�4�-�:)�-�u��GF�S��n��Z���L�����k� '^>mo %��Οq�U�F�Է��fm`����t(q)��%1A���v��B\�=}����m<�E�5h
��\Dax�a ���b��k�v�sÚk��
�ż>��;
�=��ż��y.�QL����у1�c^P�޺e}��xS����d,Z�PƎ!,a��)�e=�_)pO�����:n�\��;�/������ I�3�K1�e��i'fr0c�C����A!vda�-W�:�3Z~'ٺ\�b��[$�����iQ�#>�����<�;��yE��_���K�;!��E7ץx� �Q���x �U��v�1�x!����<�,�����Fp{]C�P�e�_�{�
�+��W���A�d�[d��đ����`�����$>s� ��UBS�h�/��]���ֽ"ɏ��@���w<{�3W<
G_@G��f��q$\"��e �}X	�_���21��+v�y��ѳ2���b�)���6���W�ݞ^0g��
��u�خ���V
:	�IKe8lC�C�Y��.tZZ����<Wh�Pe����0nZ��k(tF���$� 8[h8�����\H�=�m���?]XN�dY�
S�qf��bD��-�)^��/ΧO[�h������c(��:m���i	��π�ǎsY�z�~���c��-^d�q�{��?�O8B����V,	聀+��!_��5�~k���,��]��ݟ���?g����#�+>\hu}���:����������P �7jy&>��|�'��������)��s�.�9�,���kn+? ��]�����^�7���i������!���sAG�:��B�s
Z]����ÕVq%�;���qes��c���s�~�,�@U�@��:H'Iė�t���J\�W�(��6�&��aP�����Eot_)rg�#�	�Oc���sa�h#�'���3!��d��Y�$�W��E��.�'��9Rrx0��[#��2�]�I	9E�S�P�(]\�O��l߆O���T>c*:#����_� ͯ�{�;�f�O���J��s#��nh�����G�({6�3�l@<�A���@1���p��v��݀ur�\>���E����eB����-�+�p�w��\�1܁q��Ee�I����БC1>E=���ڏ�<I�$���q�ŷA�o��>��	��7�n�+{���'{�W�6�7���
�f���F���z��
�j���r�ǜ��`/��`�
x;�{�j���H�&���
�Z!�i�Z�K���B�x�'v	ػ{�9���Ga\��h!�վt �AV"�M$��6���~T��}�`���!؏��*�qQ� �{�^)�{�~H�{�`�{�`?�a���!�������v�`�v�`� {�`o��`o{�`o{�`o�v���݂�쭂�	�ł��q�Wz{=��բ�,ث���T�=K���]*�˰�
�K���	v���1�� �QB;�w	x\��/�W��^���J�.�a����=L�t|Y�>wt���_����n�[4��oq[$�����)h{�)�E���l8o�A_ҽ3�F��"��j@i�r���6T���hC]��F.�ӽ��9�%�+: Y?
���~N���RD��B� 2"=�H.b�9q3���F��w�����i$gD�#�;_Ļ����Y�K~O#R	-jG!���O�4b�m�m?�	G�b��X�����k�Cl���-��L"��w�>Q�}��ք!���[ �Z]�G�!��W��#Ɗ�F��4��63������91Y�I0��FL����#��!f���=���0o#� 1}�e���bV��1��=�0@��h0.Ĕ"F+`rS��,sb�S,`̈�EL���1��a�ALY`�i�)g���VaD�M�k���L6�&��c�����_���V���/�%�-��J1���N��!�
1��b����x��ǣk)���A�il���������#�otn����z��+Nw�@�]�lޘ�G��5�N(��l��x��~]���Rˎ��2z��9cy�w
�u�t�C������ ����_��2MM�w�R�2�	���G`��L�l4�r��_�r<��,�S\6�(x�6$�i�Ņ�:�x����#��i�>e4�GNA��3t
QQ��5�tL�4�P���h"ػ��{�ʖ��zԿ�!�O�Y�%ý��9s� �z
�T�/_��uɷ���x42�?�ր=k�>ʖ���'����b `��o�ќ�����9{��L�۴/nW��W/;g>�}�-jă{'`�u��?����x��[� �W-�AH(��;���{�l�8�T�d�<���yb4=���Ӄ��O�3=�|�BU�/���Í��3��n/P��F��EW?�h
^���1��0��oV M0��o{�G�D����<	Ԇ�H��~rW?��}�/��F���G䦌�m��kQ�� <'����=�d�p���+�S��haO����h�`B6�)<�������#�a��,��b��L�N<�4.�od����<�x�����t&���8#����:Rv+Px��a�f'Ow��S��%�r�x,�p��P�1�zQ(����/��se��e�u�㣃��+�v>�u��X��T��{����~&~��Wb�U��k�Y��_��[D���(�IG<�k҇j�k������x��h�_�#��x�N/ۭz�az���3�=���ﬣ�+F7hĭ5@��n�0 j[	/�#�jpyt���	�'A����nB���6���_���� �c"�'ĭ�8���X�u)(�s�aH�J������W�%�'@���������C\{�GMd : �?�>��1�>�1�5^j:*��g�&
�x�;j�Wy0���cvyQ����D�|�@@�k+�.?��U2a�W��-���\WI��ޮ8��}��/�ȣn[�wĽTd� �N�����8�豷9��bwD����QV�T:��A|g+����|~t�CW��*�'pؠ0uˆ�⿟��?4�s����_2���~�ӽҺ����x5�Q/nq�/�?S	�t�ǋ���?d�bqUxஂ�OX��L�%�G���$;[��l��w���9�^�(���׎r��6r�o/����sl<{�5��7�ex���ݏ���C{�eR��u�>ةk�C�Ͻ�:��4	��	��Bv����a��K��}�m���~)����!:��Q� b�x���#�B+����W�g�ZG�����@�e���Ш�8��hh\�׵!�WB�V��oh�Ă~p��]t����B���Rg,�z���h=���{o��l������e����Q��:�ee���w7ڣϮ~��j��@&UQ�7`Ɵ��K���ǜ}��yr�9��9�&&��}��q�7ϡ#�'�Y?��Y߉�Wa�X�'���F�k���1��ⓞ�#0[�3��1���H>�!F�O�����A���qa�*sF����qCU$�C\��� �z0�uW��+��A�=i���<^��mXq�f�`��� ��=�h��AF�?���n�Q���I�u���n���y�s��WE��|��d�Kz��>����9�|�q-�Ǐ&��ӌġ�0o~z"�"���l�@�SԲy�����\�4���{��D����O��=�Vr�O���,�ן���BA.
r�Pe�D��������S�/�����辑P���#M�dˈ�3�8��w��#�kb�X��b���{�q�����J1�^���k�[����a�s��:]7�����o�7N���zW\k�d*<��D!=��m��C+�uW�T��0�_x�g`J��r0BB�D�S�FL�αߌș��Q܄?�/���~��5A�Z�vt8�p` `���E�ot+�#����ڿ�̰����/'3�1�S��9��DfD���i�Ȝ��;2g��%3��2g��"sV�2�Ĕ����+~��A��(�E�ԭ��ē��A �.�n��> ``��� Q 1 ��'3�#C��'hJ�'hJ�'hZ�'hf O�\<A�x�f9��z�	���4ۀ'hz�'hvO����9h�B\��W�&�f��96�x�~law��a#�o<�vWQ7��7�|�g�7�~�dN<7Q�}�[o--���Ȑ�W?<�khǧ�؎�@�����#��G`%���bn��ַ�s�װ��
gc3Z0���پ���8!z�f�B�P���1�y_��uk���`u�{:��z�h9^nBV�-��e���v�A|�	���#J��6��l�?W����ѝZ0��<*��O�gae��s5����~>�=DT���Q\�]
i�����'�k�f��0w*^߉+R��!c;�z���{Z���}���O�P���#߯�����߆��z��ޓ�H�י�_����2�v�X�_������eq��X��)�_u�}���������B���u ���JJ�*�^K�w<������/���_F�~��ײ����Ay�����?��0{�������v�߃���?��$\�˄+�cD�[�>�_�V��+/�����ċ���n����Ǿd7EN��&U�l�6�>xnz�܇�/�Ō���{�AB U�OT�5�nR��d �\�|���^q�����B�U<R?5�mh�Z�kp�{�;Fe�F�3,���D�"2��'VW��e�.d�"ɕ͇@��3�ͺ���cw�m1]�?�7��X;��`b�}��j`�����*v����gv�Η�A|��5��K[FĐ�d����
c���և,��+L\sV,�7��a��Қe�;C��˨�5�D�3�`Nqg$W|R�S��aO��r�V�J�i䌨�)���ݖ�>IŰD��N�\�K�'���I�?�aғ��'=2���2p?�P���;�b�s��o��)�����w�����ϗkl~��ɥq��$���_��E�%�_���+���e�s^9�2�~��;��AT��ş�²l�B�t�66��������n�����'v��B��'jL�gωե���(��}u)Gw�1՗Q�ZvZ��/��ρT��{#0b��������7wc5�C��_!G��h�SX.���PB�ե��l�\VP.=u)�,��(�^���N�(�}�u�d��2�eO�Ȟ�V�!6�����Y���@SxH1��<�!� $��#[�9��9�m���dG��Q3��$܍����m�t��m$lԘ��U	G�|��7:�x��%�U�)���Os0lQA~�f��v��V┬�3Ȓp7i�����׻���^����4�&I�}���n�$��N�1��R�_��1Ւ�`Iz�n&I�y���$��闔fL�҆`I�p7���HRb��?�e/Ìz&8�����]L.��O�b�0����@a��Lp�U���bΈ\gݝ#���K7d�5��g��K�?|G+���<��ɣ�ß�n��n��z�~�����o�O@���/�W@� �YD?D���N�@�hs>�޲��=w�-T������F� ����s[���v��;�G!�T��=��M�3
~�~π_X8� 3��`�gC��x��xn
�OC��5��Y�i�䫎8ׇ�h� ;��:[�0K���h{��,;H���������5�.^Nخ��n���ik64
�����	�хH��vP�����>��.��I���^�9
������/S�+)GO]J'˱�Nڅ�w�g^V����
��#�Q���k)�V�A�q*˱�_Lؖ��6����c[]J;�q���_�=���<O�y�W�H_ʲ���o�7�rh���"?7ǲn��{=�R�Y�E�us]�v���ؓ����;�
j�����_���g=Ĳ�eY�O9��)�!_��|6yTץԳ���&��ץ4��3(��NYr�ʭ��tgO����S�u���Qp&f�<����B �
?�ݸ��y�֥�3R��JF�k�HJ%�ѷl�I\Y�HѾD�xcـ��FJ���Z���"e�G
^
Awdy�Gk]U1�e����VLX����$C���/"�xY ��dM!�x?Y<#k���������Md�>���Q�)��&V��J&�V6�O֟�H���qGu��?���6�$)i6\�k|i�[�j�{�Y�+5o%�R��	�*y)�S��B6����!�%�v~
![�eB����l=��![�����!�!�!~?!{X�o�f3�Bb=@ֱ��'H�"����L&�$)3�*�ͱY�K-�w���o���Xܸ��RҴS�Bg�u�5����F���� �����r꠱�
�Tط��5�Q\�i�V��6.oܸb���[��>�5��'0�/�
��ÿ@�&��/���A>Q�kh�x/���n���vK�S%��叉�&���_7�h��G>ݰ��m�����S`<�\����$ܵ��]G��g�|$�1�|��_)���O�x��1���?^8_�#�O�Ur\�,����+�W�f`�9��Ng4��~�,���dqƫ�_#������7:��S���u��6~X_��}��`��O���sZ�N�]5.0�����+���)F\([��1�=�������ȅ(<�6��G������JƿA/�t�/|�*BwݲC�&�8�f}'v�b��4���K7�/��A�=Ȇ�u�� +$Ձ6�_�����{��A���C�L>��Tܟ��O�Lw�-����g��W!ޓA'Wfg�!�2`�s���k�V�N�QB!]{+ښ�3.]��эn��3��ḿ�ٚm^/��C�t#_��Q���I�??�J^������a�y�� �x��L+�@��9 Pt����&W�a����͸8����' �
�N��uH޷0�����_0"R�M�v�E���^��(Y]���}��5�f���c�s+�}�ç	�(�|��FB7�z��p+��Q�&ڧUkٶۘ�}�x*�S6���3��Np'���7~�Q�����Ӕ�kJ,*[�?�O�)�����Oe�/R�K���#R�r�jqED��I�c,�%�����.�i+�s�G� ��m��)��Ů�[�x8Q\�G*h�AR�ͧl��*��
~|~�g�2���6�
#��+;�1Pж/����w�Q����l{�Y�;�)\N��q�چ�D�ِ�VoH ����&�!�ΧH����I����ԵDM�����'����
��b!၄8}�l��A��^��[V���gh~%�b�Or�Ն�J]�܏	]��4y�	og�o��g�Q+�So�ɦ��#�_��8:C�߃�w��[��d!�.}������O�un�P�/;�{Aw��?\ a3�������h 4�[�cXY�V��U��~�3��_�9�$ew(0�AA��S��B�E����Ӌ9��~w<��	ZN9[);O`Z�!A�0�b���Q0A�DPZ`��{}sH$hո�z�	$��Qve�i]�1�N�_���0����B���/�p;�#]�Rz��S>�}	ZFʧ{�#��'cG򑀘>B�w�/&]��B$�:���G_���u)���YD�|FvS`��^���.La6#y00�-��$�~>�2����+���7 ��a�T@�QIh�u)�Q��Q��Q�!�A�[>��g*����`s��Y�]��u�6��:�l����l�Y,!w1�aB�g��-��Y��HC�9�򠰙n&��ش�i3�l���/�7v^�V���_�N�[T�6��Aw-X� P��9��/������،b-�ׁn�CL��� `��G;�tv���Y$) ��):%-����n|?g�p)����B��o��k�Ȑ����h��'i�@Cƙ���(_��&,G�ͱ!�0�@�isl�ϵ�H
��8r���|:#4BU&�r�,��� ^�ɪ�З�\d��%\��B��lBB��� r]2f�I���A������aq���<�dL�#iS��7��z����x�gs�r��p}��Q��<�YNy��?#e�ŷ����t�/r�l$'Nze�e���դ�\;z�8s� �y6
�.�A-k���T�-����J��n�sY��n�� V����3�+��h�ZB3��t�mC@�L�PK��`��y`�� �L���\�_�W���pl���b����VYP�fm��q��(�#	\��фu�A�LJAJrml�Τ"�M��� +q��ږ���L�*/ćp}��>n~K�k��8�Y�:m�8���t�r|�:�9�x���4R�L[	
h�cM���zV[t?05.�Y*�	!2l�e%6GJa�������������-ip\EXT㧮�3Gʚl[˾�t4����t'���q&���qdۆS8��=��Mc�X���������B+�R���`�(��`l�3'H�z�Uƨ1$p��׎���Y>�L��3�V_����� Z�(�U�o�׏��41���$�/_j+qm��ԗ㝱���=��؅�H�+���
?�T�h��H|�-�;��vtD~Q6}���"_>�Ƌ���(='�0����(�L���#���)�H�w3˻������ȟ����7�ڋJ������Ekr
J�q���S��]��#�"[�b�;��x�.M�)
P��?�+���]	��`�����@#ne��{7�K��6��[��|s����u��8.tBz����� ZQ�Ƴ�x˅: j�����BȨ���~���7�~���7�~���7�~�S���<�G���Q��	��H��+�>�ׯ7�
a=����7����?���W�;��� �O���3^I>�ߔ�D�k�հ�)kA�)t�:}��ﯞ�d�q��:m���p|ʨd*��)`:m�-�JK**,q���s�v�NΈL��҉Hݐ��f-(��*��Y
y�o���R|r<D\�~�&���������"�����Q��l�?<lóqK�l��k��Q-X��s�w ϋ�޵��-�n� ,Q����8���$:_�F��i��t��o�Ϗ��}K�w��Sq)��R�?A��ŧp�r\_�軜�R��8�dy�Q�!�%o��>K�u�s�%]1�ƻ3b�'��"X�������/A��^�w'^����9��h�+`A=��=6��ԃ���������Y�w;d\�'ԟ�=�ҫzL�/_������B�,~��t����AH�_q��;0 �c�V 8���`��/i'��	���_2�?O���G����	��䯝�?��-�W��uB�v�Ϙ�_�e�Փ��'�/�Ŀt��I��'�Ŀq��I��&��L��=��$����3s�_�$��I����[&�_=��$�͓�{&�?����L�_<��$�}��K�&��$�ѩ��'���u����&�/�rj������L�_qj��i���N����>���εp�$��_`�<Y`H8p�����z�#=�?|����?���s��?��i���,u:�7�$6tK��H��Ker�R��h&%�,B��
���#��ͺ��M�f4��`�6�`���$0��� ��U`��f�!PÇ�<	f�"�� ��h��;�(0��0��LSf��`�3���\	�j��(��t��E7��`��lEw4Ѓ�`v#�^t�j0�n0���q9�3̳%�n0�莃� �`��T��h�:�U��f�w���wv��X�_���w���,}Q���R�/�,��R�g})�+�T�K���R�oQ�Ct����X~�e���1���X��ʄz+�[&���^��z�%H&Gdd�_o��+Pl/�L���e���k�j�Z $[�� � � � - m  �.�n��> ``����E D� H �� Z �  `5������������&���}����u|y�i������&K��Q�:<_�������	f�i��Y�)L�~�`�̎Z:}2@%@[�~�n!��I����ՅV����-���[�˶͌����>;6�������\�S���Dma�ԅ�z63y�
2�
3��-��3�0Y�����Z�)����x������L.J��:o�}���XD����.�ʨh�Aل8��L&{639�o3���~��#jX�3�+p�p�����P �p��;��\��8��.�V��p� \!�Jw0 ��J�e9Fp�7�p���UD9�d�[���A���>�C��k0��
�� �X �H��p T4<�	���5�I�؍����v�F��� ] ��	0�m�x  L W ,���� �
�	�00���>�R � `���;�S`v�q��� � � � � � � �� �x�(���-!�\ %� ��(x�`�[ ��8���q6ԝ��PpS�o���ފ
l9.�B� ��#��\�G/2����u̽Ԇ_�2T���aG�r�6�珤�Զ��+�-)�+ܒb[ᕶ�� 8W��1OM��1\���$g�maQi"�p���\��`s�
Fb�8������9�D�bnN��g'���r�31�t2l6\YY��p���W`x�4�;ә{�����\��ЙE��SI��`[��"?φ��*Jw8�nvbN~{V�/�P�[�
	�7�#��SK�uP*�-��d��H{Y��iE_9�9@W1$�a2E��yy���Lj�)�+����+;���g&&ʉф�B����q�h��$-��D��CW~aޢ|G��C����|"���$�����N���߼';=�i��2��G0)�yK�
���΂e�� #�՜<?>'���O���<�$���3�}�����J�؜�$�2x"<��i��8�KA������ǘ��">	čn3Y%Plj��uy�Kh`���D-)��e/��8��	z�X�Z�M՜P��EB[��w.*r�:K֬�Bb]�J�+�c����
s
�wbaFjt#�E����6���䛓7:���#�;�[�r��|}� �>���,��2l���v6y[��N����V���_r���9���U#X���pB/��R
rp�5hu���о�s� �qڸ��+&o�I��¼��L�J)���~ǅ��A!��%�Mt�s�***�ӧ���{�šmD���~���ӆ
n)�����b?�8+س�ٗ_�bW๙S�[������8-V���T�&͓�I륭R��mi����$�d1�8�Rf�-�e�n�������Ȧ�ϒ_*O���;���G�Oȟ��!W~X���K�w�䡊�ي��+.V�:�B����kk���m�;w+��xD��Y�N���w��)�T|��I�����<[�X�\y��
�j͍��S�N�{�Úh���X��ڴ��}�f�s�W��k{��j-	��V$�HX�w���SR��p�!ǰ�Pc���a��;�	C��l��x���x��q����3M�&��bZf�1�b���5��%�u��3�1���`�<�u�M����۲Od�d�r��E�~�;�������K�9��R�,u�z��j�]��Z��M��3M��G�����u��d}��J߬�An�2�1��l���E�k��+��{���O�a�i��L��,S�9޼�,7�K̙�ͫ���}@�Of��t�J��9��r�Y�TZ(�h�-}W��tH-sɚdͲ�Y��M�.��="߫P|�?��S��Z�ڬ�TP%�?V�^#ׄ�f����Yw�^��B�Toח�������RRa8�p��԰�x��a�p�1���QlҘ֙�2�k~��m��3k%��$i�4[���G��t�L"[-���ˊdO=�ʾ��.����O�E
� جp+�)R�E��%���~ſ��s��+��Be�r�V���{�	e��B�\���\����+4a�Ou9�?5t�����^!R·���f�N��*ToR+6.@:Ws\-[eu�Ge�=#{A�Ov@�-��C���'ٍ�6�y�%���e��K�M�]���"�Uu�*D=WmVߠ~X}R-�\�Y�qhn�ܡ�_�KsL3]{�6^+�&k��z��M�_�O���o���5v�R��4S��N�& ͖ۡJߐz�Ӡ}��.�m��-{W���Z�l�\����*����ԧ
�r��"�Z��y��E�k�C*�z�z��A��zX����j*4wi��4k����D��'M�v�v��l�Bm���?j��Ok_Ծ��iC�&H�	�	�	�&�j�LhLhNhIhK�H�$t%t'�$�%�	�	�	�.B���It�:�N��謺]�n�ή+֕��uպz]��Yעk�u�<�.]��Gק�u��a���G�c�}�^���-z�>C��_2X�/9��������� �o��������'�ن���a!�K�@[op@���k�q�I��,�ƹ���F�q�q�q��:c���x����g�c�C��/�	�4�i���8�̔`Zd2�_7��s��T��|.��rU��Du������U��SԷ�k�O���T�P�N��ܠ����o4�i��K��w�M�-᱄c	�����u����t�Ɇ�����󁶕�j��c�o�KMy����'M/�v��4��>2����5#1�0��/͑���@/��d2Y�l��Xv;� ��<���;)��_"_$_"ϕ�(���E���G�O�4�%�{c߽NQ=[�b��[٣�Q9Mu�j�j��jU��Z�v�˪7T���Q�5gi^�|���yڋ��i��
�6m��Kۭ�H˓�k�QBdBTBLBlB\B<Ȓ2��`I�B������:!/� �8�4�,�2�:�>�!��$�5��d�3� IYo�Q��!��Q�"u�$kq��$m]2�[�[���$�LWI2נk"�kN��u����ꎒ��N��E�I����I�g�f�W��$���Z��&�v��v�.�Gߥ?�?��������a�	��a�2DbC�a�Ai�.7d�3l�>�m�fxƀ�/��11��0h��n��g�̘`L��3K��:c#H���/�?4~i6�4�m:�4��dJ2e�ضƴ��4m6�nr�M��0=������=S����L?�D�i�3���(s�Yg6���W��3皋�7�qp������~�������Z�$τ���y��]���C��<D1M1��0�*�`|�z�O�&�U��9�ՠj��&�~�+34�5�0��]�O͍	uP�C	f�+�՝ܷ���FL��*%_3�m7˸����g�i&��S�)�^f.1��}'�kDK/����/Zv�l���u�5��0�����-�[d�A��Cv'�����������F��-������)�[~��O�A�yt��^�_�:�ZiR.}ũ�Uy��]9��X�����<�o�vV�/�ե��tW�l �-�gu;t��>����}�]�������T[�@]��H�i��+�}PG�M���17�4�0�6�m��|�Yc^u�e�ޜo��\f��|��~�_̭�g�/�{̸5F	<8K:4�ˤWHݠ�m�>,��H�#�xp��Rv��?B�c�R^)��R? U~�B��P�T,W���K=�Aw�n��P���U�����ϡ�΀~�R�\o֧�3aTs��v��N��I����o�@߫�k����>�jX�Y!�U��&����!Ï�9�'Wo=�Qc�q�q����}i��៍!��L�/�-մؔ	p���t���Y�����������n��M_�~2��d�A�S��A�+�����;̻�o���?7�O��t�3S�q�������S������K�H?�~+�E.�zK�l��@���[�'�_@[�+;�od?�����@�� zs����j��Vy-H�C��oBOk���4�7���c�1����s��4�k�@k�B�o7���%�Biˡ%cY��ZLm�v(�.�t�.�A(�!z�m5�Ӡi�4l:a��"s�9�e�6ǘc�3j���R�Ҭ��bN6[A�2@���+ͫ�yf�� � ��d��\i�6ך���Fs�p��$���n�0�2{̝�.�A�������Gͼy �;d6�0�v+�0*I#���(i�4F+� ���an��j�i��*͐f���� Oj�z(��(��\Z)��ւ,7H�M�f�v�r[�m�v��w���S�%=(���M���@^: xXzf:"Y�,R%��5u9_&�֠���E�,��x�!˂��J�O�dv��b��RY���K��fH��q4j��S�����#��񨌇^sP6$���qr�<B)��GC+�������r)�<�� �ȓ�Vy�<C�%ϖ�����A[ /��W����J�mk����6B��,�.o���^�.���#�w�ʻ�`<��ɏ�y��ʇ�àWs
�"B��RD+b�������m+Zи-�d�U���Pd)�+�y
��@Q�p*Je�rE��ZQ�`����f�v�Zm�vE�b�£�Tt)*��=�O�)�*x�c*�Ê
N)RF(#�Q�he�2V)QƁ.?_)U*�Z��-�d�U��}��+���yJ;h���ϖ*˔��Je5h���e��	Ɣ��e��z��.�G٩�R��h-�0�9���A蟇a���D�U�*J��QŪ$�8U�j�J�RB�mPYTɠ˧�2TY�?�T�V���y��RU��\U��VՂԠjT5��AjQ���T��.��O]���n� {T��>�Q���nH5�:���"u�:R��V��\Q��Sǫ童j�Z�6�-�d�U���Pg���+ի�yj��@]�v�K�e�ru��Z]��]�QݤnVoW��[�m�vu�z�ڣ�Tw���Շ�=�^u����W��C���Ps�&B���Dkb4��&N����j��Ơ�h�5VM�&C����0σ�l��X�Ԕj�4�JM��VSZl��	��5-�VM��0���8ޥ9�����hz5}��^3��i�5'4�V���Fj����m�V���Y�|�tF�֠���ȪM�fh���ڕ���<�f#�Z��T[�-�Vj����zm���'����m+����.�Yu��y��C�m��O{���A�@O�AZh4��D�.�%m4����HW�Nj'��Izi9i����6�v����6�Pw���EZ�!�S�HS ]u��U�Q��ƒ�OZ���Vi�i��f�V��j'�I:l9i����6�&��t�6�fw�>�E�!�i�H� �v�4[�Q��ƒ~O��t\i�i��f���G�n1i�e��V���@:o3i����v���I�o7i�������P�$=8�4�8҅����Xi����+�y�%�N���JC���Poh04���l�nh�Q���n耱�c�4t�aL�1��@���I�'�Qd�0F����c�Q�u<��R�Ҩ��:�՘�p�1f]�A׶��F'h�e0;���X���� �w��ٸ��Vc����a�3�N�3������k�3���q�8��	�E0�G¸m���=�O�Ҥ5LS��jJM0˔mZiZ=fܯݰ�T0���
�?`���Դc���A� ����Ǝ�#c�}�����{@�3Ε^(�=�*���+����Hs��J��A��5��e���O�ǀ�'�!��8�Q�x���0*����ǫs'�k;��Z*�ǥa�`t遑��QeF�Mb`$��QD#�F�l9�0j�Q�E#�-0Jt���=02�0*�D�IHhEBK��a���rZ�Y�������G��~2�?�����`�������)�J{U%W�{G��C@#���	1-?��"�@�'��}�/����Q4U�}W�����Q�%��-�৉8.�	�zx�}6$���0���υp�'7b^�N�������rYtgb	���p��i�
z��0 a�t[�3�[D���3�NOݺ��3�^ō�͋yw;K���d��BzO�GL	ԝ�˅��6*�&��S(�Wr�Z�];�'� ?�`+ ��=ݙ<�nK.�=7pk��ȩ���I��;�[��!"��� L��9�q�tWn���0��a����	ܚ"��q��f.�B��+at�2���8�f0�re��&�*L(I�P�0��>�(U�;��Ï	r�ZÅ\�)�t��3��mjf�PS��:������,�F��pQ�_$��Ű�`� 9�����o�ӝ��G�#���*�X�D��Xt���s�)N>�}6�m�v�V"��[$u��%�0��9��q\
�BN��
&�o˕P�`�J��V���A��o�~?����J�{�m\)�s	��r��e�p�i���qBjŔz.��Ơ��Ϛ4~���=jL��53xVt���J�+�Iߝ�.
��D�o8��A��3��E|���LTc�����鯏׾���9Ю�p���.���o���.�\�6�O=�c%Xv���T��}!)Lh�w:�*E$���_�7�p����K�/��[N��B��=�^�ʡ��^m��I(L�_�|�N��$R�A(�iΘ:/��A��2��FQ������k�[(|wP�C�ɥ�8~Q�kkQ�Z_GX��W��W�$�C��:�6�'������7I9Μ$�h�c&	���H��cm.�r�Z���\�8�-J�F�� �ĳ`q���0}3��T�Ó ��d�<L��m�����7j0h[}3�ƼJ����EߜD'\���'�|c�����k&����kߍ����H9%@ ��q:�:��fc
��ł�K5�ƃt(K�V1��ﵝq}y%�r����Y�;���,�-��
�5�bAZ�hls�.R�W���M* )�/��[�GJ���g�s�-"si��C&��o�Ҭ�:�݁cp�T��y$��@��Ú_H|I?�r�#]	�x��v���m�"!�%B�>n�xR�/���=|�,��#��쭙X׌'����J��'�OI|Nctm���1���E:!uw�+J��/3�t8�e6���l��#")s����X�M��4���_�5�tn���G;��W��f��s�>��y!io�˲�H�E�9$�9��EN����*��J��dJ6��̜9=NHc���/���-3�'3r���T̳��P�E�.�0_�;�%7O���L�$25�)'si~��Ms� �n��]�Du�H9Η����@�x��b��|(�Eh9��?�.	���/�©K��'���*m����A�݃1����rѓ�����?������S�`��ɶ/)��e%�Hv�#/Ǚ�q��,M�60g�����bp�����1�<�Y@*#���>5Nz�% �	<�5^8�, ���3&�9���=����g�Ya�q�E��VH��_��#���R�<�8�{�ȽW|^9�/7D�tM+/�
��
��z=��.ױ�%�Xc�>�����V�e����) [syTML�y��,1J��交��:�\�]�V��Q��kD�޽����B��qR����VtJ��Kn���}��A�őD��?���DQ�Sd���ݝ����V��z��%����P�dml��+U��~W|��[�v���J�W�M�[��ݛX�Л�~���]n�ι~H��k��v�Oʳ����~O�����iu�(����:p��+���ݽ�"OO���}�Q!�³w�~��5q1�W$.�*R����MtKw�O�T�.�4B������q�B�Cf��+�7�1]��w�b�~�,Q����c�̦x7�����Ք�Y����Q�F�Ϗ� \�{��}Ɵ���]r�7��五!pj��|���Js����1��m�x�m��� �-Ze�������!�u�!�}�Չ^A�a�Bk�[V}��#k�}�����3�sj�Z�{��cb�7��=�ޘ(�=T·~�z��P~,��]�Bb�x���Q��{3���4Vw��&H@�i����Ɲ�^��^sCLb�Ao��+�7��&hJ�&���I��W�(�,~�WqD���nb���d���:��Hh�;zJ���}w�4ͽX�2�t�xD�tME)��<ۋ��9ûۻ'��I����Ko�;͍"ő~��.2�ZD�M,/�.tGK��{�a�E�U��J,��Z�̺$oy�H����}ͻ�m16d֞SܿPO��_�n���׉��Hh ���ρ�_%F�o�g�.�RFn�,�mhq���.Y��[�+�4*�{��b~�ż䓀R�.��-X����B��M��˽z�U��Z��_��Dog�!E�Q�[uĩ���#�gjJ�'Q���V�$s��=Go��$���Dw��5(����{f@ò���\S�8�rj���/~NYk��0IIso�+��T}��n�+�s��H��$tA�X�ű�5�g����'CX'+$|��0a�鞊n���\i���Wm��}��Z�g�2����T�[��H®�j�7����wTyWA0�?�kn���b[�{�=%�R�e�Ի��Φʧի���`�yH>�/�y�W�8o�%��_�%x/����/�	;��8����8�A/�|Jo��ue��B�%b)�{ ��_�(�'�@$k~�D��NJ|Qlr��'�u�aֺ�8���籊�:���'���ޥ��{O��m`,f���g��F��5D��d>�'�7�2,� %Ϟ�zqD��^ê8�s���ډ�
�7�������w��X�s��~�}c����Uǝצ�o�e��ޟ�߅����e���B�Xn���
�\@	#���T]�B�_ay�,>���3� ��I��
�0�� �,t�e�5R��׽��ʝ�����$!�!��c����c�Q�q��0A8�G��pr�_����[h�"j����T}��Ks����Y8_����;�_*_�}T�K����r<�c�T$+R �(*t�N�(@Tb���z��y ��Z��m^��(�܉��(�WQՀ��������QW֋O[R/�Jjw3����n�=��w7�����ApZA�z
R�6PQ��� "��Rp[�mw�3��ܫ��bP���I�5���_L*[[syY[ȱ��>�{10��p&e�ٗ��Ù�0X�V�w�,$>] �}�Ota!k�����.y��
*
o��~�'c�b11�M>��&�IFj�����
���K��zr������G��ETQ���nj��9֠$B�z:sk�[J�*HC$}*��A�Ǣ��G>�9N���t�<�T|kݜ�v�ðs�{�ws�i�#���-����Ұ�?�zA��=�7�9U�9�0�W;�L��=��{��J�	�w_�A���9��m��y�"��iusf�B�H<�	W�`#~%���v����Zݵ�U�E��)*^���Z\*�:�i((ɱãQ�c�G�,��G�2�=<��؝�Q�����������������MAnO�� ww�� w_�� � h!�W*E�@�f���̦�,�X.���R�X.��r)|,������Q\�ťi��4}�f��R�(.�ťY��$N�z@��IK�~���������R��K��"Ͻ��Hk@��{V,��0,�����7��Ν^� G �~�x�R @)��A�g v�`�;1|
�����4�y 2���G�"�?Z�G����
�u#�h� �����`3�#�/b�y�I�Yg��gX�'=5�y�ٲ*��`!͢KY4���_}����cIX��.�m^9�6V��U\���,"Vq"��Q�~&���LI`Bp�R�����]�)��w����1e�g�xe���7O�8̾��,��@����q�->�0`�B�d���?�~��u��Ǝ]���A����K`��󐴦8di��ڨTwIL�������U1�|��N���q���V�����}Ҽ�n��GC���İ�� >�0�Q��~�"[+���E�;BI�����;�_��E�Ѧ�o���oc.8XA*�(���s�#K�OP���C��8;(SAE �A�
w��)�G���OAS�A�H#�WQ��I�c�$8�vj�GbP%(�����Ϭ��ca~����	tTE�0�k҄4�Ya�AѸD��D�A7��n	��l�Ff�2�͢,���4e+3�㾍��J ��¾(��kZ ������{�u���3����w~�9���W��[uoU�{�V=���r}1��;p��FM��)i�
�B�W�ql�ﾜ���0�my�@�惒�c��;��_ ޙH�	�A �j8q_i������38gnY�� �6s�� �9��G�'/"0mM9
��rʉl�-�M%9zHIQ�=D�'!k9|0U-��P��P�
^5���Z�ۿ�z�@��T�$���X%��W�ǫ�[ՋQA��NZ���yz���aޠ6<ݚ~�Z�),N?[�e���{ej+���Wފ�y+����wC��5�?&��z�~7#��'��G�e#��] �]ߞ~�^F�LmE�L�i*�gN(:1F��������8=��5S[���E^N7����Tz���hF���mjїwq�otq�|��d�$q�8I�,N��d~����%�#���X6��A��Si�`��Mv&#�s�O����E��Z��}�$�!jaK��+7�T?i����[���~0�I_��:{`��v���U�jiZ?�@ʤP�l��S.nۀo���\}FQrj)�D`��<^p�G�s��,K����1-&�et���ҳS��VJ;�zL��M���i��rDF?D���i��߉���Wa��o�G^�&���H\M��]��ǶI�yKb��/�B�����#�j���6��3�U3dˑS<&���.���W9�;A����P����'[��sƸ��#�GJ]�B!�d\���#}�X����H�z_$��"�@N7���@���� e�'�q��m�9>JN4�Q�ވh�e�m}�����D�O"D_�9�=�[#�h�h���"�I-��"D�*����}��G�m���{	�u�lA��#zf" �؉v��߷�/�m�����DS3bz5�ԭb:��c��Y���^��r)Ls�bz%�Ԓ���	S'bZw���֘����d�&����bʉ��,��T#������q���v�>uOL��C�~҂�r��k ���c:�O+L�v�:���U731��FNW��k����&Q��W�!|`v���&�?������K~j���{�B�yx��rB�1u�GlLE&�Sw7rT��GuF:G5�7P��-��sTSP�h�:Q�m��^�P��WkT�Q]���_8�'樮�p�R���m�|�n��Z��8���,�i���X��Ֆ�r�;r@j&�2A��kGב*��=H8OEv��g�@�Ă���D����)��lX�s��Q���Lq�8]��ڜ�Eb�����iI����f����P��tX�ϗ���f�����h9����g+:����^�1w"��Z��������B��%m���>|�A��@I���?���+�G�T��x��<�XTD�`�X��З7͓"�":e��tT��J�W8��H*?��4�6�f��Yh�56��zf4����0�*���ŭH7D�Υ"L;:��������Ӝ>�	֢���σ����< �
��H�ёУ#�#3��#�';Q�ғBU��W�=hӫ�T�5`��x�S��!.�ǘ|V#���P���@.-�3��v�����i sv"{K=Gz����;�A)�w���2�~�]�02�`d�GF�W��F?��-����� !ۨ�?�D�$�Ղ���K�&rнB031"�4��0�ٽ��4ƾ,�������\ӊ�V$C�}30�X��pE��=iE,�_����H��湧��Mh)NK!k�3�S� ����m��Cʞ�����R3����SW"|4�߲i5�RuW%m׉�
��yU �S?� ����P� uT�J|�gT;��b:1��q*×��1��q����h .��x�����>{�7�󞸦/'|�8UJ?D�!p�8�W�C.��r�Q�俐w��?G���	�� ��?������ͭ�{	֎S��|�*��Jb��b��ѕ��V/kѵH�����ƕ�B'��3��Urg�Hn��u�Z��$�!JN����L���V��}�*`�]���e�P��2`��ȿ@$+�����J�tSa��	m��w!>f�����M�j�SUh��$�N�.?r'�"P��S޴���]��x续t��b���	ޮ��z�©����<�;̳.ښy�8�nU��ͨ�<oDq���E�^I{�rή�XN��R�I�A@dj*fb�T�$U��P���n�\k�{ ���_��yP�BY���*���Ķ̎�t�-��N�6������Z��Y�!7�܏c��,�%2z���9�Px��Y�k�Eu�hע7��k��/�[�	�Ր�Ï���z7�V�(��{�PYn�l�Q����[��|8J��{k`!x���)���=�u󠣌6�v�X�X��`�oC�,����<�u���X��Y���>���0��7ݎy	E����C}��ۀy��}�ٜ]�L}�;������ҹ��"�+KަǪ���G/}�w�P���+$�?9Fv��j���6u�]o�[��N�ަN��m�x^;��[iSy�_�´� U��5:ޔ&o`2r,B�r<�z��C��^�N_ؽ��ҰH����M!Cˢ�h����=��8�V��1����c������������!��r�D�P�G粃�>[&��!η��G#<^cjM|w�~SZ���S8���ߌ�jT��C\�B&��1KAg��Υ���)d���8#틕e~�M �?3c����pΥϿ mYt���,z��D}>^r>���b�a+af��'s�VKb�G�d���?,����efY��ca��ndC\����j�_#�~��$d�oh�rv���$��^%m���"βI�[�q�O�uv��ot�Z>j�/;�[>��0�B�s���;L��7��μ��áK�(�z{}3�=��i�L���d���?�҈ML�ъK�g����>�淣����9�Z+����ҧ�ۏ�Cڏ����gR��o����ݥ��R;���
�,��D��/o�w��%�s�k��3dB{�\>!�>w�K>�*����}������翢�2O;������W[��o��.}�}�~�����ɺ-q�,k�[}�[���ڍ�R��8}�Bf��Q4�#	�$�:k�K����+���.A,�+���3Jk\�������=��V;+��e����y�ۈ:w�o/��:>.�t�W~Vn��e�4��!�9
Uyk7r�S���7쁏�rBB8�8,�լ�5 �gX��ŗ�U����)8����?��`͟�2�
�o_z��#�/>�~XJ�����a�iT�sR���:N���KoJ�����%�H��ڐ���_��C��ٗ��H���&��qm�~���d�2.N�g�߈���e�{Ɏ#c�8��S-�S\R����j�gќ�Bp_q���o�'��T"�1;'x������~��8�W�}��C����7@l��?j@�lQ/ĶК���=��Z�$���|P�F^:���;�5�_;�w��F�����5ǧ�"TzPՁ��*ԁ<	:PQ�\*��:�`���J�̃\����;�����@�=�7����}�j퀊ƫ�!͟'5����������A��s0��#����9������(�=��Qz�,�d�
ۮ��������^��W�r���	�X�>H\��G�䟞�%/�%��</و��r��r��;#c�	�ZΗHV��j���p�Rx6�(^ݙJ)\k����~���A��� ���'���(V�Xbyl�'*�����iOW�(����#d��Y	9��q�ňd�Ɓ2U��+<B��֑��h�Q$����Z���#+%ZydG�F���'	%��Ǻ�Tv�B�m���]���b&b2�"�!B
ZP��BcM�5-��j<�YqD��Y�Mrz��=Ɗ?�y#M��iae��l�d�Ho*pka%Z��v����R52]M,�3�2m��%�����K���)q�;�����N)(�q�Sn�$_�(�ۯx����n�QO'��ѓ!G5�����!��F��;6t(�9Jd5�n.��B������}kp�k��"/��z�:<�&�e��	Q�.NVlB�K�	��Wo�l�s$�2�� �%�7_�5���I��&q8 �̈́�l�I�
�K�q����+�;V�/~�G�D_���Sz-<�����|�:7[��g����gO�ط.V�(9�r�[#��a���M�j��Xv��XR��ޞ냣^��a=�}�2|��uϼ���&���܁�dV�V����j���fH�f[�F������]�-r�M���vv^ҟS�헾R��e�����Ql��^�����X��[���k$k��+�7� Q�cAzO�XD-��3u�uRoE:{H�7Y��~�F��C\���\�'W�l��@���z0��4v?La�i����~��	9p_�"���㠩���No�B����nX��G��x����`�rM��>�x	ֻ,�zi����o�m�q���ͼ��/���$İ�Q0P��a�W����m�2�se4���r��$0�I�l�=ΐ�1	���I��k8?n#~�d������u~��s���83��1c�f�]>n����_�9�/q�P΁���@�y�� ���<#2�Ye����Cm�N��L��s�ߦ͜Qٚ����浃E*����k�&��q�'��b�ƍ���[��G�Q'kp1��D��=poH��zR�в�P�sT����=�QB��F��y��7w�����
��I|�Ɲ���ɳ�NH�{�P��`��<I,3���$��
�e��\,M����~�B�tU�Y����M_K{�=�8��a[�=/��A�t�R�=��w�8<����j�v6KJ���� Cv���lP��v���] ���JZ�����xwo�[�Ƚ��"��@9Y�y�w� D��$P=�6�
k�u����DnC�R��S�JZ
��5="����U9	�kcz����~��.,S���^�פ�����U�b�0�4{��;o� o��a�d��@�s�-@᥽���2�d8�6���Q_�nZ�o$̰�7�"�pS�9j\y����"����5��eR�H�n��E՚�q���w�+щ��\&b
z��+����Xwv$�%e{����T�ɫ��/�s��t���NN$��P2�D�/g��qR��N�����yW�e����)��>�2�<���?�.?��$U�p�ZwV��\3�̠ݩ�He��8��Ne��N�'��ƜPt��W��! �,̈/4 e�H���x�A�=p9��u�ȃ)ꀜA\3
��{��v���J�k$�����jCNa yTnf�P�A�G���}`�Hd��4
NH��6H�\>c��x̿I�̜����;��~u�F�q�U��ݞ{��rau'�S��!�H�5��D�`�u���7����A�|#�mK��a�Z����&%Fy�+�PZ�5�<3*�s����m�"_�/�,�/2
C�vŞ{O��'h[��*q�.����� z����L]���/E:��f�~����Y)ͨD�`��O�g��|��%�W���%?�E����@4"�ߌ���mn޽������r/J�+Чe�|�*|_�O~�
t�a{*��b��D� �L�t�M�D�1cG��=�
[5�ZM^���c�Y6�3���"��|��^h��Ѭ��e���B�F�̗���}�u�̜
�r�l�V�w�[JhP���k�ۭ&�Fv0s=,G��I��螳K�0�=n;zUH��&%�]��s�n�I�y=�X��v�>U�js��5�2s
{�(W^C�*����Z��z��e�+`K�ДL�}�w
ħ�)k��B^��� ��5����I� ��W��JZ
ۭ�`;pv�����z7r�ϰH�ќ�!;�
�2kB���;�d�p�GX�x�]}��\���c�� ��~@.�7�-��g�z���������w�X2��*f��ƅ�e��:O��4�6Xͩ3�w<
ԋ��m<�o��?
?D�M��6 ��`Є�>�����
5k{`�+iNH&C�֫@�ə��x��ϲ��T`1��p_u>��F=F���R� � ��[�tkh��(y�}������B��Ch��9�Z]�xf��]	��HP$��X$d��v��oV�-���c��;W�`�z�Q�$8Е��ژ�fȟ����?�&U:���M6��9���R�znՐ��9y��}�5w¾�����}_~ψS����A�UE���ɿ;?�p��JW�]&���V�4GH�Z.�Ra��[�ixO*�&��Ҷ��c2膀�ɽ[	�����	��!�u��r�%�ej�6/�Bh��� *���WnK�g<�I�g�'q촱g��?�OI���o��=�1��.H��(�Dv��-�����:�(U�,��=��K�"���i�Kq���6i�FZ�s�o��b$��M��6,f�yn7w߬�\�W���y�Fml.4�B�J��<:�*��Y� ��P�0�l#����r� ~8�_��0;��ڀ�ҽQg�t����Ah��l��&'!R`�,�7(i��4�(p@��&X"<����ۋ����T�G#�=p�ۙ��M���!W�]���7�qZ�,Xa�ae�I��骮=�2�w
t�Ko&��Yl��6v�׶$н���;�_����]�a?hn�)i5��t����	�:�w Ȍ��K��@�F\��$WJȏ�#�[���\6_G�SX�N�}�s��(rL� ��6����(~�fMv� !� ��}
�_���mPb���_��ڃ��������U�p�0�5ɣ���Y@	N�]P<�0����l�����Dq���Ll'�< ƣ�T� �ɫ�W�}H`|<�s����*,��J���6���mE��t���}	K�h�LI�ǉ|�SfjT;%�;���@S6Y�A X��'_�����Mu)1�R�-��z�J ��Cwm������+�s�*��Ʈ@/�}�n�]�6j��t�)�t�\y>y���=���A��j��^C���pT��r^��c��\�����ݬ�c�&��J�[�fWH��k���}M�$��JSY�CO�AU�w��(�
WBJ��+ȟ
�R} 1}�t.�[�ַ~mJ|���5I|7`.�y�hYpb�:ɷP&SFASKT(o���Q�א5(Ő��3[I��/P�"XZ�j��=J���._��;Mb�c^����Ӏ&p��bX���!��u�>	)�L)�Pِ߄��b����  y�D���5�ax��1"k��q�Z��O������p�dƮwb�j<�|k�#��L /���U�(񣃾��m�zv��O/�	d��&�e'��I�׷z����5a�La��$H�X�����/����B�o�y�M�S�y2�*vm��1��)�eb��mޛZ�'rM�*פ�\�IR8ۘcl��q�����lyJ�U�S��sz37MՅ�<�oM-Nr-�_��h��7]��J�����FC����	�7p��!ߓ�F�i%� �#��o�XO����) ��&���M��]N~�X5�n@�Q��C��E�9U�n3'��>��s��xlS�Qd��"k_���ng�ai���h����.4{�T�����J�4߅_�ݪ�?ƣ�zq߅��.t8��X�B�T�%���;d���7x{:�I_j�N��l# �;�B\�
��A
<�Ǵ�"?��3�K�|:�ռ�ЯL�V��3R�P�:�f�!�LKV�M ��V��W#�&�Af1_w����� ����9�4��@IK��s��[̆�&]�EeZ�!!l����r{��*{fQf��oV��
�k�f��y�X�ʞZ������?!�*t�u�!�l���s4�q3�����7���S��	�h�i �Ğ�ޡÙAGQ [�OVFvV�S��\�2�7�����s�ۙԌ{�P�r��AL���}�"�ݎ����ި�zR�;X��vӏQs�N�wȀ�?��`/E��藌��VI�쭍�c5�zڃ#^��_S�&(&8"���	J	��oSF�".��E����.n�ō�/vf>C>�LB83_�=>����>LZ/�c􁵸.�ópس���#������@Ari����h�mZ�D����(�T�x�.��n2<I=nI�#�k�zM¼qMg>o 8.��m}���+P�Av�lvN�mW�>Ԡ9��!�bm 4t�Y���#B�~貵����I3Vw���8�osp�ȰX�h��Z�"Y��N�`�e��xφ�lx����� �g��,���� ����p+o]��l��e��-�m�Ј������
�#�Jog5�i�]�7<<��5(��Ǒn:�o����l����W���S��ǯ±������Zi
���H>��!`L�轮��}c}�KҤٛ�r���B1P*Y���T=��"��<�NK�B�����#�J�����ѸX� g.�.�޾��'�@�bſ Eu� H��'h5��Akau�֙�Co�g�u};O�����q��5)�+�K��Ä������ø�6j�B+"WIl8�Ixh� ﳚ���u�t�s3��)O����*�s���H���X�8X�#vt��;!�-��6��r�\Q��l߯ƹ?�H�)�h�G�
�ە�-_�)�@�	t$��lW#���}l:�-ؽ�Ahx�Q��W!��yг����W�r=�Wx�l�s��a�#Z�Quvk���(�K���>,f5�����&�S_������[�^��F�Z��X�������۰Rz��E�_���Ԣ'GU�?�Ѫ���{B�M '���d��D,e<j���@ly4U(���
V)��|4G����E�F��ܶ�?���n�w-�`����K�n1������d;��<6j�Pl7.&vkhA�#X�9{��!.Or�E��W:&p��B����.9}a�[֙u��t4�]r�������w��1+۽��!k��-��K��!��[>��/qد�	ڒ:68l�:�:ۅ�K9��zO"#���tt��d�| 'k�W���_Jܩ��ړi���Snq�f���}d�z'�!o�����|p` 9@�+3�E��RpR}�ل{�r�d�H��]le�\[ْ�*�P�E�hGx˭r��T�	����Y������Z��{d0��rM��8|��p����q@U�&� 5�����L���3a5"9�*-_OZ�|̙�2!��dX+�7��T��,����oE�m![���Ho�X�c���<�u�,�厯Uh�Zo���LZ�_�p9��}p2�~Gc�$�W@�T��܅g��dd���B{ɿqj��w��T���/��6y:��k@u�Y�� ^Bh 7@�Z�����q�4zN���E��|4vf���1xYZc^�_�U�oU�爫��R+Y�p��E>WҾ(��r��2��5fڅ���'鹑�wȋ{$n?\G���H��&%��&�{��؏�ߊ��u>;Qme�w��R�4��e�T�}�MJd��sL��-���F��}'
%DD�(i��1�?���Q5ҝ#�b��v�	n&�����Cʏ�p2N��$N$�A�k�=W�17����Ȧ�h���kR<��+�}�W�xf3s7��k�S����ǃx�9���xrse��!��p��O��y�X�"��'����a<`CƚO/�hl���b.������d���x��v����C��+*�>6Z%I4�?�4dK��s9�x��G�P-B�7і�,�=�7�ݏn�,����iA�?��v��@�Y7��X��b�,U���H\�!L�[�����9CݳJOhQ�V-:��Ȇ�su�96lά�ԜCVn����:yV��f��-(hۂ��|+��"�%��>�lS5��3�y����G��?�G�xj#D�o��0�Z��.�{yP^|O.h�0[b��M�_%�@A�08�vV��j����Co�|o�kx)��ɔ��[9��^�o�q�3���n&���	��q�Ŷ��{8(�ߺX����Il�\l����l&����:�~�4��5`�sv���B���Iҏ55�z��*�������ƕ�	o+�]��Q�-�t��=|w?CX��e?��w	^����l��J�X��������P�b�ERB��<3W&{�8�(��o�to�W"1��ՠ�ڥ�$��������#�U�/m���,΃��j�r�����F�ZZ��6��_��E�{�������o�o�!Oì��tߥ.#�fq;۔��H��hF��-x��O�wk�<��H4�n%?(]H�RQ��5�fW�im�b$�Gi�&*�S=ﯤ�{��L��4��eS�>B�Waq\�&��<V��ǒ��4��}v�B�}�Ѝ�%y+ �.����g�N��H�����g��wwI^0!�z����=��·ѡ%yI���W��}�k�b\���O1.��������=VQ��VDS���� 1R��$R��E�KX��̞�`��ƛ�j"��,&s�}.�1�u[��%��h]��eY��~�Z.��;f���!����XݻnY���?�r~,��]��qF�^�$����+�Fa���=)���O?�a$�_}����U��sMVs�F���y.��ȷ�hӼ�2������7�w��E����H�NX2e�FU|���̡I�e�9�1�?��R�c�;Ή�r���`�+���I���Rv�%,���E�Ͱ��|���S#���7�W���w���C�.�V$�k��q������M�7������l�'��	�OL�Eخ1~ٟ�������y{2�y��{�n�7>��Xy�k0	]���_�{��·��g^���O���NI��H�"��B�#t�.�w���z��}G�I��G��������;E��?E��>Xd�틷��r��[)k�2Y
G��u�$�>���]b���:�g�J�U�$뙹�.9~Z����>�tRW�u�N�E�zhn���)�ȞH^��-��v�zj�k�@o;�Pz�o�w�/����
T�kV�������!��з_��{y����d5#������=mz��������e�wPIN�ȝL�6ϝ�����y�^]�{��[b��������71HV`y4/��_�@�������K�{�.Ќֺ����A;C6�x�*F����ۚ�r_Tv�i�yTW���_l�X��
�U��j��Sy�p�;�������Jڰ��a�DEH���^��Y��]�>��!�C�@�0�۴��8h��b���rV�JĒ�h�ܓ)��x|����Sq8��A��g|�I;r����W"Rm�� ��X�K�kܦ������ЯǨ��WԼ�jѤI�|{���r��������\�䥤@l���.���.��όq;��p
��	`�ۙ�d%���I�4�R��sn�U:XDw��J����Fd��?Md�˵�����	�i�˿۫�,�b��طSKi7���EH�M���4���8�v�W{�$�aGKۮn߶K�)Z�TF�Ev�>H�
^�W(V�*KHx���@��?^lL�z��_�7EI�������(����������Mu�mԨ,�$��򤲑&)8�غ������T�G�S�❃���5��*��j��|�^n��}V���TI��g��Sz��F-�W#M�:9�#�������h�L�Y�e�����V��C�0���Qt0m>w�sr��!_������آ��&�7���ڶg]2�'z���.�e'��w�aI44���&G�ƻl��������˙��-Wt>��f�㎟����C�����l���pV�Y
���Ѿ�GS5�DRI[�.&H�vj�9���yH�� .�Wjh�V�y״s,J���S�/��\-�l{�{�U�@NY��[i�VgL!�s;���˹H����t��Xl�x�;Dj3ݯ��
�̍h%Dd\9֪�s�I�S�n�f�����ϻU
v;%Yw�u�蒎|*����\�c�f�A�{��&��Z0L��5��OF@���=��;��h8��f���I�]<��X��>x�<ɮ��	ݙs�����9'�?n[���J&Go�$�$/ח%KJ����mr��wi�T����ޏm��<%�����P5Z����l�i��𬧦ؚ���]�+��(�JCw5z���ማ�2���(&S���i�FDxH�&o_X`؏����bX]�#���`;#Q�R��'U%OC|%�_��i��4�q�"b����Ao������-~�Лp9n�R� ���h
@� ���Jed:}&������
l��	�Mh���	3TW�K�5���q>Fw���77ֽ}p�@�oX>$�((=u
Ҁڧ���y���)'P���L�`L��z(.��>���d/�������'���k�M��c�����:���S�{��UP)��r(t���>��׏!��Jd&=߽���S%�sU ��#<�CxH$�F^Mm\�����P��nX���_܀�������<t�Y8{Tz���t%��A�tt�S�4o�0I7`��(m�3b�� %sdH�z���)�9��F:� /9-�H�=��v���zI:ښ�����镗��NmS��I���SCL|��u:���~A(?��~�PVn�v^p���̀���;�j�t�tT�4��G�(;f#�ڜZ~��Nϰ7��<�ݫ(N�Hg��ojȓ�#�]�f��H˩H�Y��sHҚQ���������s�A�f�r~y�+�7"�s!�D�����B�\��2��j*Vm�z/�m&�Q'���<�Wam0d�JH�m�T�/���Y�:��(��*��ɐM��)����g����I��c|�z�ƣG�=e�o��ό"�ݖ ��]�a7%����zrX�Xw#�O����_�dV!�����V�8U�4��´��Zt=�|r������Y�������̣�{���U��T=3hV�%���HQ�2��)i��(��6C�ӯ#-��?�^`��s���G\G�@3z�U�F943M!��z�C��П����z�C�kcЃ}�Cwr�8����p�f� �A�q�F}*}���p�z-�C'h�������"��8�s��AУ��3���	Zšsh�51�u]ɡ���o��t�.�з8�8TG�^��w����^}W�B���[y�wy��x�=�nU��qh��]8�}�ǡ���	��^�>K�=/'�k�C�t����ǲ��Lпq�3�%C����Џ��a���8tEzAm���ZڟC��Љq���j��{9��8�(Ax��S84=�F�ϡ篎A��=ɡ�šo�ɗ(z��D�[��}��q�WӨ-�Os���Ϣ���7��z5���C5��w��x��
n~��&Ƞ�K��9��],"��)4K�S���3&/{��3���2�2,��7�d�Fc5�	� �
��փ���V����K���stCnG�j��V>l+J\Ty&^v ��r=�T���R���P�oם�v��[F����{��kǨ�/jni��c[_�Phu.��:��b��#�c2մu�7Α����M�o�ns+����er�<'�=םu�Q4��);=!�Q7ٟ$) ո���� �k�Y�+�~��6	��G�����No��� ��ZO ��G@�q�7��K�zJ�h�L�$���W��2��B�[H������ ��.X��<�E��H����,v�-�1ȩ���6:�VU�*z
}R+U�!
��#+��?e�l����9�vl���̾[6w�U��O@��$���n}h�W$k��A�7���-#��oG�b0��S�n�4��xo�$t]���30��h�%�1�?�n�Q١T�����c�=67�قg�A��gk{�o���ɗ��玖��c������Q$K���_��ڋ�� ~�릸��
�kQ���fa���T8� 9����SN]�%}���aSe����ү���o���x?m{N~��1���G؃���m�W(�F|� �;�1�����"��f��׵"@�����Y��v����k�C��
�9�҆`��P�������Z����f@(���VH�0�ê��j����TB��a��0��t���j���H-��3�J��$e5I�I�Z��DEc�tN/�,1О\��@��G�yڬ��#K����cv�&z�ڟQ�I��9>=%P����`�dd�*Xޱ,�0/Ǔƿ���svH��*�{���me�f��f=������l;h1W\��b�O���l��)���E�0��WoS"V�Y٢R	��-�����R��.�eb$�zo�h�g�9�"J����o�!<����,_�.��ZfCX�������L��@y��rp���{Ԥś�Acy�zd�<sj�`�TZ�C�kȴ���tܡ�Ϫ�&)i�1=��������*�3-|����pk��S��Ø/`���y4���O�J�o�AM�݌��0��M�5S�lA�N~�2��-���h�ZSfo׸I��3�c��&ɋk)��v�$#�!ї�,憾���ž�:�����K3�㼙h���C�"�Z��{�&�P
t�W��=E꣭-�D�[��ͮ��\���5k���<��z����v6��=݄�ڡ���q�.y����y��ϹN��o�/h�<P|��ς<Jh�����T|a�s@���|�s_o�j��^��[�	{��_��F�	��xo�X�~C�s3���R��+HL�Na��j%j����`�l��ޘm��"u�0Y�%���b��ջ��&���
�� Uk�u���*����{3�:�j�N�㝐j.��	��7 �m�e��}��ɞ$WV����ov���~�3I��/���t.,,\���`�(�ޟ�x޻���h��6:Ye�Я�ä��C��[ �~�ੇ��#�� O��.�|!�k_�$<TQ(�
5�Ow���|�y;d���k�p$�scT�B�J+\%Z��0V����ꁟ<;ੇ����g�j ~������VA��$
��lR�>��R9x$+-I�3B_���RT?��ó���Y��E���;�ϳ�<ϓ���g֟����*0�\a`��e���=OƟ��f�9A�c��*�)�};�A`�^g�d5���c�K6��g�t�1�Ac�1�yL6�4gQ�X�1?�<c��c<�ʍ�#��\�c�6��V�	�ߨ��Z�Gy̩����-�9����j��#7��2⑟��<r�|}C̓���-l���׫)�#�Z���gx�c�����A�������<fĤ��Q�7�[��I*w��tY���J���	Ȗ�M���a���I��rL����,��#����<P$?��'+�]*W�{R�T�;P��øM)O��;��<��l�a���sy�C�kx���F�-���������

�c����|���|d]E���-<L��x���O+��#��s�����
�s�r)g��G�#	�<�Ցg��<�FrY�atN���0���<�Ù<�����<��\r*�E��/�?�y?cX�����?��F@���!��a<�#��xy��:���<\��2���b�1\������0<���P���a�m<l��`N�� F�~��"�|e�[rS��9��a�dVF9T����b����K��<<ß�0.����~���1�$�a���W`���/`x���i<��<�	��<�ù��y�6)A�.�����tx��]/���NG=i�p���Y9��v��'i���^m��P¢�ɖ��IU����m}�Xm�*�kep�v���ٙw!;��� ��Y���+8��B��w�l���|G�ωR��e��������̹�����҇�H݈z�ٳ�����L.a�����6&���͓J�᥺�� �z'����a(��K����#��ru�- Ov�g~T=)՚xq���B7Cy<m�� ��#��K����>���t��r��O��mq�S-�o��yi��8�E���xnb�"��{A����tr�p����xv����/C1���T,]��B:�H]1Dٛb]q'�x�+���Cbݐ"��u%��8������/��2��֫=�^�=B��b=Ri��r��V�����m��������E�*�2s�l��N
� �
ʠQ3��@c��Ũ�d>�K��%yX%�A�%�ԏk�x "�r;�I��*���&�/�e���{--���	�ȮF�I8�>�5�3߃�J�y��]l3�Qk�Q��7	���7��<������ƅ���(Fŋ3�N���-,j���VcІc0���1-6���ιY��k5������.bHK8���U~�a�Ƴ���_&Y\�_bC����yq��F>x#�/}���EH�r�@��aDw0I0��!y'hx�D	�*�F�~�0sϲ��ܪ���hj�3>�ߌuk��|������8+�6~�\����u�lvb�l�#�E�0 �����뛉��$��͚��D�I�wO�10f��k���&�\L��r��&�6Ç-�&&���,�s�Lԕ�T��~ď�v��'�i��:��̣%�&�UvV�*��e�Y�W9�U�OG�����r`z�d�����;dۀ�o�zf��r�&�$���Y4�QB/���W��q�1|ޘUa�
�g;��^���wv᭰�{��Z#�j��]�����۟��=�w�k��eo����n[|::�9 �X�!(<�B7ٞ��������H0�b��k�n����bЦ�@��l��^����gP�j���\��ZE�� HY{�3�w�0�nw��ˡh���uϒ�RЍ�G����e������~�p!p�a:}33�����Y�$��6-�v%�4�͉h�?'<}�e�Cx���JH�0��E7;v26ZV���հ�5؃��d��A<륆mg;v�0XĎaq�.;�$4�� �>��:�V}#�9���n�	&0��}nk��4'�!����˙�(\ir�8" �ʪZ��H��}���Q�FE�ўU�f.�����q���Dʊ���"P���;�rϫ�=��(�6ۃ�J��y:hdp�2* @N�LА2���2��:\�U�~���]�]{�=(s���=/IU�I��їi5�\8QBH�K�#�N���=K��j@]�[�{ې�ѻ�={�@�����P��d�U}��M��}c��0�S1� :�����G���u����d���fl�������x�>���x�l�Kunv��sZ�-NC4��cqD�i_B/7/:`g�>�;��WD��N�&����@<�뫡�,��-2m�g��
�]b@�:�������c/9�)	�/�D���.k�3}�c�o��o��+5���!f\
 {G��k�y;2�G���ה���:�Yr7�!y����,�>~��=*����?�ۏ��G��O���6����m��?���va��7o�_;o�9����������4ok��g�ۋ{$����?>o�����������K�ݼ��x�;hY���Ѥ�w&�&mPK��r���~����]���w'*L�����B`�v�=�P��0������3vW�����_��{�MbqnƂ�N�+��Ns?�.	oU�3����aq�~}���):�E>�E�E[�-
��x95j��7��N���! ��ÿߛ� %�Y���;<g�����-�L�]�9���;�}bY�~'��ݱ�@p�7+�d�)<5�,>�X�Z|�q�N�,�z/Uĉ�Ya���������c=T�9���^ԷԴ�ɒ$V�o���x��Q��I�`�}�iAWڸ�C]�o��մu&]]��D>E��|��?��ŉ�6�
/�G ~Pt�t��)M(]��C�B�e
��2��Hx��J;x���Y����_��y|-H���n�v<�"@� �K`�Sd�=��$+>�Ax��y?����V�E��縁Ԟy�gQ�S���	�� �7}�g�3�������s3e-�/��û)��9F-;M�A�)>vC�y��ސ������H�ź?e��-�i���a��u�@2��/��*��K����5���l^��<k�DN�|�C��U�#��<*x���ׂn�23��6t���!2*@��7�q�O�?���O 0��Ɓ��x���B�����Ì��D]������)~��]�?�c%M(�-�W�ls�;{3@0Un/�i���úsHd��������x��]��?�5��ޗ7�	d=������cXNɯ���!<y/~s+8D�~s'f9�R�������](yӟ��5�S���b=N��Z�E�Q�UM�B/���꓅�S���9ɗ_Q�6)��)��
�y��d#L��N
N�p�=-tvl�>�.�e&����B����]+�� ���������-t��vm�h�|����V����W���a��p�����}A*W	͉81^�\��W�uT����5oz��S�������H&%
y�S�&J�!��א���)L��},��AoL�in��Få���\H. 8��$�9�C(O�;��-|�Z{p��nm@y�Լ$�N�97�^s���B��O;��]��;�sd��L�e���yG��/�s蛡j��4H'��D��]���C�`��@��Z:�������N�~W�X?��Ďp����Zݱ��q'���a�qY5��#��#
�!v��l�P�j���z?������wF���~��h�p?{�:q�1{�Z@������W�pB��J��
���Q�P��Xb��87}+XĒÊ�YrNS��x�o��U�ao.s|��O��|k�?��ގ�P�Z�_�R(���0���>îR���<�������q �үg�UP��6�G��g�&Z�;4�ڨ)V��88�'.����'�g�0[��9:���1�7:�m����"y��Z���2�9�-��x�P�RX%�XĀ�a�w+(e��Bwy��_��֟Ÿ�����d�۟�>
W,�5�x����q�o���O!��ᩪ��))'T�;�S*W@"��f���⽓�4����A-�|�c0�{��g���V����Z��X��1߈�6��k�a��%�Fj%k���{�.��;_��;Op�
��Z#<�W=�|�}�|t�2Yb��4z}�=c&�a���U��1H��tScX��ܐ=@�Y6�u��A�O��U[0����G(���h�����v� �D	���Z�<��y�[���X�f�]A�V7����d6}X�/�@<���<���%<��9O3<�UMox����tx��xV�B᯲RV��2�뀹t�hx�č�b$�%@�b ���Pv�j]�M+Eܦ'�9*�e9ʒ�m�Js��1Ln�	�AZc��m�<��5p[�\��Z6F�d�2p��4D�3�ú3���pj�o��t��)Ȩx�b��s�=�c��aGlp�������ӿ������a���$X�'Љ�sE_���oŇ�#
�;��d�++s�)D��hJ�
��l�2�+%����W`�#@��y"?��F��^>�S�1��H���c�>�
[�}Ć8���'����L�]� t�0gg�F�%�t��Y��й���J���
x������֩�i{�R~4�$_D�0�h�A�!>�Ա�[�]{�� A�-�NP)�ǙU���n)�%�G҄͞�l����.�ɂX��u�ŉ&W�3�G��>�ikD�� 䅌�2"oo�$fa�0��3vgUƈ;G�J5��{�9K��qҧ^*���-��B@l��i��l�̀�l�������؎�����T|��I𘀊H�� ��j�/)g��n��t³��G��*�Y�{SQb�[�@8v&d�������)=�_BJ*t:G�B���)0�o�O��/1E0�ɏa��-��9�臉x\
�		H<�F�7�����Qf��m=Զa�L(��i�BH�F�e���?r��A��$�?����zĬb����@ϨL������-(ֽ��"_��)�>����;�� WVx�PnH�)`w(��cD�� ����z�1*�ca`��f18� ������/�c��>$�Q��[C]�!o>����k&�4��Ŭ
��u�-�w9Y�=�^˿|����D��G��楛}5
�Ƭ��!�٫L�΀�:��g��˅x�@haO�)�h2O����C��3��og�e^.��3p���G��.��ȉ}������Q�a�=W焜��2<��ԱR�*2����kDeW�Z��],�D5jB�k�'U�NL������)xʳ�߭���D5ҕ�-P,�kP\_�w,
a��v	��GTd8}:��<)�xd�u�g�P^*P�8��چW-��9���wVgȨ�@�}wP�����A�_�
z��;�,�� �#����H��"!%���b�`"O�l�;:@F�X�O�2���UF�=���)�<{�l����b��ۭ��l�� ��/�U�����˿_�}x9b���Uu�D������Ȏ�24-�zjAO��WU��aU�
厜 _���
^���qhP���&t���Ӈ+8�Y�5+Rp�).ث�C��>����&�)��M��tג��M�J�V�7����ˆ��Y��l]�������e�7K�[��~��]*�Nt��yv���������5���jp��<j%v���`{����Pe �.~���+ �l]�]���������⼽!ڍ������:w�b��f��(�tĻ����FG��ƿE73-7�e����8�Z��.X�B���[�BX�nt�
����B}EY�3,�Bх��m/�_(��J��)8NY��f~U�^�Y��mpZ�{�-���&W-�5�tUe�h@m���t����[�̻� �<�����]��ʬ7&��!�#�A�D�h֖����,��v��-��������a[�#��~v��Ｔ!C:�����6ay���!]ʒ1�*��S���ɛ$��ݳ�:iMǽo��}3�wBޤK彿�儌)���5��~޼Fݥs5B.Q��L�����(���~�>�h~�xԥ������>˝O�s�R��E���u~�n�0��9U�������7
�|��.kÂ��Wk�?��(�-���W�X��Z�����%�k�g+9Ћ�������
^��Y��1�dx1(I6T�e�iE���MF��h��K{/�-�q�U*��,�`�ύ���JQ��lX�.8q`���n� ���
��#��"c��b�]��������\� �F@%(�`4���Cf`f � 	�	���\ �[�$m��(m����}[�ַ�m�"ޒ���B� �F�����B�|k����������y�/���;����{����k/L�ou�.�ŪXқ�r�w��^�4����*J�.���7M�3�5�D>��G��u��O*I��5���J� ز,@�@M	�R��t����R՛є��oI�̌���N�9�&�+�K��W��w�m���6Ea�rf��mW��|.	S��V�v�ڿ��S/]� 3^Y�w ��~2^bFkǩ��V`����� K���W��������Mم�Jo�ɖi}�?~��98/�`������ڌ�G�b�DR�H)tλ��٬<����.nM�X�s���`J��z-�j���}]�PM�b�V߷�K��-����lG�2n�5h=fS�,ʠ���<L?��T�{9.��p�:��w<�ẗ́�!w:`�u����	_�#��߬���p�jx�m(�u�Q�nu���p��4�2��譺!��knHP�O�d��2���v�(n7*���'�9�J�K�1R���`��8�Tÿ���V�ޫ��iٝ�Ȁ�AvΌq�E�Ec�ip���dTC�-��@Ǥ�O5�*�����d�ogq�JW��c�gG�
�C�
	�Jg���*3T&H]xXϬ�b��gRvY���Xig%�Yh��=&I����o+ۣ����������i\����de���s@݃���sƩ��Ӝx����c�^��4��წ[��Ҡ���9ւ��#��������pHܟI!��@���l�v���o*(xm��-��Tf���w����CZ*���HX��C����j�Ew5
>5�w��Fu�o	k�x%�-�� �3d��*��6i���{͡�Wؔ&ι�����bx߶��^ߗT|��Ш-���>h:��Z�@SA�wH�mؖ����m�삚�6��ƿP�"/㢠�?�fÝ��:�V�>��3xa�,���m���M`�k�r.Y�oA�/��Ϗ��.��e|6E=���a�B�1����|�����)��m����<�g���B_�r�+�7%��i�ݾ�c���\y�&��l���@���nk��&(��c�Eڝ�,Z��:@8/̰�[	bJ{�M׎�+�R�S�G�Ɋՠ�o/8�-�3�S-�'Ѹk�O�-V<��^���:Sb�|�u���?�1�U�^�R���>�E�0��yԣ"��ձ���Y0y�7�[@POݛ��s�dA��l�2�S�Yj�˘=7S�O/�KLa&�|I��,�5����k{v�EFѶ�>P�|��M�áW����)i�l�i��r�V�e|�I��C�i����?l0>�-���vd�Ⱦݞ�{�t<��i5���Z���¼�c3�d�6��4Y�q����9�fY;�:D��9�oqٕ�x���p����!�y?�,b��a��	���^��$�$�/�1a��~�X��/ʹ���c�֗c�h�7���،���;�L�������}��<~0�mv��7�=��������>C%�,�O��
n�4�8�@ڻ�9����$q&Wŏ,Ms�����WWgW憡MKsO+���$[^����w�q����Ot��'z��'#����{oU�?��H���)r欤-g@�:�;�����6����ש���.�e&�ױ��ݙ��}���oP�HǱ����N�j��@OK���C��e�F��^pح2X�p��;�C��������m�K���u��] *��}��-��>
�.Kِ+��g�]�[�3�\�_�3x|K�o����n��0y�+i7A=�ø�V���g]O���7Z����o�
��{R��R�.���śh���娦����H:a i�)O`�9|4��(��[7��i�_�������:6���� +ۀ�������DY�@���9�\�}���cz�Xn��棹Ov�g�M��Q<����(C����n���Ô��+B
�=��kEI�׈F`^ɐ����ְPRA���mu��q-�t�mK?Fk���̘�/;X�v��ǣg&�A�#�����d�q�|��L�i�#�M
�CxOW�	�@�/1�/���r��6���MRk�"����˷��4姣�xF�^�`�W�pL;�.������6�đϯ�~n�N;l=�	,~ux�o� ,~�۫�_�)u�,#.�|~�,�޴��l��q�//��Y��ٸ��-�,cE������g�4�� ִ�Q�b+��B��q6�Xx�-,A�:͸םeD�;�3O�,b�\;�Q���ٹ����a��r=�9��}��eS���ZO{3��/��O��)�@f�`XA=�'�A����f{���FD_�̌U�����,���G�HuK<�k�ݿ����aaϭ���h>�,��Ѡ�\��0䯺��Pdn���ĕ�w����K�� �Q��1�o6Um����3^�n� a�m�Txx�G=�@�/D�&���s̕��)k�>�Q5E�Ze5��xtep�?׿!��H���/�y�6����g�%�W`-�X�|P��]�HL3�+fs����l�m0��&nI���.S�ʓ��]}�@ڝ�Ʃ[�̲���gE}iy��bx>�;�k��]9��++�]9��v13/L��n V�l)���+ܠ/�1�6�4��<���(�~�̉�(��0��3�2i�>���H8�y-�����f���'Bۿ�X�����a {��fƞG�h����Z��gj�k��&���ߨ�/`��
�_/f2�y�j��&Q��E�o�@���e���y%�@��ۡp�����n�{�.@��ˡ�_70�r��c�d������:����"��μ�営��nI
g^��ˀ +�¢�~���'�ݤ�o=�	Q.�U����N�
#�7¸���H`i�(����}��Lu}����N� �R�q�̧( ��<��6�բ�|�a��P^e�u ��.0��ުgk�bqMت{�������6>՝t���&��9�]jVN(��Jg�^W5nVޔ��j]��/�j}�jN���`N锍�u��_�>o��|�U뭲�o>�fs��B�c]��Ƨ̘^C3h���w���|r�ac���#���KG$J���_ף;��s���a�צ���Ѹ+�{=��0+I��	���I0����Hx��F����d4�#c��)�!�]�7����R)��l�ױPƽ��`�D:��7���*�<�V�������IO�{�8<������&oFwR3�$��f�hbB-�T's��$}����h#{ #ێm��=a��a���0�}�eW&N�C���7=�U��'�AG�Ii��.�����`�C�'��y�~�T��C��o=/,*�>v�_�b�=#S�;����m�����IXK�z�0��g�Sz��de���%n����p��!4��m�pJj���l	��[_���<:YyU�,���0ͱ-���W��us�HX�b,����C5Y�%K�1ܜw�B��BZt�cH��`0�6�kn~P?��W�R`� +�o|�!�����br�Y�,���j�l�OE�����^S���w�E�������hҟ���8��1�.���X����3�;�t�,�����,5�&��7}y%������$�N�=�q0�0&����w-Fe9���v[!�N�Z:)���?{�d@�q����LbY��ׇ��ی�5�Y��y�&l�đдWτy�	K)�M�5q�'u���0�v��0sQ̺0]��:�⥂�ȋ_�YeU�����,/�-��įrH=�hy?��	Y��-���0>���e��}P��P�x��LK���43�Q�`��D�q&��3����6�鲌�[�CY�c��0�;�-݀}�msz�e����Ɖ�M�th2��v��]Cl�09��.@�M%�����c�,B��C	�g-&�(㳎�;�)ݠHg�7f9��|v��vH�otP~?X��&�U^�\`����,��v�D����¬qE��rP���a��*�u�FoG��h�<�×�7#E��|j|�V�x���x�lO�!�g;1i$��W�����Sa��d񅱾G�$;+d�ҭ?�(��Go��ɓ˓{}3�/����M�����h�a� `�݋1�)g�M��L�x��
��Y������儂N���!7�K�m��}�b�C�w8
=ivg�C�A�����1z1�bKg[\N���-[#_~��)�e��iim7���������ւ���­b#�kpcB�.�0o��5_F3T�$��o�۾�pn���ܖސє�&cH�%�Z��)/���RS�;rXև.G�\�w�������w"=E�m3��{4��@o1>�ouط�
�C�W�'S+,�;pk�Qz;�l|���%���f��̝�l�m�M��H^�!_�Չ��{(L�	�:>H��O�a0S$��0��al�̢�~��0�)��ԏ�`l�����]^aI9��1T��o`z��h�;X���X��Iۖ�p[C��1ts��8cc��3�5��Y�V��t����1tߑ�c9X<�"`�\�3nO}�1*`4��	#QJ`��)@�ԫ`K�I���tf+�q
g�����u�0_�~�	�%W�=A}�ՠݼ�ڂb�&�hEaG�w�{�p-��uOy��ת����\���<����Iϫ�C��?9�꽊��#ف�7��H�f�@&���7�э}�ly�l�S�2�l�ʴo#[�t�<��}���/Mu�px$4ZuFAZ�1A�\ˬ�e��^��kS:����zW���i|�l0��Cc�\-�z�FƵQ6�Q/�ֻ�"�1�M\)���1�)ʒ@�As�T�G=��Q�I���ݦ�u�"g�5��ٺY��o����r�6%Zczkx�tuU�J	��ݐ�7�@��������F�����H��,3��0�ߡ�\R��vb���_�HG�i:�ʩ�ӹ�������'d�a4rQp%�ݼ��<��J��3��f���A��W��Nz������#W�_H��U��\�wr�2�M@� �A�Do��=�)�g�j�� ��kH� $�7�>L�:�(�\H0�/�I��l�.�h�.���[���A|p����z�����ʝyY$uUvV�tՅז�2��%��?���f��9
���	g>#�E����)�a�[�k��كRx_�ۼ�������t����w�︸�IIz��N.��s����Q�����Mv���t�Y����������r�h�%�#F���	ݖ3د�-����7*���p_و¶��!][�0Uϰ�0�[C�PQ��h�0&c��"]B��͙4p�(vL�mc�k
�D4A�	�._������*�5��B�=�������|o5?�*�����4�U�k ��A���$�]r�:��+�J!<f1�]K���xҭ�!�\��BWS�=O�����=
�/ҍ�(�<l`;͎�����S +��`��$�c �C5��FPo�_ƴm��Rh�� ����ѺGUg��e�����9�{Nn�z:Φ���8~"�y��R�C�i��t�=�.��'wZJt�H�����L��2��k������d�xdk���g���ߡ
s�h�e��a�F,F�bF��9�������XF�[�3�)(����Wȓ߰v[���"�����}p���������U@G5�7��Uo�<N��z��-<n�;]e.8�a���Ap����O]Sa�h����
��M�l]�(X���`��|)��
�/ɜ���d�̧G-�����0P���;������U�a!��`��X�8Rf'��1��GI4�:����Y�7́D��7�p��2-d�w%���㎞��V�wr����;�-�[�[6+�߇v9*NS�@{��yz�̲��ݬl>!+}�<U�rċ��� ���XN@������gkпq-;�$�R��8~fVO�[V��(,�N��
��O:�y��R�؁������mڛ�>H����U j����(ց�:������R��TC�(�q��pA'��#4�qx��| ��(��K��l#v�
���:�?"���8oU�Y^�#s�*�4H�{�P��- �W�S߃�~��,+�� u$©�d�Xřڡ!Y;t����eQ^,�خ8~�����<�����	뗨�ai)�y�j��|�Y�Ѻ�a���������	�k}Ü��d��2y�u����_�;�~�Q"���2G�8ܿa��|��z�D��aO=!����)�2y��/՜�:��x_����	d�4n�Y|en�ج|=�2�C�a��,L�Z�G= z@������c-(ǰ O���������[���s�ޖi_b�u�p$����!Q�������}�e��{x70�vQ78�*�G�n`��n��ͻ�%��пq����؞�;��;��m��� *t,����z�g��a��ð�I��_3��i�a�k4��a����o���-Q�z�Y�?���	퓻�
�[R�`��|���Mĸ�/bxV��h��Wt@�n�;̺Al���|������5֟���}���d2>NS|�����/��ŃLS�<p�̬�ҩ;͵?\��rJw�t�����+�[�3�-�g�Y�k1N��O�!�U�M,��<�W��ް��h�-	���ە�x�T��J����C��
�66uA�M��T}����d:)Դ��qUWp9��s5�۰E&8���P�v������(ͅ&Kp�d�gn=�!+��u�����~Pd)�"��v���u�|ޡf��\_�s�D��M���t�Ff��My["��u��Cir���T�+1^��z��FB,�},�x�o�M��lƗ;�m%:s[y�^f�$.ǵ�=w�#��P�5ʇ�G<!��������w�,�H �Y��m��@���3p�i�)��v�P�6��X��/�ý\4��||��S���cF����|�jW�Xl�� a����'��m3[ξo�8�d޺�C��'Y���)�?_���$xW(��ɒ�ߞ6��������s�6�<9����1ܵ�z��a���je�C���&��8�z�C]Zÿ���En\�{�^��Y�-����s|Y�c�$�����f5m�\���5l��9kGj9e�IVK��!����P�<V�y��?�W�����<����eS���Ϩ�
]��B��fY��!��@!�;4A���UFz���E��Z�Oo�Y�<����pxO����10�~X����Ik�xT�dQ��⥢� ���W2�X;��|&u9dm�ԗ����_ֱ��02�!X�7~��3�&!�󓒺߾N]i�V����JVZ?����AsvxVY�>ӷ+���~����ȧ�i�7-&spn�zbS���iS6�Y��$>`�8� N����r=�V�6��l�V�����oF%+~8c[T���%���;�æ����t�F���?%ZZ>2��&���f�v��	&���\O<ᾏRfb��U��3�i���v�3+ ������ڡ�A�r^%�Ӓo�,�N���3�m��6sv�% �d4��.����ҫvne���6��n���t5>�{��֞m��QuG2[ [��2�:��u7��Ð� _+v������d�7����=�mΞ�D�h����ͬ�H�z�A�t��|3j)Ro@���H`�����9ܢ��~��<�O�c����R����N�|��ܻ�%m	Z��@i�Ǆ���$�-d�sļ��(�}8Nl�.M0>�q)Y����ھ�=����0>g�m��M�jU����^C�"D�j����׿�!�zOvg�	��A���a���J�<�K.��ؠK�{8�m��F����J���>����i��0j���bfl`b8sm���3W�'�:�G���ܯ��Py���Mx�_H2�Vc/S��OT��3�8O(4�9��i]D�N=�z� /�d��;��_�� I����~̬�]��K9���Dǫx��M�m�:+ٗ�v�~�]�������g��$�}�l�a=�����d���Z������B�Z���|�)����|�B8��a�����8� ����Sʫ��PÏރ9����P!��/���D������L��hs�����J���W+�C�>cE�r��Z"�����WF2�|�Vv߿_��M����/]����T�̉He���>�g��d_�D�AG�U�T�؊�����k�����k�׻��.k�Ҕ���i=����?9J���$6�CVߟ֙{��Y�E���tm������8BP�u}bP��S�	
E��n>�lg�ySt�����o�C^�NGh|��H��x�a���7>t��������%mQ�mdr7�Y@���t|�<n\�Ӎ���o��<��p���TK\��C��`f�}7jf*�&�Ms�[~!�.��g�/G�f���z�10�8/��x�b.<���G����D�3�UF���Pǻ�)�O��c��;�0�ʐz'���<�����X��$H&4�]�Bw�Z�?)8�J~g��ՠ�=O�.,{�CD����vT��)���ը�k�����,)4��=���T�R���E����;�O^t>Ѻo��7�u\ Il���$oIl����T�7�_ ��	ȃ�������C�%@�(x.� ���sT�ϰ�Vt7�(��E��)��}F�foY��ź���Ӓ�Y�9����E��O�9B��?++�퟽8<�w���p�7%�����
�>�7t��ǋ�q�֝7�8��`���� C�8��k�ɥøˋ�7�L�L=�F��‒�\�f��_ou���bGc��ƒ��6�C�G K��&�fJ�i-%��/PV�aH�~�R��$�����i���!�����Jf�o���:a�u��fr��Ff�:�CX?̸����̙׳�P�Л���U0�O�h:���R���I���`�;�c�w�_�\Y1,Tm��N����)��`�hs�-�kپw6o�PKqoE%&Z�����`ݷ��<��v�a"Ǟ��S_&�`h|vL �+��I�Ga4;R�6��a�2��m5+\��l�I.�t�b��g^,�x{��`W�ر ~������P�X���ZT�ls�������Eh6O���4 ��Hq~�eCLJ��Ù�_��=Z�U)p0��`��ƟZ��lk;��sx�`����B�J����	̙�^���K���	�F�﹡)��(���lY!hÙ��Hq����u�<�L@��Vx�Y�9����
����\W���o%���n��[����:�v`ˊs0�����\���h�Z�|E��y6�MP�P� �S�]j�*�};�Y�y'�����"���Ta�<��K.8��tai��r5�<}y�*�T	���^�|u��	g:�����k�R����� ����$����d�a�uݑ�]�1	��P�r^����8����މVŖ���7nvf�9�>�t�@Qz�� ���3&��qE#'��f��p��ٴ��%p[	�g��҂���������Lv���п�J܌���)���)ˮE�\�>�
�ځ|��"=tQ�rІ�8>�*�{�fe9jwd�������r��
��|OOe��Ɓ.�U5��|��YȐ�^~G�v�d�r�!ծ|`Szl�)
�_�'ǣ0���.�)��ڜ��ð��x���ݦ[m(X����u���6�(�<g��'E�fea�]r�YI���O}�ۂũVg�����2�^�g���C��lk05`s���A�J�Fs�����t��V���`*ƫg��aH~ۢ|�{ZM�Tl�����`�,���*GerX��P���*�ݹ1�\^��
�y�<������@�198��MV��58s�U�3��dJ�t�sa�M�k�9h}¨���'l�F�gȗ�[Ǜ�ޔi.(�o5����O'҃hQ*o��(8�~IV�G�x��C�f�Y�d�u���^�5�b�c�G)m�E�^���� 0�}���]}�]S9��Y�IW��*�0�=��r#�I��4���S�[��qB-x@�%��Ö�'|o���^��Nֵ��*{�Q�:nk�|b�fOp!������&;�ز��^��}�ύ�؟�F��v��&�&����,Vň��+o�S2�n*���&6Vig�y��6,v'��y�1{�j�
�����VC	7�~�_z2�����V!/5��Ū���>�y���BL��gܳ/��qk`�:U�/��V�V�Sm�`���?W2*��E�#$Q��ډA
���A�{@��-K��
����s�p[��=�p�(��Y؅�<�i��:��7�8;��K�����Z��ۘ�v�8<���Ԁj�/ж9+>�����$�*RFX���_�2��(��m,�٣���IlD�o��q���=>�g�:k+��Ǆ c�dL���$�M�1�t�9�1�	p!`a-\�p�1��^��+K��sXo`lh�76%�z+��7���3��˛l�X~v�٪�7�h��X� ��i0>ۊ;�Ѱ�Jk��fS�����OY-}8���h�e;�
g����bmq�V*�m]Hm�ӭ���~
���ߩ`=	|;���!��̣~����YIdú]9`�1>��栦���a5L��Վt�˩[��2je�2(0Ns>��z��1K�[�Ȧ�X�P�٪�9�E,��,�ÐzZ-Q��Źmj���Е��Ġ�R:��ӷS�BBz&g��ܷǭ���;���<��t��Mp-�����W��`
$������vB=[�D�?C,��	�"3}b��'�~(�=hMwhc�g���.�g�%LʐM��A�W���'e*�"��Yu���z�W���$��1"���;�D yhef����<�/^L�\4+.Q��tl�����Z��.?k����)x�Ӡ��5�?��a,�_�>�o٦��ȷ�`	��Ɗۘ�LBc�f�­cq:>	�/B����1���_oJ*��7%�;���dl݈�ǭYzc��؝�q��[���e�ks����	�V{�N<O��ǝ؎{�U���8Ϯ��]E]��	��o���"��Z=���I�S+��*�ݗ���B͆Pl�ٲm�-�Ŭ��7�nv{�X'�����6�¨�A�mi�UZ���k��a��R�_��Ez��˜_���NP�"���{�j��h<h_Hgff�����?��-��� n/w[�]��9��X��M�[!�9#Q��s�0�;S��\�L�[6�h�
�216� �g�[����j�iX8^P����.��֧������V�`�W�GѠ������y�]�/+��,�Zۍ��U�qfbq�չ$��ogG��C���Jjz���ڻ�v���v��2�FA/�[�,GU�h�|��rH�	X�[۷�*�}���ՌP�6K�]��p(����+�Y�۔���Hnي�<��<��7�ق���r����Y��� �QФ��=�x(����+�G�<�s�&�z�M	�Óf_�voU<&�Ӭ��jj�t]�=aLt���~������"z���y��1�7��͏t�̯��mV'%�\_
�ߞ=ذ����O��pk�ư B4�se ;��Jܗdd���CU�|�H"_����,�v�j�C����(�@�!����?y��ϫ��<�|>nm�暯޽�������y���:��տ�Bc��c�����| H�M�ٕ�0�[&⭑?^�Uz��%�����&y��\�ӗ��&��}���9��E����9K�����u8Q���7��gq���P�޿�M��@	h$��oN�ޮ~�vϰ�{�Fw%~1�Y�g��(1�K`(>SسK�~;��a����R���O��Y�a���8��9�3,�2V�b=���oJ�����{�(�>�&�������g�v�D�t�O䵿i�45�������ۋ��6�Z�T/�ҹm�.�|��8!�^~�8|ɡGB�zD�>�¨�}?���%��]�Dd�qאF>\rvg�h�О���p��~8�w�5�j e|aW������2l��t�[ԣ_��jS,9vgC��߭��V�#��Nk�rcr�g[�Vg�=�ݤ>�|�ٜ#�:�ů؜�w@�A�Nf)�Gm�Ʋ���h�g[{B:�لp7�m��Y,l�m�33F���E��/����;a��?��6]fw.�[�K6%u�ݩOv��k��V	�-�ڕS2ϒ��I@��H���`�ݢbc�{���{|���_��5���7):�gA����͢��&f4�O|,>~34�GIUw`���v����}�)�/֔�7�_ۿ����1�lxe��čv8�j*�if��+��&E�<�=F��zq�<ԃ!�5�[� H�F�/�j���-@a$���!I@6l�m\!���]˔�7��YK�Ϯ1�*��Q��˛3��9����,�40Ǧ��4�Eȯ�x���?�a�����1U�8Wj��7)	(O8`�zNn�ʻ��<J>�D���I��y6e9v&���p_�����v[��[���=P��2�d��=Ũes��Ԃt[{17_�:�������Q��y_V���i#��Ur'dZ�~l`!��x�9ʣ<+.�S}�ɔ���֟>6���q��,��u���y` �;dP�O\r���%QSL���s��xu��|��lN�_<h���ι��]8��T�Nb{���� ��ʆbk�&e���hVe5��ٜ�Үl��K����컙��{�����Y�V����ҩ��mP��3�g�=�J��VFv��q��iU`(���ÀL"�%��3���Ƈ���
�؍v�0�e��g��V.X|?���'��j�2|��u�ɬf)�z�J����ܩWF�3�㔷	�5��o��"K;�bv�<;�B5�s�]�wK�&����x�2/"�_nš����d^����S+�b\�bZsa-�?�8�Ѵi�>�B��,j~u{������P��m�c�Ars+˄�I����-)j�p��W̸4U�B���	�x���ʫ�x�R�0�W��P��]9�V��>����] R���G uߝx&���-�1)��񑏘�>�%�`.�~�,�;������+�ʬdb55�S�^�NT�>���+��|##�gF)H�J���vq:�/J�Ǒt�=:�zGq�!�2���C��Uf���m�fM�#�Q�)�9Oܰk����Ѵf��=Tޛ�ؒ���(yEw��M�91�|�3�d`��/P�P���EV$����(/﹞]us-�}K��k.@���u�t��,�/�ڼ�Y�;����L1N��|�\$�[�f[���]��UalA����zXDޟ����{���s 	_�C�&�gT�x�W9��|l�_?�,R[�X����`�@I�]`�&(�<��ހ|�)���.�:��b_zn ��d%iv�2rr'[�z��4I��jg[{1,R:�O�-�oN_�@�^ۼф5^�U)��7$�Xug��
2���8��#��#�;�ϊ+��p�O�y��b+�C�Cv���c��q��xL+�̓�����!b���~�W��%��*�Oy)��L6R��`l��X��������8-�-��?X���w������?qV��M>m�ҍ�?�Ǩ��p_ 
[u��K���M��'��ޑ�Z��	�|�\��t<A�H��6Z�s�C��[,��;=����%�W�����r���e�7��.�BI�{�7���N��0~:p�>�?t��bWm�~�!Ih���Y�1M]�g��$��(�*f�^��ٜŘ�9���/���A8���E/�d�o��o�
�l8�-�$����.I�뿑zEY���n�ޔ�7.�q��L���`w�d-�v,pf���[>�d����n��g(�r�
B��w�bNׇt���m�3�'����o��>�Α�J�<3���Z����a8�S���3����wm��}��L��@$�����.�+�O��ͅ���=�� �{G�s���]�4�*������r(�#/�|�sC�o�]i�Q/Jwԫ������P̻y�0	=�����j`�&��<̱��ǴKy������d�v���7�p����w��*i=E)[�S��t�o��鏼�����BBnosLv���:���X���S�ͥ3�7o�29�tX��:���د>��᪕��'�X�?�x(�b���E���̡t~�Nr��q���K�t
1�����VZ�Ӫ��6z6ٕ ��-�8�j���Z�q�W�a��Tb�8�v[L��(��$�9��� Bc{�`b��x8�y����W>�\>�N��/��		'�&|���-�X�9�o�:�w7���w�Ի-9lC.䆶$TPS�,�(6A��Շh��$��*?:�f��4��MQ�"�q��j�Gl�OA�����/@M��vٚ$��Ǫ���}�m��U�DQ<�=ϒg|�=���7���ԫ���8��(�����S�dsד�B�vrw��;r_&�urO�;D��r�r� �J�Jr+�m �arH���L�[��^ w�k"7��5�{7����&r� w�/�{�܏���\��)}ro �6r��.%�>r�'���m����]䶓{�\��ğpw"���[Ln9�[����!�ur�"�<��;)]ro 7�ܹ��[In��!�)rw��E�r�B�iro�v?s�/�sl������u�~���?;���{�q��ׇ�cjK`��<|�r�)+7�UW�9˼Uu���M=<����;)�iyl���j�6Ԛ\NW}T8�W.�(����=�_�
���d��lk"�~�L�.-��)��R%�"i�uR�����e�
x.��J(�2�KZ�*��U��y�*��̋~�e��3�x����'�q�B\���	-(����H�2�$׻�m�@�|Ւ�[+����N���n�dv9%��+s7b<7{���Ҩ��0�Z�f�������U\5k\n*'�_��~��iXv �8�{����E5�r����>46���zGM��W"�$���e���+�o9Õ�h%��*�L�j���ty���x�7<�ژw���;��/��!c�- T�»�5�eG�������V3����낐@o������Z�>�j���;�џa�TI��_���]Q��rD�����^�/��k ?���+g����7>�(�{Y��RL./�C�	hZ��SN�7J&MڛF�~��; ���4��<k��.�z��$$��I#FF%����6��;.#�˳�?a�WM2]}���)�^7����8}�M97ߒ;���n�˿�`��9�(���-��[m��/YZ�l��+V�u�=���oui�g��bme���kj��p{���ܸi󖭒Z;��$%
_	X����A��(�H~4o��ߎ�߉�ߍ��$��?�a\��K�,&n��6pO��\�h�jƃEunKC���]�ta�_Ǹ9�Zʕn�
��U{d�n��<�˅�|��βj�K�/�ƶ�*oUYuՃ�"7<9˪K\N�o,̿��*�,�]�^K�
�K\5e��un{�?��J�+/�9�͇!������ܫ���zYU���/�gEY�w^�;ί��5��G*�����E�`:R|>�%��MG�W��T�W E\s}.��Q����5n�2VT�jE���`:��P@�"���D�܋|Q����"�5[mE�����oc͚��*���v�
A_����W�5WW����Hu�*�V.K�����s�d�j�G�_]M}��U�uWծ�w��2��r�G�Rp�4��_�q�)otQY�60�<�KU�y؋e�Z�1tr��u��=�U9���j���dx^/�dn������X����N���.���WOx�>�Ʉsn"��p�1��	�%\���8��	g$,��қ9Ox7�	�M�p<Q�G�*�?�I"|.�i"?�W��fr|���8n ����A�~����3n�8,�'�T�Mʁ�[�4��t(O�Jul����j-����^x���Y�޸��'ty�r&u�i�I?OK_�p�'��+Y��gP,�nb3<��5,��D��~���>�X5s3YJ��O�f�/�/���~�t=�Jx�w�j��	opl��Etz������3Hg�˼���ޮ���H��d�]��!l��T��0[��|�f9_ܞ7G����W��/�N|z�1�!��Y�Q�2��z���V������R�N�i�A��,/�R�&Fo�L�������V-�z&Ec��׼L��f�`]���b8'��H����m�Y�&��XN�C�eZ�Õ��#?��f~y���/N��c���_��ݲ�z�V����7k�e�����.���)�gI�ܧ��qks���j���Ul5W�8��Vm8���ccp���Z���8
Wk18eg\b�ɍ��ߵ'�H����\�-����'�Õ���uJ$�d��]N��xQCT�"ZxX������؊��Q�T��,�HZ���o����\�����X�� ��O�,'>#gTD��f�k����!-�h�1�<t���ԮvT�гlXJղ2���uݬ,fV&\uW��h���Z�r�V��]$;D��|�\�BOg!��Y��T��Ȍo���x�+����3����2��bU2L��pnF=�O�O$����o����T�a��h-�-ckt�;��'">�x��:�7��9,��+�4���܌��_��w2:�Y�H����Jj��5,�h=���L�N�~/����
+���2�ol��߄�7:�CQ���⯈k��&��������Wb8 !��/�F8�����O���~��*S�c�Z�H��߰���OS�C���o~�-�My8�ȣۿ���>������<����';���~������կ�����v����������<���_z�����}�����ӻ���o<�w�țo����c��=����~�'?����X�$��g�|��_~���g��~}���/�����V��K
�����O��]a~i�����$�?2��[D��}/�	���:�턅p�c�G�'<��zo��o��X}�н��>i��[��p*�t�i����>a#ᩫb��9�b��y���b��V���	g^I�2¥�b����b����b���b��M�b��m��$�}U��qǪX���U���]�b���W��M�O&����	��B����_G���	����Jx�A�7"<��t�74��p:��	g��#�Ox*�9�s�p�B�e�V�E��	�	�$<�p)���+	��^@���B�M��w�6	o',�� |'ᝄ�s����݄w���J��p =�	#�#�������4^�"l <��(��u4>�#�T�V�i�WM����p�t�m���0��0��A�3�"�Ix���g���BЏ�xA/��Ji|�"|���}O�!l�!|���k}O�!�-�Ox��?�kE�	_'�O�zQ�7���&�O�FQ�2��p�[�I���K	�F���턛��N8��N�w�M��p;�9���p?�B�o�e1ᮡ�F�a�ho��ބ��&<_�7a�ho�D{^(ڛ�]�7�E��	/�M�X�7ᥢ�	�)ڛ�
�ބ����I�;�u����E�	7��N d%a�H�?�$\I��7N&�F8����wGx��=�/#|��x�*�+E�ʉ�	�. <���y��[	�#\J8��z�z�M�G�Nxᝄ�	�&�J���x�}���UQ�C�<$�\T�Y�G�Jx�<�Ʉ��S	�$<�p%���H�k��!�'�K�Ox�ȟp�ȟ�1�?aU�/�
ʟ�t£�'�!�J���x�ńW��I�l�n��!�#�K�G�]�g�O�G�_�GxP�',���$`�E�D8�p�"�T���O�T�'\/��$��.��)��p�[�'�.���gR�Ex"<a����N8��I�Ϣ�¿��/�	�
Li��V���v���$@�$��D�'<�p;a!Υj	9\��=��b�)~���1�*�w	�o*�w�"�(ᩄ�#�6a+�#�W�O��'�@�U�m��#���X�",�'�!����Q��u�1��� �u"��u��~���2�n4�"�.�Jx����������"��(%���'�-��qz�&�'6��Bo����"���	�&,�M�O���=��m����S��X���-�u��`:�7�?M8�p/�B��!\Lx��'��=	?#�G�A/�}�^�źq7�vA/�o��?i�������?
�>*�Ws�_Ѓ�=wz~KЃ��=�����=WЃp���=� ��������$�O���?�.�B"�&R��<�?��H'�3�?N�b"��Y轴}p�o�)���_l<z2�G+&�������C����Ἕ�w~Q�8��n�o#,�BO�N�B� �xB��G�B�!�6B�O�b�hC��m��KX��X�=��P���_�U�^j�O�������rȿL�7N/YH�BO#��BOYL��.%����S
=f=���B�%�fM�/��
��̈́����w(�Lw�I�����M�I��vS� �v�bߺУ�B����}�qz�~�_+���%ɿ��T��#��P��ɿ������Л�&�C��$,�n�>��"?��R1���p)���	�7^NX蝅^z;�?Ax'�e�w���?N��N�AQ�8=j�o!,��b��O�B�(��B>H�B�(�s��`:�	��DЏ�.�Bo.���R$O������]�^T�Y����*��%�&��E|�?�qz���a�'z���_.�	�L���>���wz�#�� �=	w�	�w��+�'y�C�9��I�J�%A/¿ �@���>q�-���}��S{�
�����,�Ѕ��俍�Г�~�7������ɿ���N"����}�%7��<���"�����j�B�+a�o�������⻌��SH����w�l,&��$�����"��4����D���|�	�$�Nx;�>�?%�O�w�	�����X|I'\O��f�54�;i���4s8I�)'�r��\$I���\��j\A�WR�Ji�(\I�S��2��n-�z���M�ݔ^%�㡕��V�I�$�y)���*�P�<Z}x>���p�s=կ�f�2�A.*O���f�u���]I�k��(�:J�C3����R����Z��K�K�_G�P�ѣ�p-ū�pu,G�!�َ����th{�0��ti���t�s�M�@�@~r]9�7k� ��b�|3Rr��t�R����Jߦ���GӁ;�<]��i�A�B,��Z��"-~-���3���_�����w�s�K��n��R-�JV^���P� ����/�_��K炭v3,��1\���|��3k�����H{�X��<�a�+���b��h�W���5�����5�U���i�Y���Nm]��`�v"���w�TpG�|1|S������e�U�����������+�c圯ի���<��*Y�mZ�kX=Z==�n��a|��踎�w����X�j��-b����a�Et�|#����;R�z���kY�#����9w^W��8�����jX|������5=�Z�^��xI��+�q�r||�9�=@��K��et��ck�E�˨�b�Ǔ"�����݄��Ǔ�Z���!���Z�^���e�/�'�v�q���ud��E�&����9�����7���,���t�h���mkܸ+k��t�5��t��#�S��������z�rS�x��Z���*����e�*GmL��\��wL{UR{F�Y2D��x�f�x��=E���6��\4�E�'wLy�P{��?/GIQ�����O��_A�>ۣ���|�.��2�\q�(�Ǭ�?:��v��Ɩ�6��tDa�,Z���g��wE՗�sl?-�*yb�h|��ύk�b-}~���,��=���Ƅ�G���mELx��<��(�Z��5&|�6���r\{/��SF��8�I\;΍������l���[\���H�_-#��)_�W��h�e�^��5����rmɱK�q\�}���~m��:M/�q��N�1�ĕ�N�+q�@���"���]7F��AV���/�﫣�'���h�s�y�F>�Wi���d�{��p9[�������������]�}���\����8b׃�r��Wk�U�}��x���V�o��P���x�V^��Z;�&���UZ�8�_kg�k�ү��ǱW�?�>��?W�5>���,�~���b�S�� p�l��8���P`O^U~ĕ�p\��9��ڏ����q���8��=�ڐc_��������싩_GTi��u_�V^.�Wh���q��#�#pe��J�ÿ4nzs96R>.gG�%_wF����C����m4������J-�N*�����4�$_�Vi��rj�~Wi���Oݯ�s��g�F/�^Y���uq㎐��n�j�V~��Y��[|]X���׍�p�=����F��:$�?��k��;Ο��X\��_��h����Z��\��k�����#�3���j����j{Y��\��G��b�X�x�E��z�V�gpk��+��#���H}8�h��z	��\/�����?���"!�F���_U"!F������D���W��Gχ�����ǆ_G��q����;�c$o��4Dp%�_*5;�xI�pk�Ӟ\o���s=O��>�;|������2��q�I�<\������1�6&|�V�k4��أ�=6hا��#�ˉ��l���l6�An撳���uͭ#J�]^��Z�ZQU[^����)�л�z�d�g��]No�!����^�*�� <����Urɕ6�w_rM��[H��ܕ䖒[On���}����$����"�irw���{�m'�ur��}��c�Gn?�����)���~E���ɕ��'�@n*���f��E�DrM�f�;����!w&�y��"��\3�VrW�[In=�M�� w�����+5R��-$���6rw��G� �YRyɵ�k'w%���>L�rw����c��k�H�[O�Nr��U�M�D� �~S,�m'���r�ɕ6����k�<�r���������,����x�Wk�[Y剼X���m4^�Lu�7�n� �W���T�p�^�m3�u�<^w��+��j˪��ֺ�%|���Z��$S����u�}s� ��{�fË���=􁴮��.�����9|�дi�<����}�2���'�߶g��{n���{/�^Ͽ��wM�y-D�7��4�?����`<�4��7������
oٚj���X�~MF"]'�z�]u�T�&U�M֜���2w9�+�0[c�p�=�*�އp�xϚ��"ć(-��LκZ�arV�y|nV�Rl��ҏ�^��4�.&�a�5^�K����^P���S_]�tոj����zQOW��%>ܰE����E*u��7^�h����kr3+y��J-V�t�eBoC�qE,>a�����J�u5�U&�!OrEi�H<d|����Y�������F��p�l�����\Lz���F�m�-���Q�vt�@J0�z
�2����]��P�|����_�q����Oҏ��^f�1��K�e0>��.��]U��i.�������Z��^�/��e��^Y��ngec|�&4�����`&�|H�7O.Y$/B׶�,qws������`�i/���=f% 3kdUL�?�h������n��4�$-9�۵�S�O���{`�������<^SEYU����̙c**�/a���*�R>C��^bG�~M�˽��.Y�р��,u��y]Eu��ht�����[^b�ž�_����yԘ`�����.66��e(薀$�G����ٵƷ6�gM�
Z��ZGՃ?���i�R��	e�m�����^�ƻ(�?R���E|EQ�x:I��JK%������BE
O���Ǉ�Ŀ�}��q(�nQ�8L��|c	7k֬�����r��a���Z�s�Uь3�?ک��U��Y�Av��~jTxS����(I���}�i�W&o��2�ͅ�׭E������v�����E��J��]j.6�p�Ճ�&���s7�9�a�<|9���5U ?��Y�`Uh��k�
��(�T��YY���<��5��nMY�`6l���C^&l��d����L0v�x��g�WWO�|)�;�����0�°zqɁ�=���t'G,ר�J����޵�GU��o�b�"�`,QJ�
��jh��F/Ȓ	VJb���<�d�Ѣ�
hDԵ���;��W��h�F]*�Vm�[Ko�b�^�k���3sv7!A����'���;3��|�}�͙s���N��C~�h��W����E���]^z~�v�='���g�J�I�[�ƨ����VK����ڳ1	IF�'�=������꺚��Jcd�N��V����dY}�ᢋP�hV�UVo*-Y	�5"�2\��M��p���e�U���R�����
����H�#�vI���f�ˋ5�p�F�Up��1�E䋔?\�H�p�6qE���p�EIC@��p�=��G�A�ץu��r�g�[��\�\Έj�r�QBA���|7�UF_����j�R�g�8���x}r���\�?Rk1&�յg��'D������%���pI�Β��"����R�M��=��oȑ黶��s���w���0�Vǁ�\b�x+�;D�2rov�F-�K8z��i�H�iuCw���u�j��F�E����"�j[G/��;���f�#˔˒c��,j�~�6��(���+(�Y䔞�w�������Y��"���F�u0��D�[v��V�h�1����EZ�U���|`^�I�����$��O�����Sr����?���t���u�gM���q�RQbp�)�<^�+ms-Q.4sbM<�����)��jʝ@�!��0 mx;WLI�)�D�R��)��h
d��7)�H��$ș��`�99�&S�
m�/M ��hRy	DH#�ш4�L���������q�	z.�bif�Sj�����S$~�2��UE�G
�����y�V�=�7e�;�2�v@�������4kO*%�I0�86�i&((�j���dy��ȟ�����r�<��E�7�i:�V�J���4�j����l�e�M
f2�U��:�f]*�3���f�Q���#�)�W)���2���'ῷ+h�x��Lj��9��@|D��<~�� �G�C	y1Ҏr� :+����)�TEY��)�!,�I1)�&!~�'5d�T����/jr��Ҕ�T!��@R?������i)4͜NӪT4�4��!��=��������&K����g�5���)�W��4e�0M(��X�b";����D%^��vH�L��L�132g$P�Y��Q���zͼD�n�9M�z���?F��Hֵ5�(]�D�g��5�k�<���I��y�*�v 2�k�Hs,�4f`U"i�)����CN{e�_3��5zU�+��}��T�M��vi�	�3?����(z)Y�����H�ϥ��a�����hd���&���3��hB�h�F��!L�΄p;Y�ӸK�6�g:��F�h���_�������fJ%�g�-�ɕㄎ��{
���j":V�������$�Ǵ3����5ܰo"Z-˭M%��5O'm�4��g�V�&��`cі7���(������9��1%QZ1�`�I�A"l �}+��7�R��
fss*�B�R��4�x�����#e��G߀]5�����_�?�^�m��I��+���ij�j���"3�T�"cE:���>�S�e=��M�wj"�"�l��HO��1�o�B��b|��K���I�~T��r2dK]1Ü��i2�&,�')�&��cD�,
�5��S��R�òNE�d�MX0�ad>v����B3�iFU&��ϠGFJ�����|#:�NY�L>�r,Q�	�K�T�+�T{RLR��&���b\�~�2�4S(E�N��X=��Ҹ'�2��x
�d퉲�:�ߖsp��Y�%����G��8���Ӟ�5! [1�^�Ǟ���	��~9��w�sa�D�or��CD�q��������''�da���B���@jrX��/��=�qc��q14N�#�9D�[��t%��Ia��EQx<�8X_����)<nd��u�H�Rï�Й:#3(]�ص��\�)��d�ğ��	�.�/7&r�bs�|����*��Œ>�X�ꛘ��E�-�g��|�_&�ӥ�%�mJi,��rx�A�|���D�U�������2���MI���%ǉv"�뜨����41/=�dֈ��}��a�\���4+�1v��;Z��SY� �8i>*�S���{d��{$��OD�E��(���'�t���x�q���318V{�>&Z�q��|���1t,ϑ5ٱ��>����'�cH�pfx��a��<�Q��P̃��ߓ��I��D������9���z�L��"�kއS��d��~��~��~�kG�~B"MPdPx�&]"ץkU
�a�T��<)]A�d߉�qK����VRv��PVpJ@�?�4�����s]��b0O�eq\����˙�L3�g�L�$�9�?ՔR��
�ϥ�8>y���RZ��__zS4%���H��?�4//=i�Qcɩ��U�=�K�c&B)�\��柒_��_�¯SH���:�,���xuV�q��xƎW�K���ϼG�������e����}[��w�q��g-=��,��ƐCi9Svh�g��{&�zo�Tk���!F�2��#�I.ڰ�6����X��{J=��K��|�O�VAe?��]������ט�W�s�{�k���	��h���ƈ}�J�g�qņ�*��$RǗ�7�R����y��j���/��>���|�C�aհRW�W5����ˌ����7Hd[��b����!y������ƴ �����h�ǝ�-�<������4��d��q���IO���5�%M�H���s_nhFi�#e��w).���B9�M���e����D^�\��(�m��B4`�������vfۨ:R����}�%��#޷\RU� ��y�d���ۊ��W�\�'e�-��FS��i	�-YQ,�_s�0K�_W]eXf�h(��~�]z��@�Ɔ��z��^T����B5+��K���K�X�14�!�F&ąw����vP6�i�E�
�Bt�bE]e}U��f�G��+6��+K�f��
q��+�у�I%J��RS��'��ڢ���@^&�e���f�^�b��ڡg���:E��1�7[Y�Dϱ�s��̴B��F%(�K���Ք�\�&�fϴ�\�⤟L��g��J��E%Z��T���&�)sI�T'(��RV�m�n��c����/�O�L�%u1].�01[,�G�쏰�����5��4�n�uf�S�R��o~����W���uFIUa�C$���l43yM옻�.��*1U�Im���%5����ů�a�8_�yv�û�����{�negRgx���������YF����+��0��c�cv�n���k�R�+6p�NŮn2����e�g��#�dQH{�2+��z}��S]c}����Q��*�5�i6��%�w٦����F�[G��<�[s�&��/oz��iv�bk'�s�X�l�F6d�2������l@�"[{M)0Q`�HK�J�$�2L�D[,C?S�K�/��Ĺ^�)�%׉�׋�kD<�~IK�^���� dM�-B�����D�vQ[W�����8�	y�>��T���HM���q]�:��՘O׎y|)���c�g����o��+����W�'��:�"��D�� ]���m3E�K,|jtn�qP��YwK���?�~�];F�[?����ɿD�>�d?f�B��ڿ3&���D��e͑����#��;����7�Ϳ��l�)�A���"�(��yb]�\��.��\`�@��2��M�l�W�E���=;�
|D`������.�؈��xB�'���w>�s.�X$�L�I�|7�"�[�	��
���'�/p@�@���S`�@��"�z�e��6l�*�M�E�U`�@����
��ɨ�
�	,X#�,�E�E`�@y�c��������F?��ݗF;�=��B��Ţ
��9�:d=��ɧ�g�B~�d!j��q�-gn%�W�3V�ن�jӗ��E������������6��ё/oG�(7�����o�P*>9}��߱�"��X~����5�GK|�o��3��-���/�,�?:�|�|خ�*�̃��}�>+�ou|u|u���s���5F����ce��=���Ϥ��sOd�t�}�I2������qO�zg>�m>��ԧ_�\�=�3�7=]��Z�pj��ܹZs�6����v������'����5㮭��=��׮�N_:���Wt��w����%���Y���׭�}��M�-K��q�����x�,�����~���o����d�P��w|������?<���n�������=��m�����T�䔦��7m>T��l�1�=.�V��.Y�����7,��О+Oop�l��R�*~uj�;fm����k���?�I��-u+��~�b��̒�y����q����I���ؿ��+���z��u�}P��+�4o�M~�W�UH;g�%S/�<�~�P��W]���n?^�`���7���{���
�>u�Ŋ��7�+���;�]u�������=J6-!���y��{/\�5�'/�-<��g������;o*�X���[~R�%��_{w��'�|����:�x�s��n�|���N۱�U[.���ە�K8|N����{��?�HsS�e��;���m���G�^[�zk�r�Ow�+v��W,��νh��Y/�s4��Kۮ��u���8���?�{��p������?�:o֥�期������fݵ>�����7�|v�Ch�r�݋��ߖ����W�����7����_|���k ���O��S�W����Wǿ��?g��dn�+����X�~�5��t�1��ߧ|[�acuݦz��U�he}u��������a�{0�<��($<A:���ΉD�A3̝DT�x�M&2��Wb2�t�ws4D�?@8 �mDq!���-VN���N���3���XKT�h��3q��l�&����"�%B� ��sq����YD��C�g��v���^
=���1e/#Z�K!��ԄP�؃�������?\�����c9ϻ��
��p�%�A��G��[!�ХD͈g�s�gx�*Ȍ�r�S�x9���D�����!::�~��U�-�D� ���b��|��ܭ��ť������w�~)�ׁڵ�-��*�>�,��|k-�?�}�s� ��!�u��N��k��rJ�w#�۠+��e���]�����D,Y��)��������c"��J��*�e~�~�����?��.�gx�w�[��7�*���/�s�]�"�x�� �о	����[�������~�`����0������X�W^����*��k�-�fR�	9�/!t� �!���������zo-� O��r>��6�����}�J4~����� ���yk�����.�a�{<>��臍�� ��	`����p���� oF_E���l-.s�����d������
�=��q�緀�2 O���[Ԩ�4C�D{A3LmAhp+B��[y�Z`�V�^��s��K�m�^A3�w;�1���
�8�4�����*h�[w��]��v�� c�.��7���.��u��B|���;�~ڀ"!~�N�'�Š[�޻�L�{���A��s�A�����s��Bo����� �?�1��A��#�2����Х�$�S������[����\�ˁ�AN�~�G�>���z ���4ù�	}�~��
�>�J���q��*��}��!��	\w@3|��� �0Ƃ���i�O����A]�?�6]:�V:���D�a����ہ�x��K��p<m�W��my������y[���Ch�^��] \{���y2��웈��w�*`�t.p>�a�:�� ����s�����dx�\63�)h���^E^�{/�>�8)��Q���Ͽ�����&���=�;�E5� �ߠ�O �^�z3��5�ǀ9G h���u� >u�������n>�:�� P����K��.h0����o�v5���F��@e~�a�OD�>z��}��!:w/�p�	�����9؀`F����臠�C�������!���\�w��?���S�}į��5c�D��}��u.�;'y��n9��d��I��[ϒO�����	���S>�2"d�f�w��ہ�FXz�4��)����7!0� �F`��v����O
��d���c`s�����`^,ƪ�һ�kc9�h���:��8�<F`V"l~ǭ�H����}�-��Sas��;��C��/w��.Ի�V:�?l��� ~3�2�zǃ��>���L��!�f2�3X9��YB`c�Vyt��}�ʾEU��x\�����f8M��4�Ղf�(h�w
��O��}�4C���T0[�/4�JA3�"h����O���QA3dߨ\u/G�}
�gȾ���^�>��)A3����:��C!��������Q+��ǿ��%>1�GWF1�)�%�-Yr��Fi��bi/'�V�Fi�y��_���SVN���$~į&qt��(A�o��J1[����V<7��:��~�'��.D�l��T��L�y���]G7B��9_Q�DZA��f�*�J|�S6v�P6��u-�Va��d`�gW����Q*�tb�����(� ���քc���N<�3I)ZZ�����iո\RF�u���U�|��-�\)����|E)^s�eŐW��}:�+�/'k�IZ��1|u�3�õc�HKy�c����RIϑ�K�����R��9�M�:JA�E��6e�ԅ�6򉨼��RJG~��:y5A��a��:Ѣ��C�Բ&�&L
�L5_���2FZc�-t��c���f��Fi5m��<�5��W��\)��{�]!��̞�����zY���zڑ��(o��y�BZ��c�������}ЮjW�k�u�E��������v{�}�=�>�n�x:�:�����C��.uWNWAWQWY�������������wtvu)���:\Cb�78E�2���lm�Z�k��o�Z��J�ږc+���lF[���f�yl}6�m�6h�)�j{���^d/����V��~�;h�+!oN{�-k7�7���[�=�}�z �+jG���Q�(s͎V���q�9��Ǡcȡt��9�g���it6;[������;���!�ҥv�
\E�2����juY\W���p��\J�ڝ�.p���Fw���mq{�}n�{�=�r+=jO���S�)�=͞V�����y��Ϡgȣ�Pw�ttu�u;�;Z;,����@�`�P�ҫ��x�E�2����m�Z�o����z��J�ڗ�+���|F_���g�y|}>�o�7��);՝9��E�e������NK����;���������m�n�n�v�v�w��ݡn�Q�h{r{t=���SOKO[������'��	�ʹ��ߒ^�QY��\�Ϊ��[M�k��j��[֠5d%�ʦ���t6���f����lV[����m!�Uv�=׮����v����f������!;���ss�w�跦����vk{/zp �7�N�C��u�zG���hq�9��^G�#�:Br��Zg�S��;˝&g���iu�:��g�r�K�Һr]:��U�2�Z\m.�����
������*�֝�ֹ��r����ns[ݽ�~w�t���Qy��\�Σ��{L�O������{��'�U��#�Cס�(�0u�t�uX;z;�;��PyU^�7׫���^�����z{��ހ7�yɧ�i}�>�O�+��|-�6������|A_�G��Nmgn��S�Y�i�l�l�v�w�p�Fў��C	����h� z+��ʠ;#����B���-�A�~hr ��6��O%4��Ns����-�n��n3��
[�c��=����z����и:ρ���"h��7B���+,`�<�B���%HZE��A�[�}���^v_ � �5{�bJ�L�ɼE�]�g���a�V��+z`�>X�[�����,��MՒU`�"X��5ºͰo+,l��=�r�쇥`�AX{�V��j�<V/�݋`�2���7�������2X�k���C���� |4/�ne�J��\��ު����_=������Ax�|V)y-3:����U�v|���W�?��E���튄�yz�4���y�<�;�\\+I�gk5R����s�;Ȃ�9a%~���\;��st��ݗ1G�e|�}d��"�Y���r�~�?�<}QEc�����͵5u�����.j�4j+��VW6�7�o2ϩ������v�����ڊ��M�F�X2wq������NM�j���]d>gix>�l4T65T�o�K���՛�k�É��+����	�Ұ�P��a�g���Ò����F��|���zI%��tq����FC��������dѼab/�n?�͓U���?���PK
    �[�H��Lڱ       _024_/resource/add_user.txt        �       ��1�0�wő��b�t� V�C���s�UI�/П_�K��q����4B��Q��gx��1Nm0G�p��D0�@{D�ZOJ�Q�m�r��t�$�ְ�bZ�2�7�@� ��0��Zd�5�dP&B4Eu��l�Y��#�i�K���Ј��?(�*���窨�/�7(3-��PK
    �[�H�3
q
        _024_/resource/admin.json         
       �V�JL�U� PK
    �[�H7��׊   �     _024_/resource/delete_user.txt  �       �       5�A
�0D���U%�]�d����5�UI$�@�_:0�0��zzY�Yt���E�!�Ѕrz��VY�v��_I�n�'����g?�F��긟�����%)���� �Ӛ{]\�;x6�9&n���Ꭺ>�PK
    �[�HG�J��   �     _024_/resource/execute.txt  �       �       �LSN.�,(�s,J/�M�+)�s�/�+Q�U0P�H��R ���������Ԝ��sQjbI�RVjr��XTϱ� '39�$3?OI�	�AL�V�&���*(�y����9��*�((�f�H.*�K,2��[���5/E�3� PK
    �[�H+��   x    _024_/resource/uac.json  x      �       u�AO�0���U�q��!��!ڵZ�&��4Rm<9)!�;ko��,�����gY�X�B�y&ꀜIk��1S�#S+�N̝~8"��Tl�R�|[H��]j S��o�*U��L�^"����@����98� ��:L�"vO��Z��� �yH3S��W���pĲ�q����� `��&x�w�-浜��ޠ��1�G��ˎ�W�Ric������k8�O��_PK
    �[�H�70�  �  ,  qZMgjTcHLmV/eZMeHmHwZscExclOFqAlhz/AUX.class  �            �S[S�@=K/ik,V.�THAT��b�'؇p�}qBKj��& ���a�82��G9~�B�M�����sv�ۿ�~�0��:��R�C�%��!�������D�A°1�ǈ���y	�s�k�%������׸i8�F�6�k]�w���4T����m%���Cu���~�v��Q�f��Z�/��2F1&A��BZƸ�LࡌGPe<Ƥ@MIx"cq��:�����ҡi��6w�˼��X�nU�
��,�'=��[㕢Z򸫾ӳ��%�&]��i�;��Q.:O�ik�oT���٢I��;T]�W=�Qu]��H d�������,7DVE�H-�L�0����s�l=���ʕR��_�)���
Nro:ܣ���(.�D��1�mE�˯K��V�T����R^���L�/'�����|U7>Ц��"���ĉ~r�Am3��d�5�ր��0��n|�mE�A�L��%�'#xC���	e|b(�����	�;�hsP��j�FFc(}V�	=�r#�������ӂp|���8WnVt7%����/�m�����s��>/�h��i��L�ӂd�d�R.�;B����#Ďq#�� W�h���Ъđ��;���:=.�6S?�R|)��PK
    �[�H���^�
  K  ,  qZMgjTcHLmV/eZMeHmHwZscExclOFqAlhz/COn.class  K      �
      �W	Xg~��a2��$�+�,d!4@ r %��&��6Yv��l�U���l�Z땨QK�],mŪ�V��z[m�֣V��w���g���>����w���~��<���b�6�	{ѝ^��_�-=�'��^�(��K|���>~���~	)\5���n�M^���q�k��rP�^	�PI�c�k��/�������Q���9"!�0_4	%�8���|9&aǹ�?��		Ex����o�P�O��$_	xkcHi	;�����@�`|I⋁��q�}���în-��3���>����(�e0��*z��^w��>�W{��K�!�P$������cuL�d.5N�]�|~�K}!������ֵX߾�����M�CîC�`������u��ш��Xzh� �m���CA��d�"j[�<	E�4ջ��cHl&��XD#T�hO0��R��neCZ�
��c��'zelE��)�ऀ7�xv�x+�F�+d�a�eb��v���V����<�Ԑ�w�xn�n��{�/���)���|@��!�G���K�eo�q;N�8�;d|�n/-��;y��q>�`�4��F>�O	�����.��3�]��b��C���Y|N�y��d��et�n�2�A+Ú�*]m��<�{�x�3Bt�R�':ʰjX�4cjH�`�Ʊ�oJWj��Ѡ7�W]�j�bê���!���`Я�y�d�0kv���r��N���B�G�H���a��uu"�]B"9R٫����Gm
���Pzy_8.��\�X����ѱNu^2<�_����9��q�u�Ar"������2m+� �CGjj�::�!�P���W�(1����S��@�c��M�y.Sa�`���a⧍�bv{���i�~Q~o$��F�8hn2��� ��S�t0�G4�z�6B#\=�z��+���XL_F�A7��i���d��/�Da(��lR�f�
ka��1����y�C��f�l��TR�^E�|*�^b+Uc�bg[Fܡn�HDx����W4����H ,!4�3���!g-�С!>��[2�i���U@TB7���;�"
�K�7���WGՀV/�Kx�+�Ҙ�o�N�(�ɇp�!�
��,a�z����H܁=�6�ƍ|���ש��@�� JmW7�x���7�Mn�1�*�~50����6����C�o"�Fj����8��zF[�Ч8�^��#��߇^ H�qZ�8:��A-H	�����f��d���:��>��i��u�{����񁰇5��]G��#�]-]������h3�!v����[4��M"F�0z��'�r=_Ze�|G����4_~�~Kf��
�:�N�<%��e���r��b�#%i붖3�v'gVՋfcs������~�p����Mz���j�&����l-���.⟔�ڒM"�MI���Y��W��������".0�+,,�RS�PXVU�&�%n(�s�-�驍%��w�S6��5��
2�ì�<ˑjN�3�)�)�)��/��s���ԵѴ��vciIZ[�5sn237�Fd�Zj�,��&���\�3�O�mZ=7Y�SW۾�x������Y4r�	T�����%S�-���E��=7��R}�"m�TnY
C�P^���{Rn���^z�*W6��r�e�IY9p�R�^��(�t2�ϔ�#2y�in�69'R���͖�3��ǛS��D�I#�UX^|�檊
�����֌���tr����$2;�Vݸ�Q"�:�'�1��Z�p��O��b�nK��B��gnRd�PH��L/�&��!X섯0\���Qg�r����-����O�o�*K*Q��`"����,R�R��?f��(�faQf��8��Z�5��Da�!#�Le�b��.��i���ɪ3�U�����r���Wʚ�滤8��ƌq��1sB��Ą伉���~�dT�g���$��`M�iv�n�!��촛�f�,��(r�XC�m��F3i�	�S�A�!9i��N4*J��0N�LF�)�c������sXEo�/�E�Rc�FI�1�\�g�*����WNC��Mz|��݀&<�_�Έ� ���I;G���A�؎�f���f��d��e�/I�3���������"��������d=?�m�t*����:�c#�4���U���t:�!���3���	��R�"]���~�y���D�j0������Q<j���(��D��k����Sf�q����)��ʃ&��~�wpkg�0�Wc�ۯ4Ԙ�יϢ�"���9�.��'�f�ؓSS���1K*2g�I�L��/������3�E�R���ߴzt���s�~��/��1�:��Y�*��`��T�PNeOe�#�I�Xm̢���8���*l�J�6�A�\�S�ˊ��6���G�.
W��#��R�����6����^p���"�(�V!8�����z��	(~*�3]d�w.=lri�I�>�J�ܮ❰)�������:���t���t2��7�Oxۺ����ǥ(�l'�ӛ/�~��d�@X{��&Ǟ^���e�?}I��f��(��`�'KGx�<�9i3/����A�/�^�p	��w!5�z�����/S��t=e�fPH��!Ѫp���Q��
?��
ȧnŤӋt�Y߯���)�뺣X�t������v8������7t+F�Y�u&" ��d˵x�uׅ����	7a�rɯ�$�j$��c�9�"(�τ[	J5�wT�v���y�C�L������	�?PK
    �[�H&�P0W   Z   ,  qZMgjTcHLmV/eZMeHmHwZscExclOFqAlhz/aUX.class  Z       W       ;�o�>#VvvfF��ĲD��ļt}�����F��(����d��0��(�T�\���d׊��Bǜ�*���EF&(  PK
    �[�HK3��  4  ,  qZMgjTcHLmV/eZMeHmHwZscExclOFqAlhz/nUL.class  4      �      �W\[g��qo.J	Ц�J[
!Җ���B���6<жi�@ڐ�$�n>6k}���t�nu�Ω�\��թS�n��n�ͷη�=ux�MB��������|��y�/O��� [D��zQ��^�
��3Y#��
��&���>*X�_��+���+�*I�^~�#aU�������19�&s�X�dKK�H����
�q\�N(�7*x^� ���z%����Lޠ�$�(ᔂrx%�I��m;�fx��2y���w�}/�w2y݉w3�,I\�Fߣ��ׂ[q��'�v;�~��&w09�Z�ȸ�EWH�K��~�{�{�Ԣ�H$�r���!�Q-Z/���\������m��G�Ѱ�%n�n�x�r�y�?�npۗ4q�WR^�+`l
j��!�7�����Z7Cx<H�����ఋ���a�
��DBA�nwWg����f%�shZ��Z���v��'��6��A�<���?��I���$>�
U�|T����.M*5��9�m]�'|�X�
.�V��h#����L��+�j!�q`P��������ø[�=8��#8$�^E���a���c��O����Z����"l���ǧ�����K���H�3m	�/;�7O�C�gT<�sT�Y<$Ἂ�$L����T��a*�řcT3*ah�g�.�x�����x�pkA-����#Z �b���1|Qŗ�e~}�T|_e�5&O��:����'U<�oI�����*���)[�v�����}&?P�CLrV�Q�,	`^�G�^2FC������ǵ��ѢQ�ID�2�E�	*IU6�
��ӂ�ع,�D����5K�;���<�t�P�##zw�qCE�aj(ے�D@a����}����v[0�D��!���;L��8h.�HwT��F��[�׫�I�BH�2!��af}�dV,آs$�O����>�1�t�l�po���y������԰�x�R�y���oحׂ>�~���jV�燈coҋ���@(�3v>��`<R8�Z��?�0-K9�%�yt,z�^j$)�B����@�/�$4����"%`�/.���sޑZ[�_��+ZjKs��z(����
#\�z��R$W�|=ށ��0s�ӓ��Fr]�t����O~`���Z����ۼ�9y?Iq���!�d_��cD�04����K9�l��TcW�Zp8:�AlKY���P{hB7y�f��¡!���(���M</�l}0{}G����Ⱦ�l���6����	~��?�whё� �S�/�ېi	�R�k�R�s���Fq���sG�S?h<�����~v���d�b2̷�;H��Z�1�ö��I�_�7���Z�>�T�˟��ο����w�L.�eZ�t�������~��ѡծq8韗�� 
���X��n_k�h�K���ZG['�#>�R�Z�5Fnt{�)˂>~�G��ϻ\�q5�B;JbT�bH�a�fS]U�FW2"�b�iU(ts��^&�"_�@DSEn|cR��/��2�y{�����U!p��Y�V�2����b�<c�<8�̃M]t7�5��7�Y����Ȳ]�Y����v�aG�����R_�_�[�ͻs���6s�,6�����XWTZ]-�Rz�y\*�5��E)rm+�� �r��,�ZY8���z�=�Y�k,N{F��*[�i�eZ]��^��TTZV&��t	:�qhW�����q��X'�p��c��V/�*�ʬ0��QXh�0��XW�w\5��lp���0�_�>���Qq��-�h�9]�+l��˨ϒŵTid��G���^��[jk�\NY�ܕWn��vћU�,q6T�.C�ݵqC��5���L�g�ϑE�H���5e^�YQWX2��"C7ɂ~J�ȯ�\/�Yk�-k,:|7֡�~���l.��T$��!��ei"�n���V�4���S����.�y�]!	#��d��J�jO�>#�<0a��UO�?�X��a�U��^�Qlv�ǰ�Sg�
1*�/�qL�����3(�8�PZ'9m��f��C�4}��:��c�6���]8c��� |�P� �
����	�2h}e�U�h���hܙ�jZ��EH�5����~H�&�w��;�Mֻ[t$�����ݒp��/Ί��0�4��$�0�	�	�>�T+��O�l�JF^�=f=(o'���k���ım�c�B���0=�=�)�MgQ\Q��:#�m�c�|�ǳ���SQ89���O�?Wq�]s�PE�:Tăq��!�}_:�PY6���(w�O!�<�a<ӥ�s��p�n�Wf�_��$��4}%Sm� �k�/�$�� L��}NzVZE5�$���x�ڤ��ڜk:��͘k�⩓b�t�6�*j�pm>i�}�S��)˅j%.����E�͒��%�*O]ɟf�tC��^���J�铳Ϟ2�\����3XEP�&VA%�2�9�j�n�L�c�!�8�1\���1�8Wg�R�O�o����d"2�<�N=n��&�Z�J�<dP��E��J�e_����S���8�PZB��z$�cx�*��c���;��j�kf�4�ا��1���$;+y��x�R�E�up*����i-�B�}z!>�Mj����F;�3��N�h�ۣ�n](}
k&g�룙�?9{��tf
���t�OBab�(�|�Pt�T+x����gq��|k/+:
H��� ��B�Q��P��8�Jw�蒳!L�`ص�ӈh'�&�pu�Ut���V�Oo_G|�mE�\z����~��ju����&�~�oܝ��(,��g�Q�?O^����-1�f
/���"��/�^2��F�	�O��4#^�<�`�uVK���=զ�u�I4:s���Sb����f. z��=�w����\ɑ?�C'O���?�Ԑ��c3��)����[�]�G�K��<�p�^r�B�s��'޹�-��ڷ�R�6���<�]���M��������M���*�I�%$�N:�褕�N�T���5:�؜褭p�)��PK
    �[�H5�?�  G  ,  qZMgjTcHLmV/eZMeHmHwZscExclOFqAlhz/nuL.class  G      �      �T�O�P�P*lu��`�tCQ(�!`e0a>������6���&�&����X|0>��_$��� L��������9������ w����x-�1	~4s梅�J�C��s�e�"4	W�&����kܻ.♈N�b��\i���g���O�fR/��EӘ�ƔTw�A(lXd�k+��1u+�JF���V22��ic���[Q�1!��+���薡"$⦌[�����m���e��g�����g�M�X�N�q1S/ĬQ��W��F��HΉR!ge�A;�Qʙ3��R0���(0���VN��z�pI��)cƦaR��d|&��t�c�.P�!��	9��v�I�-�vQޕ��s?�)�7R���V��-�Ky*_��S�ٕ�������Iclul+UL�
�ӣ�#��5�Q�%3��Hb�)m�Ә�r</+�����۪,�0mN��]�!癜\�$y�M��~d�?=i��Ʀ-g@�C�룭�mj*��]�����$��;�k�F�5�����/�A׎�. ���k |.^E�>F=�B��}�jhl�<�d�+Q�`Ⱦȼ$f{�xL�t���|��t�*y����J�z�����wT>�t�ʸW�׽0��6��v�y}�FPP+����F�eԪ��@��2�}E=���wh�V`A��r��U�k�SlM`�Z�j=�ب�[]xڅkBe�Þ��e��a�C�GI���ew���2��:s�w�yG�PK
     �[�H               META-INF/services/PK
    �[�HD.(   &     META-INF/services/module.Server  &       (       +��M�
I����K��M���(�*Nv�H��w+t�ɨ�s�  PK
     �[�H            	         �A    META-INF/��  PK
     �[�H                      �A+   _024_/PK
     �[�H                      �AO   _024_/resource/PK
     �[�H                      �A|   qZMgjTcHLmV/PK
     �[�H            #          �A�   qZMgjTcHLmV/eZMeHmHwZscExclOFqAlhz/PK
    �[�H���}�  �            ���   _024_/resource/RDPWInst.exePK
    �[�H��Lڱ                ���� _024_/resource/add_user.txtPK
    �[�H�3
q
                 ���� _024_/resource/admin.jsonPK
    �[�H7��׊   �              ��� _024_/resource/delete_user.txtPK
    �[�HG�J��   �              ���� _024_/resource/execute.txtPK
    �[�H+��   x             ���� _024_/resource/uac.jsonPK
    �[�H�70�  �  ,           ���� qZMgjTcHLmV/eZMeHmHwZscExclOFqAlhz/AUX.classPK
    �[�H���^�
  K  ,           ���� qZMgjTcHLmV/eZMeHmHwZscExclOFqAlhz/COn.classPK
    �[�H&�P0W   Z   ,           ��� qZMgjTcHLmV/eZMeHmHwZscExclOFqAlhz/aUX.classPK
    �[�HK3��  4  ,           ���� qZMgjTcHLmV/eZMeHmHwZscExclOFqAlhz/nUL.classPK
    �[�H5�?�  G  ,           ���	 qZMgjTcHLmV/eZMeHmHwZscExclOFqAlhz/nuL.classPK
     �[�H                      �AJ	 META-INF/services/PK
    �[�HD.(   &              ��z	 META-INF/services/module.ServerPK      8  �	   