PK
     	g�H            	  META-INF/��  PK
     	g�H               hERVpYPtfIqNRTl/PK
     	g�H            %   hERVpYPtfIqNRTl/qHYgYZuSZInssdeYNkyW/PK
    	g�H��I�E  -  .  hERVpYPtfIqNRTl/qHYgYZuSZInssdeYNkyW/AUX.class  -      E      ���N�P��j*T�7qW ��[��A�$b��J)XlZ(Մwr�BM\� >�qZ�QW,�̽s�7��y�x}�����JC�BY,Jؖ�H����	ɚ߳	��o��n��u�v�dZ�=
	9�14�M��ǵ��!��$CB^�e��XtMo��u���M��|B; $ԢN�K��39r��`[x���	���qK�a�>n�ڮ6>5F��S�&��m4o�WZ�����^^G�I����(�2
X%���./D�,H�E0�IP��n�����8�KF�	��_���5��m�;�id��
��%���x���?�Ȩ�>PK
    	g�H,IwQ  A
  .  hERVpYPtfIqNRTl/qHYgYZuSZInssdeYNkyW/AUx.class  A
      Q      �V�Wg�}�f2��T↸�$@��J5�Y� ��d�1�	b7�Xk�}�[[��GBO�i�ԇ�=}�9}�s��f �}������~w��??��>|'�{�؎79x���9x͏V�/!�6{%��'���H��NtJ��~I���88 ࠄn��8'���ts����W@����pDB��r,����c�p�!�3��H��D6�ƭ��M�1�C��̧��U����G���E2�^#kX����Uo��ʚ	�g�~3�� �d"s<�7#}�w��%��{!�褚�-�PȨ�xO�L��y0���:���V�h�k=q����#�eK+�����6\':�-�,1*#U���!h�e��I����(�<J�S�)��V����A��J1T������bY܄΢�I�yc�00.�22�"+�DN�9��⤹�<C�r���E8/c�������L�9�0��U�#eʡ⬙*ft5��'t�SQ��u �������5}�ukӝoP>I�e����̼���Y*��[ݺ���4�e���괾�oT%|k��^H)/�*�Т�R��Y:��JY��&�!R>��/���v�i.�-RU,R)0�)G�|U��v�/���Yj}ˊ4�f�;��yg5JYӫ��Kw"�ť�I�*��c�+�[\c��tC�[˙_�r�3L[�k�f���l7ɌY��%�^���lA�S\w+���������O�R2F��&=τi��d�e�;�3�u�xN;b����Ȩ�iim��e������0�v��;��Y�~#���è"�J�Fy�	+9&��!�A�����x���hdPV䨯�Y�U��Rj��x��h�n����x��L82�Z���w���Ơ#�.�W����p��|Xp�O(�z��~�u���{+	��Z�o�VQ�!�*q����r}�=U�!@'�l���}^�4\U�<�`h؟�}]Eg7�_D�שp� �Q�u{�������V�@�E�+g�:�E�6�5Z�x�{<泯B���D	ԇDEn�[B5Q5�R�����D�������h-�~9ϭ-!�(~��؈-�n�Bdu]	�K�0���-�Ƒ��5����ouZ�7C�x�ݏ"��884���݂�XWQ�y�A��-�n�>��+�M%l�r�N���&z��~"dN\�7*��?O��63�E�.Vǚ����]l��J厲N�E�V�f�<	?ov�o��E�&Y���a��2��9�{�A;����b/�@.c���@�@c �&�p� R�#��m�i��s]Sd8��n�̀M�5�4<��N-D��n�7��]�y!��H'�.�1��mcW(�/PK
    	g�H)�  �  .  hERVpYPtfIqNRTl/qHYgYZuSZInssdeYNkyW/AuX.class  �      �      �U�SU�n��n��д�FS[,�� ��B1A)�`H(���n,]�a�Q���;�q��f�iG�3>�G���T�a�=������=s��?���=!p��wpEĈ�"Fe�1̍We��(���6ε��84ɷ׸H�x�s1.⺈/D�`�䶵o��a�
�m���N��[׾�0������0\��0�� �Y�:C0gU5sU��b�%.�v�A2�q��e�R�-��Z,�h���Q����0��o���]gm[��Qp
&q��0��R�>�V����1��#|̵Y�t�9.n)����ⶂ,"�Um����U��Q<��Z��*թ5��q�h9+���Fc'8�tg�Ҳ̶�/kN�XGc��RǍF-�Z���A����U)˭�1���f���ި�^��9�t���ɳc�����W�-غ^lTFC���r�W�~�P��<��o��htϓ�Gr�W�|���3�}g��9�y�V͹o�l����v)�K�El��e�2�Pf�[�B$r���զ��lew�+%3�s[�����z��jm�j�����l�L$�Fw�F1?V�R��S�+Xâ������8�G�t�|�<-��d�GZ#���7	w��		_�Ґ@���#c�t����ԕ~	DG��Oݼ�JJ���%'�?�``���=�l0�ɑ�dx0��|�?�����Gͽ؃w��	|�15-�O���ZV'�!�O�B���~B�jZ
~��\Xt!��C>X����9,7����\(��:����?K�%g����_?���urT��b ,��+I��TaXp1��l�t��C��K����@�e8��.��Oq��_��xq��ܒ�!��Eܡ���%\�����9.�������"�=`�x�"M~�l�����~A^��D|�	�cxv���	�g��� �!Z�7PK
    	g�H�g�4�  l  .  hERVpYPtfIqNRTl/qHYgYZuSZInssdeYNkyW/Aux.class  l      �      �R]OA=�ݶ�����v�l�/CHl��b���cYXf`?���4i�h��G�lIM���Ù�;�cr�����'�gxZE5ne��0��f��ᶅ��:��2�Q��a�itJ��+j-�Ó���bSCE�U%�3�'�f�a�i���	�b.{��%��`(+�&��FS6fq���m��=][�qSWU7����D$�ɣ�������w�)���d/�!ٛ*�
��m����*<ě-x��������-�8"��\�u��=u#�4�	%�8��Yp�x�G�3������Q�6��<nol���l��VS�iW탏���)��y��X�"�3���q\*e�KU������2c�ƭ�J�Ll�[���n�g`_�f����� 	�a�\�|.0kO�a���*�#���>���D�}L��Qr�0�`~�5�Zz\z,\�"d�PK
    	g�Hbs���  T  .  hERVpYPtfIqNRTl/qHYgYZuSZInssdeYNkyW/CON.class  T      �      �V�_W�>r�V� ���'Mb0��(�b�D���.ɂ�%�b�}ߵ�m��Z��b!P�֞?������v^���vޛ{�̼y����n ��o�Д�����O9���+lŶ|4c�-h�fA>����;-(�.�9Ⱡ��XP�&:8�+�kA)7��trt��.�����@�=��h�K�q��rpH�����#|'�,�_���֎c��V�Ƞۯ��F�a(L3{gXU�hn
G��6�:��:wR<����6-�p�ZPV��XX�W��0�\RuG���n��ï�+:�_rˠ����}	=��ɛ"{�؞�Lni�t�kw���M�4ff�����y[%�G� E� ��1�%�b(�#b	hs-!�an=Fq���8t.�`(�q	#8��h&��UhM�Ր�p��C�#t��NᴄGqZ@H�cx\���"Oq�������j������y	/�E	/�e	�p钬�Ƿc4�D��a(�^:�Y�t��LO�v�ԏ�:��a��J��ۯ�FJ܂x*�;堮�N2,���2T�ew���t2]IS�r��Ǒ�q#�:T�+�E������h��=�pP�Uv�r��v���b�=7�*$C32O5�agv��s2����g�}I�~�3rsi���T��t�l�seՑk��hT���祑iy�Xײ��s���t�1%B�Ĕ�*�Ue��׈�i3}QzXuǔAe��)���7'4��B �^yH�]����Xp"֕��)�� ��4�&�t[��9�/5��d?��	oJ�x�xR�AU�+���U\���2� �+1����?5�po�W�-���j���qD�R�j2e<GwtuG���g�۵_u���>O$)��=�6��fRf�v�~�d���̌Tm6 �C>�΢Z�;pKx�$��j��y�|E��h����K��ߺ�)�+J�^WV_�P"���j���5+�"�R󶄚�Ʋ-V��ܰu�õr���t�2S�_W��]#ڐ����As��|i���f�>�%VU�$37ɨݽ�.��a]�6UVU�#�/XA/.��1Yy� Z)_��lf�L�D^��ւя���2`�8�I��Ϝg����q��!	�&�c�7	�4
k��&�`�4
�~�$���(L�h0Z���k��t��h���-�[�'S�� �4JI��U�Y'��Dyo[�#V6N��RmI,&�t�K�ߓ��"�\j���),��&2�#�lW?��be��+13gNb�+`�݊$V&�j�S�Ěs��u�@�����k3��$�uB�.��fv�D��R!�{���W��L�]I8�c�h�`=p�n#�P:�h�9�*Y>�&�cU��:䡙U�cl����F�I��y*���ӟ�l��mD>�b�A��E4B��ǆtqq�<�h�X���:�\�I�	�M�0�Lc�MGUK��~��s)�-卥vh���qo���"5��PK
    	g�H��p_  U  .  hERVpYPtfIqNRTl/qHYgYZuSZInssdeYNkyW/COn.class  U      _      ���N�P���R�T���4q�11����A�ݡ,6-7Mx���5q��Pơ��X��93�?9g>��? #�d�*c�T"%D%��'�c�N	���2	Ѣk�&�h�fu*\$���T�+�f�ڥe��t����J�26$l*�!�`q��U���h�f�4�):���?����!lϭC�`�pO�N�-��j2Ż�J��_�څ~�R������7��3�L�t?�ky����8P� A8J-�"]S��6!�h$yHA�@jd
��|*�W��mț�>�rFϾ���{�Af��d��]���1�2��f|"�
�2������>���v�_�ۭp�PK
    	g�H˿4��    .  hERVpYPtfIqNRTl/qHYgYZuSZInssdeYNkyW/Con.class        �      �V�WU�\�1���ce�,-�ea�P��G�� ,�ca��aw���U�,#z��J�,�A��]<m�:�N?�CAK���` `��{�~ߏ��ޙ?����j� �7����<T�`�Η9Y-��9g���D�8/���3wb���Y˗�<,��	�:Ω��nN�ỽ|���<�C��y"���/4���>p���uD9�TizU���1�S�X��4U�g���P�HROT�t���:ķ����0��Q���V=��Ê�)�q��/y�����*Y���(\��0�	b;wk	��˰���͏g%-#�Q�P�f	-8,�mBhpD�c�`X��#nQ&�]T��,%t#��=|� ����%<��=!�I�Hx
��A�Q��ۛ̚ND�1Sө��7�$������(�{H�ej�!���.X
Yf}�R!��"�c��<�T�nLX��1�`���U%��!)��Z��ML2���GS5�˗��-&ej�*�SdjO��P��_f������1�P(K+k!�X&���FS��B�(_���/�miN+�_.�������4����Ԩ����=����WC�0����9���ϏM��G�F⸡�jVr��#O%)��w&�?������H��~�~��j�Zs�D�vJ�p��/�_ԂyQS\Uf��ah�x$kܦ��z��*!ʩ�.�"t���b;A@��C2kn ̥4�N-�T�H�ͫ9[�r)��q����`����Ӌ�p�F�3"N�$E�+FE����%<��\�<����X�W��3�o�%��(�e�ǐ��(fL7�2��B�)��g�u��#<&1c�㡎�x��!yH�Ku�5'�ɨ*��N��KА0�F��h6��%��/��p?����e�@«�J��*�P*�Z�F~C�N5Ҿj��ի6t������R>��r��[tx�f}��V�нc�l�X[�ÅO	��Z_��T՛�b��*���4�"�s_.�!fII]�G��-�^r�=�� =��ı�ӵ� �ַ� l�̫�Uf���o ���Z7��^�8��,^.Α;f�� �9�eYw�}z���g���u�x>��WҰ��.�����,�U���}r�L�]i��ixz*29g���@��ڛȭ�e�'� _y>#/�ܛFAb����T޺�R�sܪq�H(�^�U(>�W��s�[׹=_��������=_Α�4����!��D~;G������s�Q�����g�؂V�K&�A����N�ހ|��4J��D�4�V��<l++Žs��oZ�.d�x��#�9���7޵vQ��3��'	򳨀��Y�pa!w���9���G���r1��PG���i��`| �Fˉ4&�4��G�I���h3 ��3���=ڿ;T#�����=5��:�4�^{�x�͒�I������<�]|	$��
��EҜʙ�.!�ױ����o���3x���#(ѓ�b^�'�PK
    	g�H�m9ΐ  �  .  hERVpYPtfIqNRTl/qHYgYZuSZInssdeYNkyW/NUL.class  �      �      �R]OA=�--��*� ���DmLc��e�.e��.�.D�����sZM���zg��"��a�=3s眹w��ϯg 2xE�#��'�9�8d���a#Q�>��(��(����a�|{,��0��W��zڴ��M��1��^�I�{�YۡE�g͛5�[`�K\L9�rq?�,2HK����nu�Է,c�CO����a"YTЏ�0n)��;
�b��$��N�+ƞg�5IL0��[���o3([0D,��8u��Ϳ��4�g�cT<�9��Q�_��ʽXL�tW���X�v�!��Iג���{�e�UWv�׊{�+���/�mX��ڎV>X/�k��mh�G�t��
:�*4�h�$Tѽ�.��{y������Y)x��T�*�D��gS�aH\�j�M%g���ѯ�b���H�~$k?�<R�8� ��l!�G�!���	�'�H�Stj�M(��j���!��]ĮNai�gr����� �\r|�a����.�%�"R/�XG�q%H&!�	��-!�lC��&B��ق(i�ڜ4��ɸ�Ѳra.?(��1�%�E>I,.��!�]��JȶJ�89�@��o9�C2oBJ-ǥ)�<���5 4 6 5 ��g)���W��>���l���ehM��=��PK
    	g�H���x�  R  .  hERVpYPtfIqNRTl/qHYgYZuSZInssdeYNkyW/NUl.class  R      �      �R�n�@=�4q6�)whJ
u��By,��RUm��� [�q��:R>�ϨT��������̙�93��o�?���p̛8_���8�{�jzQ�%������X3q�a��Z��BE�
�u����!ò5N2��N��_?���6���P�G�Z2Vr/�t�T	C&��V��1�2�}[�`����.���q�j�'���ؓ]��	���r��E�v����|K�l�&�V��|�ɪs�D��B/V�؈�y�̸��D�_L�Qԇ��s�(���Z�G��E1s�����ց���6��@>s|�3��l��~�so�m���Rl�>ɱ�"��"����X�=�d�lI�dmm)�pe�� �
Y�G�1�>"��}����1�/Ӱ9B���G�&G�BOL�Ǌ�M}i[q�g�]�![����/�������Ml5e��
��i�W�\��A�r���PK
    	g�H���	  3  .  hERVpYPtfIqNRTl/qHYgYZuSZInssdeYNkyW/NuL.class  3      	      �QMOQ=�3��a��P�~!�:�'a�BЍ��6M˔��>���T�S��	��u��&���C꽥IE6.޹�s�}�ǯoC �ptLc!��:����5�`���U�k�S������+�����M����#��yvxa�ً#?lm���NS
�J��T���Ya�����BB�ɳ��~��tp>g �9��$�f�Ģ�[X2p��e�d'-+�HzM�i��ďd#�D'��u�t�wc���Ń{7e c�!Ӓ��pTM�f��ڄ$�5�����*���V߸;���qy�8��ݖ[��շ�n�)��듚S-t�x�b����*`	�π��J���>���h*�00o �#a��}�@���<d	�&E,&E�٘%M�D̍��Q� ����P�&t��HD�&x�1�#�������I�/���7U��V��pCUT�jC˫��p-�������UHR�S�e��d��i"�����g{��d��Ԕf�}�+��4���C֦8	�PK
    	g�HQ�ѭ�  �  .  hERVpYPtfIqNRTl/qHYgYZuSZInssdeYNkyW/Nul.class  �      �      �TKS�P�n�&�-��XD|AZ�ъ��*����Gk���FB*i����\����hq�q�?J<�� �qܜ{r��}��s���__��c6 Z��8��8'aFB��l��JW͊:kZ��8nڦ;�Ц�"!Q)�JA�2�c�˖���ש�d�HF�YB��vt0�e,�.�e�Ћ�5״Ԓa�YP�j6߁Ar����u�]ǴKӵ�Ñ���qd��k^��� ����Z2�yW/�.8z����H>���4ck�����N3�DNXz���׈۩DR�����c�CSB �q�!��h�j !\k���p˕"�S� �8w�NǴ���2Ĕ�)*'B�Q}D��C�[ib2b\7���kv�-�_R�-�>rnM��;#N酲�LQ���$d��G�3��|���(�Ѕ8�ݓ!~�N	z���M�g�2/�g�Jr==�`��O������v�Z4��ꛬ��Y�b:UR��BY�C����i����9�</=�3��৯AZ���Gx>Û��� +7Lc
������-�n�"��[���z�x��+;��Ԁ�%s�Uk�P[��X���㾯%@����KB1?����!��M���F�w����hx�����l��v1�c!)>�P�go���o"���}�Zl����M=M��/$��S^xhEs;`��9�D!<��ľ7M�$��PK
    	g�H R�  �  .  hERVpYPtfIqNRTl/qHYgYZuSZInssdeYNkyW/aUx.class  �      �      �QMO�@};�C�_��������RE��h�s�8��qpL?���^�p�RU��QU��T-p�;3o�{��������(�ǌ�,��5kࡁG&<7�bు'��ײ/�u�V,�	�F��	3��A[DRt/��~����b�X|��M�k7�R�0u"��$��:��cߋ��"����b��3���H�3��2����	�m'¬�Nc8jn�aR�ʈat��� ��	B�qTk��N|P?i���d�=t;���z8��n����#ޝ񫲞��#z|��P��^�2�A���i6%r�,��@�αU�F�f��gLs�]���0���������$����Uղt���ЛJ�����$�j*r�[V����-��^��s��IyI�I�^��t�Ijb� ��~�)L��O>�+W~"[�s���[�\*� PK
    	g�H���o  �  .  hERVpYPtfIqNRTl/qHYgYZuSZInssdeYNkyW/cON.class  �      o      �V�SU��$d�eK!m ��J��j1�jI�M	B7ԏ%,aa�Ɇ��Ѫ��t�g|P���5鈣/G�/�7ߜ>���� %����s����{�g���?��y|*��z�G��sN�/xQ�}^�A?�^� ��x��.pΫ�zM��q�EN�)·n&"����"�=�׽����xC@���ry>o��d"9=����y����PUD��+b�h���V�	5��ӆ6�'g�`�������ʺ%醖,�ق=f�4u��y1�� C�$I[�[7��zVN�٘Y����vnm�m�X,]MkY[�L��q���!�`�T"�{�%���A��HHHb���dh:@��GZ;ǌI�[�%L`R�U�0pP%(HI��S;�Ix�Hx�IP��*90- -a����$蠋8yhf��rC53����ah���\�l��G���ӡ���-�@�~�d5 VCho�p^`�Wyq\$�jo��<�xj��%=G![Ju�bӆ�׶��AFԜfҡ����-p�"��3UP�H���ք�;�UԬ�t����8����]�����;5R>�ae2dQ�Ӫ嶂ݡ���*�;�W�-k5���Dt4����ǐ���Ё�CSCef��B�pC�>�f��Rטf��EG'�ʈ=[J����e%��
c�����hJbamRN'�ը4���"
�-��i�Ѡ7J�et,�S��iz𷽈6��yK�'�R`t����}|���{�J�V����r�3<�0<M?��Zw��&�J�8|�܅Q�����M���z���J�Q	�~�tQ��^�i�џ��8�p#=E�q���Kh�\p)W����=E��>�A�o����'�~��c��p�E߶�yo��"7�}�"�w��N0rѲ��?qa/����JiP$q���D|���5�� �6N�~�o���>�_�{kϜ��۸W^�!_Y�:41'Q��p���P�/K���S�A&��8�<z��7��.S���3�"�>�
e��-�,Q��+e^7��n��˴��.\���u��K���'�@m�&:�a��#K�"�H;�N�D�G�I� ��+U����q7��z�[e����h�PK
    	g�H�M���    .  hERVpYPtfIqNRTl/qHYgYZuSZInssdeYNkyW/cOn.class        �      ���O�Pǿg��V
t�SQ�[���11��K ��'��ʺb2�^|���Q��Ҁ����{���~�='���\����T�ԐGQC���@Ō��W*�(��Ȟ����A�#L7W�-J��f�T7�r"B>͛�c�U�2�������u��]���"���;�cύ��+��t<��xJ������!�$�i$}{=�PDAHP�r�0.2����,�ڄB�H3 ���g���8��k�8��A�������{��i�~h�{�A�s�?��c��˹"r���;1H^���ݮ��1�I��`��<�<�}�Q�a�E�&`�:Ι�`�b�B���c�,�x�9�%� ēZJ�U�2��c� ]"���*]߰=S�i���yn"�?��5��F��72Y�����$�6D!밦X�eo+[��1�z��m*���nSqPK
    	g�H�r���    .  hERVpYPtfIqNRTl/qHYgYZuSZInssdeYNkyW/coN.class        �      �W	xW��d{���q�\���HG�H��DI�:������)���ֲlY���@J9J�U�H�J9�t�W��R
�$�(w��g9�M�̼��C����{���=�3oW��� �6;т�r�~,�n�B/!p��x����x����(E�0����X\���.��`T�D,G�U��E�1��pD�.�D���u��*7�sC�oyT)�8ʱ	�q�R��/n�����_��p�R/�+��ܜ���f����9 �_���{��?�
�Rī�j'n�k8v����hGX��x���1���<�K*�O����@�Q���-�/��:+�3e���CS�Qb7�;��<7!'c>"Ɠ1"��'��U=�(_�m�p7�3T��Q��V#r�_���������%�Z*��3��zi�'�mY@�b�a]M�����}��y��&d]�F��JF�&"ʘW�<[ϡ�����E4	Atx��7�������5Ű��l�R�DT��Q���&�Y�[�V	w�.o��v�C�	n�n	��]ޅw3��"�%r�a��{�^��#�}��ؽ���9��>�J��>���O�G�Ǐ��\�|��OI�D����l�Nr�O���b����X�)!��=-�3�_@V�g�9	����<� ��!j��LAKtCu$����F�h*��zm\��bT.��S�B��{�o�%�\S��zsE3��Zp��S����A�G������S3��L-Y=�H�C4�e��A�u����KG4;5T���Q�e���Q_0�VP�!kda�%K�'W_�9�D�j��&9Y&�0��L�uC��:�Y�(FK4�):�W2�3�CY/-Eϛ8��s�]*O�|P1�,�����w����U\ Z�H*ҷ���H4��[�K��l�ɣJ�Z��a^��~v�$A2Fj/e����Q � �ʌ�������]�B�q%AO���������+!C�v"0�zʊ\��t�G�+�J�~�F����(�*��o�1��lUG�dM6T��/�Q��p�-����Y$|�/1�⃔�J��W�Q�NPe�:���Lfh
�u�������#��ބ�ȁP,N��;��UB��c����12�"���l��0�8-n�J�+6��7�*+�i��[�p�/p1�	*�Y���*������<_£0x*-P��r�D�V;+�����R�R�+m�<-z<��.B��Z+/VK� �R����+w�r9�Gj���_p�fhO��X�c����k�z'��Aj�D�v��f����zm�{��j�Co��j[�
���dX��1���-�������]�����کE-	'��A0t�i3�g��e��4L��%���!DF���yU۳p���PS�S�g!���~NןN�	�ė]��ZN�k�ZkB2���Lԝ����)�7Yؒ�+=��Ц���w��RZv��=i��{hiɴ�Ӻ�XDg���u��h=����g������,�ś�*���[)�ա,ք������9�5qIzz(�u����,=������[��O��X=�1qŉ�Y�����5�Ll0��c3h
���Ӷ,�TK���X���lYے�=Q��_������Z���s����+z]�,l�;��H����ܱ,��<�jdpe��4�#�8/�(n���-2��뚞�nbY�<���mbO:�<�{8���p���ӹ��d��bb�i��ĵl���I���;���fm�6�X�~\3Ӝ7QcR�x��X�ob�x��<NS�p�=�o�6vY�6�P��؉�XX.|�#�,������5<A�4��$�`O�?�Ӷh� �(�93E]���}�榰wSS86��S���&k���c���h�X/ͦ���Ѵ�i��[i���?��Ɂ��5�T��9�sq�2��PK
    	g�H/K�9	  1  .  hERVpYPtfIqNRTl/qHYgYZuSZInssdeYNkyW/con.class  1      9	      �Wy|���,i���Fƛ�@�l��r
��Q#�� dS���ز�d��$Mڄ�9Z��=Җ���)�}�w�6��#�6	GCgf�C�r~�}o޼ys|3o��>`���B܍f!I�eT&N	;d8�+�O�q�$x��d��<JJ�)cRL�L��I��dyj0�1��v�ȸ{�1��Eo��-x=�[%�&�2�`���F	��X�f,�nҳ�G��K��ɛ$�Y�[p'�����%�#�jv�,�6&�e��29�����c�N�����������ݬh@��x� ���{�>�_2>�J����-���gө���M�M=�z�h�j��vk���H�Yf9�K��*�:o�M�[�-�.Pݖ�i�-Z&��$�N&��t&ҁu���T��,0��'��0B����adtm'�͟Xk2�5��6�)gK�����ʭ{c���H����NNj�� �&R�MS9l�T��ʋ�^n�roQoJ��%&�7�n�֔�����
*2�Q/+	�9�ٲ��ęfh�D�J��	��u�\*^,qI�D��
ڰ]�f�F�8F���i2˛>"0�%������a|\�'�]�'�)�X%������!��aGpT���q&��8�R'��a�(x�Wp
�*��(ᐂ/����*��#P[>1
����{X��9�H������
���
�Pi�%|K������|���x���{�?��>��G�1�%/±{G���Ϙ��
~�_J���_+�~+�w
~�?(�#�T������ga��"��Gvĩ�&�zF3�bN����7�������j۱'�0��H4�X�K��ĩ4���m^��x�T.or&�|�U%]�zucMO6��z�_孿�1���8�x���ҖIڵx�#�{%�Z�ȮMdh�ΰ�Ik��/���bS�/)�&�9���Ж>-ӡ���X��~Y�䬡e�l$a�MMrĝ��d�B���*r%&r_;�L��ԧe��^��=e�J�<q7)�r��*O��2=��-�Tk��z���/g��X�6�W��6f�l�l켚2�E*²��ie��v�#몋2�/㸞Թ�I`�tb�ݕՍ6}��䂰�ř�S��K~�*]˔�f��٨�ZFO�k���N}�Y1-�3]�h��� �Բ��>fe(���%m��3����K�w��ަ�[�Vp��Ѻ���u�b�_��h�N+�?u������]|Ye�Z��7&	��'���K�_��ޓ�����?�T�w���$�I�;��MGL3b�0A�����o�n6v�v��;��]룽Ѯ\GW(����hx`(�Y�����C�F+�HR+(ς> 9 (�b��~���63�baU�/�Z����@QǇsɋmI�.V4Ƣ�e�V-�D%�vg��fu�R��A��t*�K�"O���l��o�_	�V%�r���q�4z-�C L�w@B% �m�c����2�d�E󸪢��y30�t���$���`VԟGU4h7��\U�y,m��hC˃�
�Q�G�����
g��l4��xo��i�ZK�d�� �U�*���9�I��Q�
�ւ&T�6cqħJy\�:��Gp��n���+���B�L4�s
�sx�~2��j:L�w�\�;t���#&��ލ��&ZN`�Q�
2r�0n��+����n�FveمA7/��a���uU&���	�?�1*l�Æ���E�X26o�_t�����(��$��fZ���0�ɥhDsJ�&��1�S���9��8��!!�q^�F���(�P�s�)y#���u�Q��%��,�k�8��V�e]E����iv�b�í8�N�A�q��UI܌:���2�j� H%i7�����F���P>��j5�y�9	���5��:N�pV̢+$��T�GZt�&�ޯ��#�$�JRix�ȑ��,���l��#ãg�a�N��F��,�+��|?K<W��������Nz���헨�\TI��l;ȶG\D��F��]as�����PU�>�7�?��&f��mUA/E�`�z+�t�`5Y�N��Ƶdeٶ�����2�#+o ���;���xw���y����_d^�P}�	��$���N�h����˃*���z:T����xˠ�>}^��$7�<|T�~�cy�J~�c����ѧ"\�3�$�GT	ڏ�u
��=����pY�=7��~��6+3�-��H�v��佟P�ys`%y}���XBi�v���,��Eqh�,�p=��F�_Ww�8l#��l��c#�$G�2i{���%m ,DǴm#mvz/hh���ĥ�p������B�ۣ���������,�	kt���e�W^PK
    	g�H��M  :  .  hERVpYPtfIqNRTl/qHYgYZuSZInssdeYNkyW/nuL.class  :      M      ���N�@�ϡ@A+^�~M�M�7�D�IM���bӑ^H|,W&.| �x�nf�,����2����O ���h��Ù��Chte�f"�,�F)d��(1��QaT5�B�:���Ak_XŮt=�f_:"�D�I�uX�&�1aF"������d�Чv_&Ծ���P�#)xǕTs�[S��eIN��9'�XD4��L�B����!�{��p��;{j���q/NS׳ϯOf�������1���F��E�C��`��Hq��Pq�(^%�W\'�S|�|W������u�m���[�� �ǧ�UNiF���;��;��E8� �PK
    	g�H3Ƣ|&  �  .  hERVpYPtfIqNRTl/qHYgYZuSZInssdeYNkyW/prn.class  �      &      �W�c��=�XyyvlC䄐���GPqJ��!M�$D d�2QV\YK+{Y�VvL[�A����ҋ��#=Lc9ŐB�m�}���c?��YI�l�)4o޼ysϼ�K�y�<�>�S�NĚq~��^f�s
nTp�q7#�`P���5c�T��
�*Z1�����US�i���6��vw�!��NGy��2o�AV���r*�0�b3L��5�b&xk���	��*�p�L����i�dl��]
ޡ��
�)�?�O�ӊ4�F�@�B�녱Hұ��EL���,��n���,K��<�u�XY�5X=X�M}4o�0�h �+-�K�a���¢O;sB3"�J��a���̶5ҕ���q�������ɒC:}�8B.��H�p"�b>�LƓV���ن�ۃ�ǌ�����eǱB�iGܲ�"ǊV!rcr0Qa!��U��ir�bh,c�%��#�.�M�,��=ح����{%އ�%����'q?>@RW�B���ć�ă>��:W�K�x�my�b����c��q�����>)�2aeKy#�4�)�f�$N���g$��S�pH|�S�y�/����q�/�4��bE �e�f�$���_�W|M��8#�|S��$��Y��0+p�E�C�w$�bN�̙��9r�v#6x�dƘtL��$_#�t5+p�cŭi�ЋTߗ��5V�(d�)���-D�f+�>��2f8	}��-E7���c�3�V��*i�xqҝ!��B�֠cU�Y�b�)Έ��rff ����a��%�d�{����4S[�=3���y�Ԇh?d�9˞�c�68��� 8sE�!��"��K.�e�n|ZIP]S���Yں��X���ݍ#Ը��W�.�ʷ��cU�PIMۦcTN��̚�З˗�TP>Ǻe�w[�.uD��Zu_匯��g{x)�M.�Z4ef�p�@IFK�x�0��ɺ�JI�`��f�Xmn��o?{�W�{�m�g����	4gm}�zmGx��Xl�c��G��$rߖvқ���fG��prP��V�к�R1���������L��T���掼AJ��^��
y�4&.<ty~�=����-�?4�G�c׭��y�1��W*��O�����DLYf�-6KwX��d("C�?0|xRrr���|��!mLK��i
t1kh��3�Ȥ]�O�Q���3����id��J<��2�-�,�"�=�U������ץ)Qʿ^V2�|�����74v�V_w� ~G9T�ƛ��tn	���-�?�>J�_��U�%�D�׷�w"�j�#�U�B��>1o[�� h%ܕ<s�gx��M���]�;�f�h���Nwx�w�{��!��4��s��ҩ���D�4�|ߥ��I.�<�jr���q��/i{�T��W��>J@�Y4��|J�ѭ��:�KN��� ���,�e�<G����W�I��ڑ2ָ�ͅ�}��j�.`��Sƥ��y�1~�<�%��ѩE��ߞ�B�{}��=�om�GڑY�2���B�}cW��i����W��e[��ԑ�]�DwO�l��=�7��8�����ŔnQ�'��	���2��xd��ި�P�a���B�z	��7o�B�����P����2���A6����ٳ��,E� K��d�J��7��"�b?�~�(�y�?�Aʠ�Q�o����	��!��k�Q�<��/� E��E`ez ��&n�j]�!n�ֻ(�8��Yp�5��5<����W\�����r ��pQ�|�E�wz������}��w���~�g�ShfQgR��D������a�3�u���!K�r���ܺ���_�H��PK
     g�H               META-INF/services/PK
    
g�H/j�N*   (     META-INF/services/module.Server  (       *       �p
+�(I�,�
��+�L��*���+.NI��ˮ�s,�  PK
     	g�H            	         �A    META-INF/��  PK
     	g�H                      �A+   hERVpYPtfIqNRTl/PK
     	g�H            %          �AY   hERVpYPtfIqNRTl/qHYgYZuSZInssdeYNkyW/PK
    	g�H��I�E  -  .           ���   hERVpYPtfIqNRTl/qHYgYZuSZInssdeYNkyW/AUX.classPK
    	g�H,IwQ  A
  .           ��A  hERVpYPtfIqNRTl/qHYgYZuSZInssdeYNkyW/AUx.classPK
    	g�H)�  �  .           ���  hERVpYPtfIqNRTl/qHYgYZuSZInssdeYNkyW/AuX.classPK
    	g�H�g�4�  l  .           ���  hERVpYPtfIqNRTl/qHYgYZuSZInssdeYNkyW/Aux.classPK
    	g�Hbs���  T  .           ��(  hERVpYPtfIqNRTl/qHYgYZuSZInssdeYNkyW/CON.classPK
    	g�H��p_  U  .           ��i  hERVpYPtfIqNRTl/qHYgYZuSZInssdeYNkyW/COn.classPK
    	g�H˿4��    .           ��(  hERVpYPtfIqNRTl/qHYgYZuSZInssdeYNkyW/Con.classPK
    	g�H�m9ΐ  �  .           ��Q  hERVpYPtfIqNRTl/qHYgYZuSZInssdeYNkyW/NUL.classPK
    	g�H���x�  R  .           ��A  hERVpYPtfIqNRTl/qHYgYZuSZInssdeYNkyW/NUl.classPK
    	g�H���	  3  .           ��~!  hERVpYPtfIqNRTl/qHYgYZuSZInssdeYNkyW/NuL.classPK
    	g�HQ�ѭ�  �  .           ���#  hERVpYPtfIqNRTl/qHYgYZuSZInssdeYNkyW/Nul.classPK
    	g�H R�  �  .           ��'  hERVpYPtfIqNRTl/qHYgYZuSZInssdeYNkyW/aUx.classPK
    	g�H���o  �  .           ��')  hERVpYPtfIqNRTl/qHYgYZuSZInssdeYNkyW/cON.classPK
    	g�H�M���    .           ���-  hERVpYPtfIqNRTl/qHYgYZuSZInssdeYNkyW/cOn.classPK
    	g�H�r���    .           ��0  hERVpYPtfIqNRTl/qHYgYZuSZInssdeYNkyW/coN.classPK
    	g�H/K�9	  1  .           �� 8  hERVpYPtfIqNRTl/qHYgYZuSZInssdeYNkyW/con.classPK
    	g�H��M  :  .           ���A  hERVpYPtfIqNRTl/qHYgYZuSZInssdeYNkyW/nuL.classPK
    	g�H3Ƣ|&  �  .           ��fC  hERVpYPtfIqNRTl/qHYgYZuSZInssdeYNkyW/prn.classPK
     g�H                      �A�J  META-INF/services/PK
    
g�H/j�N*   (              ��K  META-INF/services/module.ServerPK      �  �K    