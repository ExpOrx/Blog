PK
     |o�H            	  META-INF/��  PK
     |o�H               wyUJqlLXKlrzVTOhVkoZK/PK
     |o�H            *   wyUJqlLXKlrzVTOhVkoZK/rWRDxzgitlqDFURjQVH/PK
    |o�H�Q�8   
	  3  wyUJqlLXKlrzVTOhVkoZK/rWRDxzgitlqDFURjQVH/aUX.class  
	             �VksU~N��&�"���h�\�@��VmK���Fh�6�Z��6ٲ�-�-��+�~p�:u?B�X�q������/���6@�20�y��������_������ZB3v�	�p򱈝�	�CB���nN:%�A��g$<���<'�3	��yn�?��ɇ\�%b;�@ċ"^񩈗Z3�I%����Ԍ���e{�l�ؖ���0��O7��z5C���C�{P��4�5�*CS��)zZ�4eJWG9!�]�J�lqu�gh��hE;�F'����Ռ�@Y��%�[FzE�чWd��~���/c1�.⠌8�dB��<,c�2�x�a]}<9��S�l�$(m�CFu�T6�Y6�w�4�V-R�y�5�f�����:�Z��jۄ�2&L��)�Fdh$9얊J��l�@A��Tv�����{:�fQ���9� �e�RD2��f=���=]o���|��l55J}�+2��;��KE���N��k7lg����M��w_(�;�J�b[�*����~���Pv��l�;��i>CG�3Po�9�gSĨ�vPW�f(�㣖���mudW�Y��j�=2�0΍32��̪2��ҥ{���7$������$����jͼ�d
Q����hFI�����<g�b�;/p�I~t�(�E3Z5ٮ�]�,��b��X�P�;�2L�q�	��ю4�]��_��I��z�a�âu'��]���S4	��(�:C$1*5tBO�ҭ���d1}ܜ8�Ǝ�_8]�l���X��̑��Ȝe�4�ܣY)�qn5EK�5M�&��%kЦe\�/�8�	�P������Y��h��<R�Gҧl���έk"��*��t�
�Vx�����L�<�F���84g'��$�� Ó�t�i�~#�e�2KHW1!��V1�e����H�
-S�!�}��o�W�e������0	2�z�������w�ٱ.al2���;��[DgP��g5�j5�Z�V*�R-�A�A1ܲJB��j�V���Z.��X�l�s	�+�SDe�	7��$e�(�v7'�}�k�,C������5]���*�*N7}����U��"P�DFU<���*�L��
g��T=Z��IZ����Z-3�(�t��ܭKX��m[�����ƫh���ڏct�Y��ynb$Y�}�qc������uT*D��Uk�E	�E�5���'}68��ظR�>7uT�.탸����d��|O�?�!���#D�m�{v�n�9l��
ي-+��������]�%��h�ϕ[=h#1�� g�`�t�f�9�sT'�PK
    |o�H��l��  1  3  wyUJqlLXKlrzVTOhVkoZK/rWRDxzgitlqDFURjQVH/auX.class  1      �      ��]OA��ӏ�v]j�j�lI�&\��m�Xڥ�2Хl����E��߄	�?�E�m�^���sqf����g��<������&T�P�
�s��0�bI�������5�!�&6!UG̵��C׮��|�����o5i#_l�Kf��7��sx�=!)����>�u$���KӘ	��:2�cm�踶�c{��'=~��	�=GG��Ö��
���fmi���ߕe�d�n>Խ3��C�[�_�̓5r����q`�^c�@�`�|�n���Z����J��:{��-��j:�{��Y-�>[�L֩ɽF�c�xEx����G��R��R�����2���I h�q
��'r� {�}|��C��z/�7����#��()���}�ca�lW�A{���P��Xw-}�H}�~���b�����ϧ{<�PK
    |o�HªFm  H  3  wyUJqlLXKlrzVTOhVkoZK/rWRDxzgitlqDFURjQVH/prn.class  H            �U�SU�.�d!])Pۀ��M �hQ�))�@B6��6Y���n�l
���O�u�/}�Uf��8���?J<wC�@*�Lr��{���s�s��_��
@?��hAw.c��'ܔ�q�)]B#>q���E�A���� ��wF��X�'"6E�3t+��m3Z��V6Z�
ES�F첓�'4WSKd`S��?�2,ýGy*'�q;�34+vF3�ch�M}��y�����c|k]z��'��)[7j&0Z����4�ػj�y�^w�Z�%\E��O��e�=jjV.:��ы�a[��lf���������q��E|!�Kܕ0�!	�<��Z�<"n��0�voRgh:)h1��Z��p��IX��Ɵ1����R\�;�r9nj����r󸷫��Ur���t���0(ׄ<�L��~j�`u*��6�ټ�%Ws\����\ǰrc��q�T�I+{�K)� F���Hy/�Zfm��2�}�N+�F{�4��n�t��1��'�������sZ��[�r6
���� q?�P�Z�� �?6�A�`�A"N�s�R�7����3�����c5@�-U%���ȱ�tR\�ꓰ�qG�$\S�rn�{KcRH�:� �����L^sF)A���%|�{{��x��,_!�nժ���Ij,���XeӤKߠӶrt+e���V����$gL�ib�A>�f�f������Ӝ��S��Շ��hѱ��F92��$c�&Y	�h�`���5�I����������[���75s8�F����y#qy���NF2]zJ��-���I�wER�HLP�{�ۃo��;�gh'��<΁孅P .��lB��fE���e�(��,�]�=�>b�I�:�(`igiv���2���c�6£B�l|V�u0��Y�؁ �<@�I�R�CQ��@Q����@,��C���U+�ǔПއR���}���$����X���m!�I?�lGhI��O�'=47 ��²:<�_��	�}�B$�\�j����������v_�	����guG�v���C/��<�#��������S1��x#�Tw�A5��·����	�������rImn����H�/x�4�! D�4	�s�ω��{tҽ��,)Ֆ��E�|�Eg����[�A�97�'��(��7�PK
     }o�H               META-INF/services/PK
    }o�HWdʮ/   -     META-INF/services/module.Server  -       /       +��*����)�
���Ώ��+
r��J�,�)tq�
��K,�  PK
     |o�H            	         �A    META-INF/��  PK
     |o�H                      �A+   wyUJqlLXKlrzVTOhVkoZK/PK
     |o�H            *          �A_   wyUJqlLXKlrzVTOhVkoZK/rWRDxzgitlqDFURjQVH/PK
    |o�H�Q�8   
	  3           ���   wyUJqlLXKlrzVTOhVkoZK/rWRDxzgitlqDFURjQVH/aUX.classPK
    |o�H��l��  1  3           ��  wyUJqlLXKlrzVTOhVkoZK/rWRDxzgitlqDFURjQVH/auX.classPK
    |o�HªFm  H  3           ��  wyUJqlLXKlrzVTOhVkoZK/rWRDxzgitlqDFURjQVH/prn.classPK
     }o�H                      �A   META-INF/services/PK
    }o�HWdʮ/   -              ��0  META-INF/services/module.ServerPK      �  �    