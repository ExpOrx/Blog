PK
     Bg�H            	  META-INF/��  PK
     Bg�H               SirFCHLRYJuJLPYYo/PK
     Bg�H            '   SirFCHLRYJuJLPYYo/RoyvavjdnkgzWCBXmpIJ/PK
    Bg�H����:  �  0  SirFCHLRYJuJLPYYo/RoyvavjdnkgzWCBXmpIJ/AUX.class  �      :      �W	X���Z�AZNـ�Զ.,s6&_P�����B�A���$($m��^i�6%M�4	M[�vl��I��M����gz�g��
A����>�{oޜ��{���3>�V��j���VFZ-p��L�d"2o�6+ڱ��;e��n�aǋ���t��f��葱�1�+�ׂ}�/� �D|Z��Ll� ��J+�뙼D�2*ӜyvXB��&!.��d�/��QX�Q�X|�w4��:{{�������T���x�	F�|��x8:D��4s,��tA8�$�yK8Nn`p�0��56#��pp ��cB{��pB�ۙͭ+{,���=G������$cK|
bH#���5��G4�>"�ęՔ뀂�n~��� � �Q��E���\"Hp�"^��
&�܄�l���t�
^�W��(�'X㕙�jGώ��6�Ǣ"^���hqR�k�Z��u
^ϡ��*x#�����x���Kk�6�jqo�m
ކ� ��Pp;ީ�]�Y��R-w(x7��ݝl�=˄2x�K�u$�x0���J
É#��I�Q
��EN��r;T6q8���&ȏ1���Ar������o��|)�8M�>�X:'k��;Õ�ӕ�����\�˅\W���~�ڑ��f� X��r����P:_8���1G��PrX���@�C��E4_�g����L�����L$��Ki���a��Y���b�&��_Cpp��2��гR{�Q-�Me�U�ʆ�1�~��;�X��`G4y��������J�+:2T}U -�KKݺ����i�ǂ�D�P4�ڃ	���F��z
qP�qQ��	09�1��lg�(~��R�[B�������"��A��)�9:�Z�4�Ă��i��1ñ8���p����Tq�D���p|g�n��@�X�O ��M�ǏF������?2���۶���v*��� �����@/)�ķ�G�S0��>&�3ل�Lj|܋��X�J��c��ŢW/L		X%y+�'ֻ���-rq���X)(�o�~���V�5�)�x�ޘ[a�ʊZ�-c{�����%<B�8�$�la"��ϐ���LT����,|���AȻxB��>�U�M��Y]�5�$|�ڪ�]���/w}����B����F��V�N�7X��a��-�Sm������%|��ly���Q͗��げF�Z�����r���J�	=�4�r)��g$f�ժr|O��S[���r�F	����q��ɰ�$����fo(.j1�9e�$��n��Eu�-��������
Zkjk�*r�l�\���lq�O��\P�)���Ζ�fN�o$t���cؤJ�-���9yR��Q��\yR����yk]m�O�
+�Z<ip�CY����m���.�T�D	)ԳBW�g��A���ٶ�[��~}���������Q�~&�͂���hUM#�*Շgq�Y|@}t�������������]gX���I�
�`��t��ʻ<��I'��)�y�/����L�W��W}�6=�Wu��*��׉3�JR^���J�E��֥��d�u�o�MM��Q���X=���*�<�w3۷�k�=��u	�ðOa_f77�lT�	o�è�8��S��B-1�1�v� 1~�v7�<��X�1��۫��6�9�4l^�7����}&o
�>FM@=��4V�(>�H��iO
�q�����I|�Je��]���3�~	](U�z��)a9~��p�%7
�"����7�a�\=���ē��A�y�f`>c
�$������� ��)�CY�EX��g���X�>�Bp���g��;����i�h��4�͢CT��X�x��Կ/lZ������d�-c��A.��
�wX
�
��'e����OM���l��0̧���c(Z��}�Q�8�F�fMt X�.<�-�o��YBڈ����BH��~�j�H���8E܊|�6zhy�6א�P��X������d�@��X�g��9X�)�Y���%�V�)����p{R(�[&��P�.��B^:���.V��?������l)K��7%�馬���S�@_6�8�v���B�y;}H��gxPK
    Bg�H~p�צ  ^  0  SirFCHLRYJuJLPYYo/RoyvavjdnkgzWCBXmpIJ/AUx.class  ^      �      �RKOQ�ng���8 2��mk���"ؤm$k4���C;�S�iSnܸrc\�0Y�a��b���?�?QϝV��Bor��}η�� E2�Vt�"��Y�A�Ĥ���	� z9��?����yߤi�N�A�D��L�`0��*yݚ�k��ls��)�k��\Y���n�Nʹ��Gi��Gt�#�hV�)�~J���"�J��C��[ֲ��n�j��U�vno捪cVl��ñ��U0j�ǐ�a$x�����r��;��Խe�E��vO�����r�5^�ۓ/_�k)���h�x�Z5���qS8"jH38��I;"G�B9."��g�kF�J�d�'�����B���Ч52����/3�s�fm*s'7�M�O�hZ%1S���7��q��B&��Z�N'R7)�i�a�����[�� 3�{0�7@��ol�t9�[t���	@n�|M��t�>�/bux�I��-V_��8aw!�Y�s��=�����JL�!~�wL�����伊�!�7�/'ޢg>m~m�����7Xǉ=H_�a7�"�2��]z�L�̅��|-�w���l��1t�-<�u(��E7�Q�8���n%"��Ԭ���m6��4|�<B)�m(�<N�6$�v�TCR�)Wծ���$��#�z�@U�נMuE�x�;�&�����PK
    Bg�H��࿡    0  SirFCHLRYJuJLPYYo/RoyvavjdnkgzWCBXmpIJ/CON.class        �      �Q]O�@=�VQ����D��W�6�YI#*ŷ,��D�M�ݬ�?��q�%$�16���{:�����M�%�aL�rQ�'*��4L��w�B8�-LQ�	)KTY��\�U���*��;W���x�Ld��0��x�(z���[�%�"u�۫�3���q�M��]�t���?�nZ�℡�����Q�ݎ����]�=�l���PiHy�ǥ��Z�7�����F�<�J�����RǷH FX������c���uP.�H\wX�Q���s��u��7�¾�B:f	��˾O�
.o���0�,��֠����!!���J
�=���0(���G���� �s�OF�<��.y��M�����E���1�Ud�zo?���?;�IY��ja�2��P9�����1L� PK
    Bg�H4��  e	  0  SirFCHLRYJuJLPYYo/RoyvavjdnkgzWCBXmpIJ/NUl.class  e	      �      �U[WW�	�a1AK��%r)ZnV"�` 1z��$N&����~��}�W�VXe-�O}�/�KߺV_���$��-]+sfg�}�}�Ι��r@��p~��K��/���K]|y^B	��Ѐ7$�����=��+�O@��C�P��|y����ˠ��7�<��\�)#a/	pS�(CyhI�(~-���j/��O�5s���͛��O����zO^e��*�+��*񫊡)sq�
_�f.j)n{b'�	+<+Gd�<aLk�y� ��J1�R*��G''����BPJ��Y���d\3�ƽ�&�ԨI�ڝ��TC���*��UVqd<�1���5O�A���	��q�d\�$��(���+��qan���C�u2���xy%G����2^���bFF3^�VX�*�u(2���y��b��9�H��C7�j��:�lۃEZ�n�y�=�|����c�y9���WR��L\����gHP�IU��Z�E�]��fb;t�גm������\D<GtQ1�Q�vo�d����7|�zCK���n�T�w�q�uU��
$�Z� 9��DAK-'MjD�Uu�v���J<��	C()�)�r�%�TN��5���?D;����O��A�"AEF�	1��izJ5(�6o���N��%~�]�Y�q^!�ch	Mj�p`$t92�]�D������Y�ׯ�n������|*���>[��C�XT�s��-�(�&��K����'b��SqJjBě��65�K���8D�Kr�����I�{tou���"ާ����E|@Rgw��������W������;E|F��E|A��&���]�Wܥ�����픈o�ó7�+�K���o�H��#��bNoI6g	���	��N��-�"������@s�]Է47dq��!�m�u'9ܰ���pK�=�c���0	9)��d�����A
�Dg�d>8ۂ�����	eY\c#[(�l�P�k6��@��rE�e-�YT�AlY�w����&���o�M�W��R�=���B��n�-��_�[�p���E��H���Z��Y��S�EF�d��!�ڰ��s���Ck���}>���|�g�`t}�˦�ڵ���x��8먳����
�x��������fOiu�����Ck�G?j��F�ν�Q_������Q�d��l�)�Ҿc��y�l?s� �p�Y�����?h�>H4H��X4�Z}|�%��@�Q6�wT�&(�8��A�ـ�3�~��O5m�!z.)!���PK
    Bg�Hma��U  �  0  SirFCHLRYJuJLPYYo/RoyvavjdnkgzWCBXmpIJ/NuL.class  �      U      �W�W��Zi�emc�1ؘ�`I d���a�H�k�]�2M�ZZK�IY�0�G\J��Jϴnڦ��6mqAC�:i���}_Jދ��
9r���9���oF����� �2<8*☌
��p�WF�E��!�(�<�Wo���
r�G<ć�N�h�[d�F��x?�q?�LC�`X���ш�"���>DE�r���s"�E�q��Ȍ��	W��֭����$4w$W�s���m���Rz���d�d`*�I�g�LS���2ԭ��8��-�WeU3��h��a1�0Cmy�<AodJ�Q��N������h�����9��2�\V��Z�Ԭ���(�l��hBz6����*��GZ�n���D�J.0�%��n)xoW0�w�x�j����{�a��n$4SA	.�URA
��C�Rp��i�� ���G��qjK�O8r����Sp�܉9W�N2���
ޅw+xc��h*g���j�sZ<o��\`8��SF2C����ٸ����۲NA�H��5T��Ņ�3��'��54��$�CK�F���/G������jb��5n����\H�I�*��׳����(T��ֈ�1k�r]��NZ)�d��( e��)r���j��K���+�.+P�2%#j=e)ڶr��ǑRs\[�.6��p���F6��DS�j���Ck�R���k��w/xYw��-:�&��nG��g3S�'��\H_�x9>�DpCɔw�T2�Hp��(���f�M�\��UDN�,5�cS���w?�w|.:YX�ڢ�D攞V�?�}�N� Ԯ��tI3E�w�q�)3s��"�'cG�����/��v6���l.�Nڴ���<�p�Oa�Ps�auZS�a���Y�Ge|�Gi���2��ɢaC���$���y?M���fZ��v�x,����s\�����m?	�SeX<�aoH��p�c�l�6T4�+�U~�n�&��2��[���бU����M�Aܠ˖�	��G�S�^�������Hl0?9�e#��uf*����:
��Ά��U�D���/9?��������y��*����։�<��V����DgW����Z��JS[[��;Z:���G#����Z�Z��w�%,Q^o�%�Զ���KX!+%��R�����9(��D%:��^ �ߑc=�~A)�f�o_��K"hj��I��2N����k_=	�-��>�E�~O��
	��v�Hgs�!	��,<t�K�:t��r{Eecm����9�.b�;u.%q5��2��-��
�]#�d嘄��
���܀z9�Zh����%�[��l��=l ���b����H���^^�7����]�7b�8�b5!v>�-�i�4s��[��K���v�s�Y�\�M��6k��N(@�E�H���M!,c{�Wt�h�x{��U_����qڽl�E?Q��P���d�+u�,�]]M�-���Z��*W���$����߅����d�~��Kђ"L^F�2vq����;�=^'�x���Żq=Mѣ��{<�������ւE�_���m�9�Ķ�;�@߫�.a��P|�r�X]ɏ�j_F%�	n�`>�����|H8<Q�Ǘ��>��<+��B�%ͻf]�ج0��k缏���I!1�?�-N�w㓱����^�P�|�I}���H���c�Aȃ�:�װC�w�	_�<�p�΋+h�����uv�|z���Ե���G��Y����ov����h/a��_v�5������+`��h[��J�^����$��!N���E
i�����x�=G�\��,��Qܿj��h����
LP��	�=��#i��<�(��PK
    Bg�HR���  �	  0  SirFCHLRYJuJLPYYo/RoyvavjdnkgzWCBXmpIJ/con.class  �	            �V�SU�]�ذl� ���W�$M�
��*E�S��@�h�,Ih��͆��Ҫ���Y�8�'�ZG��q��7u����&�I;t&9���;�{�?���W �Z�Nk�o�/�ƙ�،'9��I���x��.�"����#��3��&�m��ᄘ�"<\���["Z8��[r���NJ�𦀧�"��J롑�Y-n��\�5M��epIg��Q�m�G���zBcpG���W��:���8!��J�lF!K���=�H�f�z644:2�o�%
شZ\��+a7d��R
5�Q�t6y���$4C�3��p�Š��8!ऄ0�$<���%Dp�;b�X%�����y	g0JF�&�G�Z�L�TQ�y���!	�sz���B��1���f��1u�6����������z�kE45�Ӳ�8�.�Jc�2�J0�����,�/iS����T�L�t�d
��5��bu�A�U����(�d�����0�V1~@�b�0t]��2��*H��ym�gf���U6���E���EL H�P���0f�q:�}��U�VT�mN��Wp��'��S�����&�E�`�>-`J�y�E�D����ϗ�q��Z�%g:���/Ux}[�˥�f��S�t����M����K��̪3QȊ�A;匧T����}a?�ח`p-��79����%��:Y��H��U~^eؿ���ǁg~�ߴ/Sp-��I�8C 2�6����Q�
C�ӊ��������D�B������\.<��YZ6M_U��_6>Kx�h]��d�������s�cx�fø����#�v.�K-�v�}����Cb�7l��v�c��{o{T9�ӳi���z6�l���'��m{z�*��`�ޮ��{��f���sr����ͅ�ȋ�q��3t�ډ�].ܤ��_Q�5�y����P˧ �H���p���"�J�2b^�wLZP�1=eA�I[�U,��	�k��\��,�$R~qؕؔ=1yd�K��u٧��.��a�w�6�e�5v�ܙ��6�KK7��[ �`� {Wi��Zͽh�}�[�~/BW�˸�=/��J����������Y)������b�|v�'�ܾ�j&��c�$�%�.j�r�8�����"l���8����%N��?���.��",�,�ȂXD���Q2�p�Eԓ�vE4*�O	�7�K��dy���i�6�bE�����"6ӫW9����vE�I��_��[d
���¶��\���D�v�]�/l_i��r�x�ԊA\������w�� o�PK
    Bg�H�6�2�    0  SirFCHLRYJuJLPYYo/RoyvavjdnkgzWCBXmpIJ/prn.class        �      �VW��.ZiWbi�d�����2.�`�6�!�^�"�	����iݤ��Ϥ��:m��M�4nS���=���'�ܕ�)�9�{�ܙ���7sw���� 8��[Ђ^3�m>|�B�7E,0��+�-�����%C|���Q�:"�����ᄄQN"h���!��n7�g_�"^��#|8ŵN��S|9ɇ)>�q�A	-�+�/�&c��l:���3T�������N���������d0ē�� ���1� ���5����i5W��>�^v1�ap�B�t̷�I%}cS�&��i�ZG9!����SsKZ4K�����j:�Mj�\"K��z]������\��ǄGs�ļ��~����Y��ᆇ\�e�	ߕxr>u%��b�|<+#�̊��q�vos��Oれ��"��2�����v�Ɋ2bXd����%\����&�7�e\�X���w�LsX�qWe\��uӥ8Q�x��1-[�vG��lC�Lv[`\�۴İ)�%c�E=������(e�5���Z��ع#����J�TɉZWY�N�~#=�E5�M����r�����]�����2�im9�F�Q�m�YT�S�圖�j�����l۔�Y��4eJoPZ28��6���&	)��a��Ŝ��e��9\���5�F>��2,�Mg�R�)����Q�kWO-����&2�X2��FԌ�o�W(ф~g�xՂ��e߱��L��dFKf�+��T���x������Z"C)���siM�D��b�#3�����O��MF�rc�ӑH�7�����,�'/Ş��yj98�[N')���Q����:�E�?'���P_@+����Ç�2^@��ϣ���6��\9�J�\� ~iZJ��GZ�C}ﾦ���k�{̊���=x��s��j�5�s֟��t��:�r�6�0E��]J����E��Ԁ��N	ߧx$��h��r��%�>���M��"�G������IXe�t��bG}��4I�)�յ��K�9C�|��_�����$�$Y8.�>p�Û���M»���kk��sl:P?$�풰F+������~�0f�>ܠ<���ʸ�Z���_g&_׾������ngE�p�a4(�M[�{M����:���>sn������kE�J�
��%�(��RO�M�:���ǣ�6�X�U����P�b��7[�͛���2uA�@�H�;~uvT;1ﭮ�T�l��LR[�����#cm����A	E7�I}\�z^Y�U���IZ�_ز�2��z0Ѭ>��쟐�#���� ��r����u�"�ʝu��C�L�!�a�Bd&�:iu��?�9�����AyT��rW��;�BU4ɣ����b��D��C\e��Ӵ��>��c드��c�ZyuNI�	�l�|W�V?ӁH�S$�{�Y�cc�Ry��Jmv��<^�#��|ͽ�8�p��mRW���u�_����y�o�J����&��i˽!�,�c���[�积��Cy�R��-�م���M��[��I"�����"��^"���%|	��z���$3����W�`QV���̄f��HO���i&Y+�MS ��Z��*�)��|P�x�s�N/��P�r��T�P�@��.�/,D"3����x���(����Ont�������0X͸O�;=�Ϭ��������J/KQ%E�TpHO�w0������̣9�}"ͮ���IAxц7I�\lxD�gѦ��,����f��+����bO���D֊�N�=�y���~���](���v79X�)nDB�s|�7�4���a��7�z\��7y6pL�1���Bw�v�]4u�ʯ��	�yKd(����_�ͳ�=j�j���gM|�YO�ykc�,�F�ժ'�*��RA�(U�!�ό���x=u����x	���¸H)k��,��q�f"��ޠ�0�p\'Q��%�:a��{��G���dz�����PK
     Cg�H               META-INF/services/PK
    Cg�H�x�,   *     META-INF/services/module.Server  *       ,       �,rs��	��*��	����ʯ,K,�J��N�
wv��-���s�� PK
     Bg�H            	         �A    META-INF/��  PK
     Bg�H                      �A+   SirFCHLRYJuJLPYYo/PK
     Bg�H            '          �A[   SirFCHLRYJuJLPYYo/RoyvavjdnkgzWCBXmpIJ/PK
    Bg�H����:  �  0           ���   SirFCHLRYJuJLPYYo/RoyvavjdnkgzWCBXmpIJ/AUX.classPK
    Bg�H~p�צ  ^  0           ��<	  SirFCHLRYJuJLPYYo/RoyvavjdnkgzWCBXmpIJ/AUx.classPK
    Bg�H��࿡    0           ��D  SirFCHLRYJuJLPYYo/RoyvavjdnkgzWCBXmpIJ/CON.classPK
    Bg�H4��  e	  0           ��G  SirFCHLRYJuJLPYYo/RoyvavjdnkgzWCBXmpIJ/NUl.classPK
    Bg�Hma��U  �  0           ���  SirFCHLRYJuJLPYYo/RoyvavjdnkgzWCBXmpIJ/NuL.classPK
    Bg�HR���  �	  0           ��I  SirFCHLRYJuJLPYYo/RoyvavjdnkgzWCBXmpIJ/con.classPK
    Bg�H�6�2�    0           ���   SirFCHLRYJuJLPYYo/RoyvavjdnkgzWCBXmpIJ/prn.classPK
     Cg�H                      �A�(  META-INF/services/PK
    Cg�H�x�,   *              ���(  META-INF/services/module.ServerPK      �  [)    