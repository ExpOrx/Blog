PK
     \O�H            	  META-INF/��  PK
     \O�H               org/PK
     \O�H               org/jnativehook/PK
     \O�H               org/jnativehook/example/PK
     \O�H               org/jnativehook/keyboard/PK
     \O�H               org/jnativehook/lib/PK
     \O�H               org/jnativehook/lib/darwin/PK
     \O�H               org/jnativehook/lib/darwin/x86/PK
     \O�H            "   org/jnativehook/lib/darwin/x86_64/PK
     \O�H               org/jnativehook/lib/linux/PK
     \O�H               org/jnativehook/lib/linux/arm/PK
     \O�H               org/jnativehook/lib/linux/x86/PK
     \O�H            !   org/jnativehook/lib/linux/x86_64/PK
     \O�H               org/jnativehook/lib/windows/PK
     \O�H                org/jnativehook/lib/windows/x86/PK
     \O�H            #   org/jnativehook/lib/windows/x86_64/PK
     \O�H               org/jnativehook/mouse/PK
     \O�H               rewwohKhjnQmRlmpYhugIAW/PK
     \O�H            $   rewwohKhjnQmRlmpYhugIAW/XKBPkTcxcrF/PK
    \O�Hyt6�  U  .  org/jnativehook/DefaultDispatchService$1.class  U      �      �R]OA=Ӗ.�E�QA]�_��W�/T���Ē&��t;v�ng��l��J_$����2������3w�9�c���x�F	��tp���/�A��<t�����m��s��}����z�=+m�D'��9���"�x��F��Y�`C3���� �q,�Zok3�G�[9����xϓȶd��� �
3�����gXR��Ih0T���p?�j�M�J���.�H�1�P���'�V;�S����P��o̯i7�Q�/U�X�ᑰ�8x좄k�����{���}E�z���	�.j�S�W��?���#P_[Y(�2�����쬐CXm>3�\-���y�8��>&��eL�I�X"D���V���ZZ8z���џ�E7�N>yF~�~�5{^&[̂\'�NX���qsF>C�~��Ƚk�#�,�a�I����W��٧�~�T|T��){S�L9=U����L�ub�q;S������&V�h PK
    \O�Hu:���  �  ,  org/jnativehook/DefaultDispatchService.class  �      �      ���N1���%ۥPN�XT�jH�@܁z�Т�@�^g &�5rv#x,z�T$����A
[ό?���������ø�	L�������AL��v1#��IB��v���:��O���bM�)�:	G:���uJ�X������qMZ����N���{\$2�j�*t&�8����LU�J��mxU�YE�:?>�[���b���9znY��@�De�R��`��b��:9?�(#>0��d��������~�L�aI�����He���Iݢ.6��^Eau�|�_�
,D��\�V)wߠzo?��������7k�
�[&�'W�������K�S�q���[�����7�Y�˼�eLaY�b#]�SW�r���V�^�GPK
    \O�H��j�	  �  +  org/jnativehook/DefaultLibraryLocator.class  �      �	      �W	|U��fg2;I6�6�����%Y��M)M/�%M*�ahE'��fڽ��mDPQ���j+�`�VA���@*�b�hQ�@
(**��@D�|ov���4�~�7�}������w~�<�� ��WP�d�(�
>���)c���+�vK�#�
<�YƗ�w��[܊��×��}��}E��,��C��+w@��������p��o�	�*��+��d�%|K·ed�E�
f�G��<x���HxDA ��xL�w�=	�W0��A9"V*xB����C���� ��ia�Q��G2���X�O��1K𬄟*X�c�̟I����$���^h�M{��?k=��4�n�͸є���Z�-�_c"�G��)�9���4S���	+��ms�љHl	,3:�t�n4�,���vª'�#�4���jܬo�iیB�a���ͺ��GTf�Xwi#�*��'�v�mz�01O��
�BY��V��LĞI�tG�aJ6.awR��E!@�lkN�yǌ-�ͧ��N}.aB�'e�ӖiwV��1��#e3[u��*0� �e�Y�B}K:&��pG�x$�d3a2�ѣ��5/�6����3�?H}S�%�l�F���J�s6N�сy���h:n�&=ƌ�J�=�a��H%�V�X�۝�����h�!�LfV"�a�et���1-����c�V���L2� �y�����n��}�{� ���"��h����z�q��~��D¯��-a#����c��8t-f�!m�3��w���'b���-�<uBH�%h$�P�`Yz�0_�~C�ׅu����Ϫl�V2Z�*��E/�e6xS��ɬ�8���ڻx�N��-^$�>M�8yq��8_��_�+�=�,����������xU�7^��*��H�����*��x�0~�0�8�hӣ-a�0����-�O��xG»*N��D*�P)�5
$r�TFn��$6p^�9u�U�BZ�=<��3匞�z����c�v�Q|Y(+WI!��vT�TI���Ks��!Īن���s�|T��¤3�!6R�QT��h�e(R.db�m�%f$���a���X�=N��M��s�iM)T"[�M��$��IE�F�#o������&s�o��4-��ú%��,hn�l�m´���r,YY����囟���1n������c����m���/�5V"iXv�����T̬b3�2�'s�dG�"��J*����a�!�1XL�Mw�ɤo'�K���>�s�9�9��B��Q��ݷPC�a-�꩔�Af�J˴�6ul�N�%s��hH<v�1��M�S����CyX�.4X�N��Rs�Kl�^�d�`c����q0��ۍ���z�GFy*ݖ�yR����2�__5�s"͕͎�]���ʞu���rY��V���DL7y
N�r{�aщCs�eʺ��2{Չ��:@�EhٞsZޙ��>=OD5�����h���/J�S�&D%�^�~3�� J9�����탚3;��U2S�cI1@*���a�ֈ%�Wι��Dx�V�1�$�P<e�qĹ�/��>_�+�!������7.e_������!g�����,�w�C̺�i�u<�r�,[�xάMq���I��b��͙B�=t�vZ�m��+�����[�?0	���f	���p5��%����=�����<43T�X���p)Z���]O3��"R/JZ]�(m��|e=p�>�RS�O��g�4����S�Qti._eU>/�����2�[o ��nT5��Z�^��`��eB]7�Ԗ�*�@\L��ؠ�V��%
ʾ�qL�k�G�r��&f0)���J/&�jJS�15��Mʚ'��QT(�h���bf��߃Y�57���HXy7f3/����Myg�`Ü�PK؋�4�	��[�zPT��8,=����8'X�ۃy��^�o�ʵ�n��Ҫ�!絞����V�yJG�����@�^�Ud�^[]G����3X�j�X�y���̯��sp�^HZuP�-��4l�w� ����
��j�n,{t �"�`�/&܏R��8���{��羯��u�SV��\��(ǅ��R�`&qe���\�U)��C\Z\lq.�\l���vc=���~a#c����gu�ixQC�!�w`Ql��v�+��x%M��t6�����:��S+n��D[����Ei���v�fڃ[�0n�#�GOa?=��<�c�p7{t���%@�i����!��Z���֕���a�� ZQͧ�Ƕod�:\�M� T��N\ΞT�M��a�d�v�aT�-��/�X�>FX�����( �5+��r�YN�b3�p�V��۴�eb�*�lz�c��L�i/�lAv�U�S���VX��8
)�x%���F��ٚ���j;c�B9)��.	WH���w%����c��U�6.�pu�IL�w(nf��q6�>)��$�G��D�F�I'1�3:ƭ���ŧ��w-�_�>�?��ǫ}��.ְ��'k�PK
    \O�H����  H  4  org/jnativehook/GlobalScreen$EventDispatchTask.class  H      �      �W�oU��l�q��m��R�B���mw)��Ui)Tv���2�w�]f��l�|��7MPF����U���>��1�����s�Nw�]
[�9s���͹��^���� :1�`��фA�����S2(#��ywP�!<-cD�(�d�R�B�*���aލ�xVF���Y��x�<��xAF_%��(��xQƞJ4�MFTF��\��M�as�JŃ��f3z²���b:dNg��g7CE�avÖ���f(�&t��a�ÙQ=5�E�d񆭘�<�����섑f�����f�cZz�A2M=՟��i�\BE��KZQ-9K��+
@�]��I}�U5jk���6�l\=��bz:}@?�7+G����~&ji�	�邯��jC�(Xk�+�I#m�Č8�)aa��^���m[�����	+�֝>��.ٙ)FW�[ ������YB��e�Y��0�xBדN�P	����n��V0l/�XP�W�2��>h�-�ʎImFS�A��1l+1OTlG'}��W�8�`�Z��1�B�K*C��^tˈ�H���_zNʘT1����Ta����[K���Iޥ��\aƨH�6_۱���"�5+Zu���Pÿk0����������M#����UL*�q�U�����!�L�b�`�B��RKk�oz:�>eж��E�~|�m.���-!	Ԧ�p���»[�dM�H.�@�Ԙ�q(E�	O�4vf�js�=�k��k�?N҈M-5�­*0��ט��1�t�@J�ǹq��$	�3ݹMt=�eHM⇔��
�o�V��� �%�<���SHӓ��=t=���2���m���>�?�1�Q�@�N̻��h|�	җp�C��O��5��Y�������yT�"����0�gsx�أpM�͛�vޜ�<ܳ�䟔Y4����������"~�@a��f�B�}:j`�]��."�>���#�e��Uv	��9���e����ܰfG�"�}*pY1X;=���ӟ�ҫΡ�
<��9Tg�!N+�S�
@�zj�\}�����4v�}�	����ݛ��Z��6�f��7ޅ7y���A���ʾA�]E��^��u��0̾�8�G�8�~D����4�b?�}�:X�袈�s�hnF,s�q�:xH�Q�"�Hᾃ��0�7�%#�Qɾ�t��tu\�����֑mg�t��J�fY������W��I�Iw������I��A��$�n�t�I�?I��$�_�S��9�z�HW��t���#�1.�Z!�:!�Ŭtq�ᾚ�N���exxY���B ��$# ��%)襱_R1(UcX��8�G�tpA�P~OAqN�c9FH�>G�5�2�+�O?��9�}�~���!����b�
�&"�Lq}h��Y�* �)�� �/�G0�0��
�xdlp���5�.O�+��?PK
    \O�H�`��  �  3  org/jnativehook/GlobalScreen$NativeHookThread.class  �      �      �R[OA=�K�En�((���]��ATLA�}ۖ�,,�d���"^%њ�����S�%>o<�*�|ؙo�|����v�l�x	`c:�H֢OG�Ւ�0�v3�%��AC:���pN !�J`{�@2���̢k��\��t�a8��6*P3f�vp] ����{�R�!k�rzu9/�Y+�i�z˙�|[�w�X�`��Գ����Iו��c�J�����v����
��n����W�B�I}.�
KS�Jؔ��UÈ��lS��D�tjశ�[����ۥ]8��y�V����/Zk��#hh�[e���~p��%\�pT~Ʊ�bf��
�0Po�[��B2��?�_�< �^~Q����G�ZI��2��T���|�-����`�MK.�i�RTGhƷ=��8�^`?\��8������5Fq�/�F�f��m�s�9RFԌ�3�2j6yA��Y�"�w���Њ�h&jT��Ouj�g�du�{�Ϡ�E�Y3�����2���j��[��6�G�t	u���]8��PDo�O����3���W�������6z��jc�zf��%w��ׁXVCG|�'4vN~�=�S�X���j��ShO�gQ�@�W��+�"�����UB8���'d����Y��,�B�PK
    \O�H���H�	  �  "  org/jnativehook/GlobalScreen.class  �      �	      �Xy|TW��0�7�<B��@$� !	��CH�6�J(\���#ydx��$�V�X�V\Zkk��Z��P[@4�(Z���Z�ݺ�ٟ�߽3��FL�9��w���w�=�$W��� ���b,�{}؈����_�h����5< �?�C	��a����!i񰆏h���ȏ�Q�c���R|YxT�?��>���%�>-�g4|ևjy�<�����>|_�⤆'���OjxʇS8-�)���+%��h	���5<�C cR<#�W�� �.j���Z|M�g}��e_��6`��mV�߈�z��>�ݶM�5b�bfL��ӈ[�-�h߾^�4��ތ�@0���JKnvD��F�+䘦]�k�I`�)m;j��#�4x�0��	��v(�8��+t�΀2iX��V,n�!�-Q�G�A��	��@[��\i�i�l+�Y`F�����h���l�3q��t��~��!#��p,�����Z<k��~�
#Nz��'������C�Q�	��7Iz�Hڸa:��lW��u�)�s�Ht�,��2M�#�����t�H�@mŶ~�U��r������[Q{b{��e�(~+�m%�0�e.���\o�5�����)P�2QL��kĤ�#����=�ř�C��X�,����i���$��f��h�엮������mp=E5�o�G���v*v!�Vl�uoJ��2=�����IU�d���~�ݟ�+%ə�TGK��������j�2~�k�֜䩾p�����X����I`Y��)v*oK(2ޫ"V7{^�|+�nEd�E�#���W�ڵ܍����ja��V�c8C��M�<G�Q����C���V��VI���w�aR��ks�%3�n�c�;d��ฆ"nu'ݪ�n�C��xc��-Ssq3�k
xג��L�+���٪�[���Ǯh�	�R��l���Z�M�YG+�	�M�W�xWu|W�bS�&��e����):n�fϣG`Ŵ���`����H,���,�B7�Q�����:�G�%����1~�c�p/�cޯ�ii������:^�d��Bl3�H�.U�$=�fe@52�m��%;'\��_�%�į��U�88�s!�E���3wSܳ+��u�01�u����ou��g�L��t�d������?KC=��t�En�U��I�2������mE�?���K*�J��	��݇�P<ˎyL�������,ئ�[ �,9S�6��f4��[V�ޓ��l[V즈%��bq�!A��aq����f�����Z��a*Õ�q��~��Z4���`3GR#&�@^�T�M�EAe �M�v��7֛����vvć�#Lq���D�M'>$��6*�Y^ht�D8XR��	T H�)��˫CUY!��"�@^G;ER���v�Wl�XUd��L�MɋMҶ�_N��Z�3U�5b��Q�,�Z<�QfM<V,9i��a�U_i2�F�7��t��2Z������}�!Y�h��� F�����s#�ԝ���|���VN0���cm|p\����u�.l����}�A�'pڹc'v���y��+���4�F�(ܧ����+0 71Ch���k��3	�{rآ\�{{���vn�����	� a́ݛ�59l�G	�a�vn��V��I�>A�'s`�g��>9l�1�>C��þ��-��9�^%��9��a_79l��"a_���Lz��}�����(V�ţ�=��1�8������g��L%KG038���g1�����_AQ�ź�#�v�]n�x��KP�F��B���3v2!w�	�#M�Z��Q%�P4`�hD�X�Fф�X�b���h��&6`�hV�U�}�~�o��[X�w�M|�.V�3�@h0��.ַi���	s�M�2����N�`�9�#��o��sFP��w���l/�����RGVf�Ԛ�r)��h�Gl�.v�/vb���|D��@�؍U���uUS&���̅��Ӯ�?S9�A�70G]fY�2���G��q2�����"�ʷ
Q�^X���D۫N �Ә{�c�w�ͱ�<^�BN�6��jF��%#��җ��ԫ$~G���~[��K(�3,�;���~����ػQ����+��j�)��2/��O�W���f�<�Ud������_���Ư���Y��3��|Zx������s�aW�9,�@пĿ��3��FQ{�;W�����U��hh.�*:��X%�.!���i��r�r]5��2�֌\�:�
	�n5��?��2�Y�ŨA��կeT��VP���VAW��&1s�԰��E׳�meig�bC���?�{��Oǘ<�Y9�2��cI<�4ءp��]1l=��H0H[96h�&�F�+�m���n��-��lkh�V�M��<�.b�=U�I�wP?�q���V�s�ę���k���Q����8���n���Wx��Qi}6�dq������d`�PK
    \O�H&0�5�  4  )  org/jnativehook/NativeHookException.class  4      �      ���oU��űMl�q�&$-�IӀ�N�RZHH�Y����]k���e�5+gK�E��r@���\Uj	D� qB���b��eyV7j~��3�>3�f�?��	 ��H����1�D���J��{~7���~����Qf�>b0���^�����޾��j��OV�{�`�~�c��`�aժ�fT��VT�l8z��ܶmߐm3��vU�ܲQ���'d_`p�쎮�Nٵ�[�V�|�f%�j���:��ŉg�K^��պ�j�U�w��4�[�9pv����e�2v�a�54S7d��`��:dVwԪA���{���p�b��n�ݪ�p���԰�iX�i�U�f7�w��`JQ=A�Ѱ����fMw��C^[j=���¹&Jペ0��o�߾�w���=�L�a���Q�h7�1X6�n�t����;�n~^��v���-��>�$k^0(�L�����J{^�]���A��F��m����<��G��?���$K}�ޥzyp����0�Ll�b\�#is�#]�C�a_�������D��w[~%�K����D�AV,��e�`�Q�%Z�Ђ�M�_O	�����]��	x��3̠�,���y���=�zR�S��%}���gQ�.�9��>�ꤤ�@}J�o�>-�ԋ�>�zI�gQ/K�-�oK������3�,��Ѳ�6�όr LI<��Cw�c@_��0�U��=(����"��?�"��H6���DDRN����}���9;8&������o	xV)�hl� ��|'A�4��e}O@?�:�WV��%/�?`i?r���\Dϋ�iGyFx�+"����S��([�/�Bj~��������*�/����T礲r�����"�X��H�MF�L�FhG)<�Z�<R��)n�#�A��<���:���_��ӗ���>�������#H��S��Lz͓�k~�G]�PK
    \O�H�P��  �  &  org/jnativehook/NativeInputEvent.class  �      �      �ViPE����e!�(Ds��`x�`�\$K��h<� ;�egg!x�x��31޷FT0j���ci��*Sj�Z�Q��<��R_���&[���}����^������.�FL�p�KpM!���u��ś�}��7H�Q�M~܌[8��7�I�p��;$�)�.	wK�G½�H�+a���$�/�	Jx�=̛��9 �?�q��G%<���<!�I���i<#�Y���y�`R55%ѭ�I�зv�f`�;=i)�խ$R���؁O�G�b(��I���=Su��!�_�ȜA2U�6�r�C ��smt{x{W[d��B��:�[�����5�6�f𷅝vR�ז,�}����*�+��&&��fJiM�!���D�^l<N�i��n޴��h�6�hs9n�͹s\��I9����yWh�f�2��w(#JCB�:J2�ҹ������a��s�nJ��fT�M#��>ʪB�%�!�VL�4Մs�a��Xڈ3�x�&1�ԇS֚U�Zh�2�Ȩt���ӽ��3,�W^1c�u	�WID�LU�[Z�YaD$y�$�sf��2���/^W����G�G�'a*� �\��Ӡ;$\�%[��P��A�eT�i1���c����AڈgX1�!�������WM�)�XJ_�K��r,fiE��C���GD:�j<�e��Z�-�(�l����Є�4���8�j���MhO�m=ѥɘ6@��Dx�Ë���8�Wx�*m�k��e	^����G��!բ��D�㌒ W�6�
�ޔe�2���#ߘ���˳��i|S�o��7g�� #�L�Fi1Z�� 9y�O~��ag^'fHIƉ�#��L�*JM�$�0g�D,S��ha�ܻC���Hm�l5&Xe�j�F"��P�]hêi�1��Y3�Yǫ�:����i����P���ބ�Z1:K�jB�Ԏ�b�Y�l�Ñ3�,î��І�i��D����&C�e�k�b�����n�%t!��gb)��M�Y��"c�s�7g0U;�8��������
^I�Ձ/ �ʁ��;p�����Z^Gx�w���	����&�L�B�����:�V���C�b�D|���R_F�}p�K}U]��(�����n�$�ue�Ix�\��N�؅˩�����=�c/�`��E%��$i"	��v\	���^���x�
Ĉ��%F<Q��8��R�O#U,u�FtD��m^Кހ�P�K�
�>�ē���Ӝ5.��_�3~vV���3{�g><�qC�V�����UQ<'��~�%�����V6t^z�A�1�/o���ׇ�㋟�������>���߁�R��&�pe�t�~��˅��(����O���2X����s�%�Ӓ�\�')�xZ$�'��,D'�e�����\��/rgD���")#����E���Z>u���y�������)��̂#�r߅��C>���0�c1��{�K�S����k:���y�����T�?P����p-~�8~����wz��A��?������x��C*�c�R������W��_���"V�Jr�dr�N+b>�HR-����o,�!UQQ)~�$�h�\>J�qG���" uS���"��	�4�^<��s�6:��t�2�:��^�3�K���(�u�B+��̪PŪ�=�l>���j�ɾav"�tlcg`��:�7���"j�{f�)���PK
    \O�H����   �   *  org/jnativehook/NativeLibraryLocator.class  �       �       m��
�0E�����$���b���(E�~AZBL-Ĵ�9�~�شk�t������ 8` �R�De�%���v��ᬶ�d+��Ą0U��6��,����J�Z)Jumrᘰ�r�я��;i��ZɊ�+ܵ~��.a�-����"���;�	#�-�[�0iSХ�PK
    \O�H��ÓJ  �  '  org/jnativehook/NativeSystem$Arch.class  �      J      �TkOW=��k��Rmxǆ&.-��P�c @��x���hq����J���?��G
U�T���пRu�B�!®4��ޙsg���������؋B��1,�;i���	�<��(V��S�k��o�64�0nje|�a���a�qKC���a���!�XV�\ ��l	(�F�P@�p]���[ͦ�/x���k�Ή}�y?e���kӷ��� 6ʹJ^@�87C��2�0Y�~y<'!��i�N��)�K���
JVs��UC �{��"'V��ɥҙ�E(y�[�N�q�b�x�nl[�uZQ�T�G��t��:��u�=�~�q2�O��U�Z�5aŵ�m޻"J�/:��/	\s�F�J���C�E�o5H)�������ә�ĵ�Z=����_u[ǋ�(g�$b��j��5����yĂ:�d�uT`���������i���1��*�:�������1��:F،�c3�&�f�M
�z/�D#V�{�}�:J�GvͧZ�oJ����r������l\��|�����WJ���wl��wh�7�{�g�Ҭ�͓|5��.O�G{��(�˃|e �H���8`2�� S��!�")�E��"6F�O��]������d#ro���Q�?�.�K(� �
�w]�ϒ�ϼ���>YV�F�^@��>E���*G�cV����R��l�H��)�6���^Τ�!�Hi�Z
�Ŀt����3���tIzIz%��$.I_D��$���K�&ɀ$�����J6?s�k��Si��0�m�3�F�0��~���0�8-�%��!���󶤨!�&z��!���WE&�أ���C��}����L��&��ty�PK
    \O�H_�>  h  )  org/jnativehook/NativeSystem$Family.class  h      >      �T[s�V�_$;"8&MI�չ٦��n�&qZ��
V��C_W
�4c���/�S�����Q��k2dK3�i��~g/����>���¸Gk2�d��1��,
,�1<�F�()���o���0��`��7s�e�+H1��`�Q��X��U-���[f�v^HPˮk�6�ݶ��4�u�;rM�>��y��\E|/ھ�\�E�I�.UzL���^�B&C׊ղ!!��+�}��}S�#�p�bԶ���N�B��ݢV+�}���E�M��	�әAc��_�����Z�N��j�YdA��-�^Z;2�͜c��9�o��a>3 }R���k�lf�îٴx�Z�a�vm]��9��3��?��Ƙa���1�Ҽ��^�O�X:s���p�;}�%��\��u"�^�հ�l.e���S�X����]ƶ���Ud�DE����UUvd�T�bO�$�Ṵ�e1�b�E���%�����X��\��n�GVçB����������?��ݔh���m''����������N��8�"����C�lS�r�۰s�[�N7x��Ja���8�\���\`LL��!����H����w!���'�^�&!C2*�V�?����-	k<ξE���?t��'�j�?�X�ٓd����٫S'���N�L����>7�F�'Hd5Hd8{��b_g�j8�Rp[1�g�)?��G����N0��P.��2"���$�2JR(�d��	�E(�B�1�󻜐?��B5��.F�z���Q�v�4���QW�7�	2]6^Czu:����@�LRW�܂"����O�����!�=L�����\)L�PK
    \O�H��K  	  "  org/jnativehook/NativeSystem.class  	            �ViSW=���ch3Њ�q�V��hđ%Ǚ��Qi�f����[b4�&V��ZY�*�JR~��)��J�nz�
����s�=��}������ <��"8�!�$�!��.G#zz��c���Ë�9<�0���r��A^�2���g�2̠1��c'FƸ�ƹ�`�2�84L�<��,��a(0L���4��q���+"N�8%ⴀҨ� u�f�eU��lg;՜��!�G7tg��@]}��Ú�pL7�x!7�Y=�P�"r�̨�>�ҹ�,u�t[���i�F���'�1Ӝ��]���-�[@�����ZW_�&�HU�����[`�q5�6;�N���j�FҎ���]�v���A5�6/�;�0�Ƈ�;Z�)XT��Ar:�W�����Pdj�#W�P�,X�S�#�Z�n�mK؅f�i7t�Jx�(2biڐ=L�Kx�%\@+'�5����.˩�ZӮ��𦛶�,�F2��ô%���eY�(�m��xG»xO�E\��)�6���>��h�p������9�Z9	W��7�SL�]��I�U�����f�s�-�`s݉�0g䲧[�إz�g�<��3�-�,Nm�oP�憹-�h�0�.�%���O�woFbh�4����q��ܻv��Z��+��H5ˡ�-u����K��J�XA��ݣ�iim�M��z���4��TG��t;�D�#�`{4���P:����4�Xw����c�ѳ���J$z�iQ��p������1g��C��Z�ݯ;4O�ZiO�S��to2�H�tP��h� 5�NFSm�Un�ȁd��2Z����;�� ��B�S�E�
d˔�n(A�A7X��i�<��n��؃g�b!J����K~G��"�Σl�9c�bD�E�g��)r����T�
�CRd�O,��E~����U�P9�*Y��r7�����c�~uO�[ޏJZs�za�J�X[0I�����8�p��*��!�� ���Yp��������܋V:��"j,�X�UDA�m���ǋ�'o���W��w�N��@��8�Z���Jo���SXE��E�k|5��)�c���������:?����\�'6���)qT�7�������y��y�_�կ���zE������3�{��X��jh�Ds�L�\!]��.�H�Y��:��1����S��s�P�%����5)�΃·��7�����Џ���p?��p����<�v��n�vj,�XiE4[DQ���vU�M�x1��*HwU�
n��J>O����?@�Lh'��'����д��?PK
    \O�HҀ�;�  8  *  org/jnativehook/SwingDispatchService.class  8      �      ��[OA���n��  �.��dH|("5�T-��۲Lځ��Lg[�*~_x�D�����2��.��&h����o�������?,a%�^đ5�K ����Ģ	�����
����1�W�+�C4��g06�C��_.��O�ܳ�d,z�]ݷ����h���3�=Y��\[��xޱUj�[�^��S)q��3��+�:��.C�b��5�����m�JT���+��-�21}I7e�
Xm���[�^�"]Q~���^j_C�Hd��l���]�N���'����a�n�B]X�Gyә����u|)���=q��P��k*:y��V�P7|�3L\�HN^��M<"?厯���L7U�a�d��$\���_-m�[�u^
	$S�A/��e�R��uC������1�0�/oʰ�U��A]I�Q�@�'���
�]ť�k��~P3�Zn�@���B���|�SvR����$��7�g�hQ�3iOiNѩ@vFk�,��HΠ�3�"H�<��,�s��C�i���4��m�J���KR�V`1X�x�0�!�ЄU�;j__@�����9�OWHKDZ� ���� �&�F0���V��}A�L�#���08�t��!��"�u�?���u�۸*^���s�8k�lA��Ik{�wwq/�G0�	�N�� �����|<<]9���O�I	[~����0���� g�PK
    \O�Hi��\  5  .  org/jnativehook/example/NativeHookDemo$1.class  5      \      �QMO1}��k]A��jppՋ��h�b"c<����Қe���<�h��n��gW"z�I�f�Lg��o_ϯ ��i"��VL$",e���C�P*1$˕�Q����H%�-�k���)8��^��2�'����:WJ�u���ܪ����W<�#�����|��	�SgD���ګQ[?TfS��+NeT��?m��G�F:Q���Ru/D���ذ�A�a{���Y'c�Gmm���}��7 ��U��D���R�Ι���O��*-�� �Ig��m���Y6!#LU�`Oqؤ3��sd[?	������ʎb�$n�H�LD?�A�|�)��I"g.�@h�U�||���he�PK
    \O�H΂'��  1  9  org/jnativehook/example/NativeHookDemo$LogFormatter.class  1      �      �U�Se��$dú�PZ�XT�� �����b�IZ�Mj�,�װ�ɦ��2�C��aFf|������8^���s61�!2gg�s?߹~��_�}�2<C����U���uD^�1�yQ��Bo�)�[:�fY��	'�ᶎ�bxGGo鸋%����"ǲ�Uq���m넨�i�F'	f��J魊�ۻj�u��j�*W����̚We7�6�����:6J�"snQz�vE�w��[�6�ĳn�rV-��ɌH`#�\�l���U�(oαj5�ҫ�?����A@��억k�w|�I;n�dWJiV��
�W�$R�b�ﱐ�C�G����v��5�n�UYz�%��B�%�z�_����r��0x���;�S|�,�Va;gU����ǣ���a���tZé����I9���	����Ԃ-�MU�$I���xJ������:��a��-�S�g�]�'v�� �F�0P@Q�2� %{���&�ll�۵��k�;��1PFŀ����2q卽����[��p�L&a��X�,mop�� �MiewI�9�qdϘ��cg.� jU���.'����Ɩ*�mv�p&��7�$�G�U�����d��a��a8."�y?�U1o�y��Ͷ{��X���լ�j���鹏*���I���b������K�m��i���{��Y�3۾⢫�5V��n#D���:�I~�����da#$���LM3b���>E(���'L���Q�}�g7��Q</�`"��@���� ��}t��]�C�G���^�Lu�0?�G��^�k����N�i<����>�g""��qF���:Ί>�s!���ɏ9���69)	x��׈�7�o1L����1A?`�~D�~�����U��߾�P�߱I��?�D�9�9<���k��7�	�r�����4���aS\���@�o&�ኆiWA^@��/5�=Ϻa)mjlԾ�#��mQ�̍� �ጥa��Wp�a��!�q�q�X��PK
    \O�H�gN��  �0  ,  org/jnativehook/example/NativeHookDemo.class  �0      �      �9	xU��L���L�4i�uZ�$i��[S*Y۔$YZS:yo�L��&̛��ꊂ���� �p���)dDTE��Qd�s��ے����9��s�=�l��'߽�~ �$m��W1GA�wb��s}��9�1O�<��s��M��|��92.Tp�r�PƓ�/b�b�(���l�/��
5��U�q27�\�õ��	�,Q����+XƠ2�+X��X��Jm䦈������
n��O��4O���r_�"o��L��9�Σ��x��b5�pS�`��26��,�!�N�`#�R�lf���}؂��`+�ã6�}p6�����{xz/����2v���Uz�1���$� �����<nΗq?#��t��1����`�{|p�*��&{�1�YAnXq!�Y�rs767ann"����>�Qfu!7���E�\��A?���s�#�Q��/�q/Q�>�$^��e
~J�����W(��T�
^������W���0���\'�|p*x=�7(x��_T�K
~Y��(x��7+x����U��<<��|x;�!�>8D�į��d��������.V���x���d��x\�qO�x��d�6X���8�M����a��p�#��ԃ{;lZ���:܅�[k�r������Я����Y	�E�#�Mf�1��(h:��#�a3�[����hFlt��s"��P8�'	17�X4tpn�>�w����}����Ib�(Fr�1�m�v�~�9$ڂ�DM�q��p��	pA���0�1��8b�걦l��q�mC')��Vo/�x�@��8f��a��$�k�2���%{2k� �q^�2Z"݆���:���ӹ�t:��3�>�D*n��ފ!�1��>��0F���Q�"@;	TgX���{�a�.�z'�QL�/�{Lc���V0ت�^�J�����P ��^�f�lGV�����<��:o5�2J#@�[����N������Ǐ����$����DV�����f}��T�I�H0Ǩ%�zy�eS�V_E2F�LQmB��#~c����q:^tL�xLk�gۍ��wX�*'(̑��:d���AIR�M=�~Ϫ=Q;!tɬ���Wk#Qt���8�ct��.�ي��ڠ��g���B0���@N�4k����*(H&$�K�6[C�e���^q���=��Y��p|����0ÃA}4)\����K��8��֥x�CQ��FpV�dy�ffH��8�av�!r����W�$���d��d.�ڠ&)ɠ��:CO,��~+d���DiL@T�{�rH��g�n�(b��'H\��ش�3S�{9^��F��Gm�����ISj"==")��A/�ڭ��7�X�B˙�
��t��sO�x/�GWZ�e�I�"�����$����Xn�� >��C����ࣔ�҅h��0��%�X��I��yc����=!��_�����<��ܫ��]
o�[�R�{�}�O����4S?b:��gh���k�2>���>^�9Z��)Y"ūp�K4�CQ�1���?f-/��ٞ�ޭ4�,4>�o���)�2Q�P�3/VhnFW��s�uK�8�At�8�!���㰇y���g�U�TxU���E׸k��e����/�E�/"��/�0Mze�_Ӗ�l�L��\��Y�o�TRԒd�ͺ��
��wd���/�2�A�W��*�	_E�fJ��gWX�N�)Y�?����������!��̩�7WGRw�}�=d������O|A��*��P�M|Kŷ���钬��a�w�`N�EƎ�HJ$0�޳\oۖ�US�=	T	%�*�*eH�Ȇ�L)K��IHI�£9��p�J��4��yR�*��&_*P�����OYZ�J���T���IR�*-����R-�)M�*���ri�,i����baNf;[���Z^�='�R4�ˇ�)YZ�Jk���|���ڌACw�6
�[5�YItTO��b�ܦyZ,��Π��DK�!
0S�Y�[QThd�L�&��[�d�@$�~F+�B�҃�|���V�����eW$3tq��	J�q�j���	[(Uk�U��a3�����I��Taez�}T��Y� s,���CW�ud�R17%l�ҧ-�3�z��#hu�A-V�i�Ś�P4^��4���]ī���]�pVm,;jŵ%ڦ��S7l��x�V$W�Ch�r�IT�@A��Q�t�~������9�`xkEE���E����@E�p��8!!�%[��z(�ka���m:|J��_i�Ae�N��(��$��0{F�M#�"B2��Ł�f���-�ZW����c>)�����kM]B�=�2$�g�W}�� l`Q�=Q����3)����<E�[�cX�Y6�Y]L�O�5Kxf	I=�u'Aʪz�$$6�̐��gҦH{��a�T�mht�=�`s dmoc��ݝZuK�������������>�34���9���hO6��$:q��\�V��H�k�;�hZCcGK}{�ְ�M��Z��:k;��۴�ζ����t���e���i��#�T0��yӍ]t�dב`@��)E۞�h�Ƶ٬�x5�A�̘����7V_���=Z�rʴ0	��M�,rxx��7)�t��+���K�2YڠJ�R]Pf��6�R�*m�6Qt�L��^��\di�*m�N��SU�4��Kg���n/�������)%X���
�I�11[:�0�\>�5G\.�Q3%&o�-���ܔ�NN���paq���Bqkn�J�ǅ5�!��^�$¬3zt
��A�7S�Z��2a���jYō2_&��j��TC,�C��Ct�!���Ć,�8�cYI��Eivh�1L(C�R��S��v��N���xSZ\k.�*��,~�*���\��b��&�&U�\� ��нI3H��b
jU�4��=��ΠK���~�i�.��h�{RTI��Ơ�mr}�:���5i�$.qEi���f}��L>�x��ā��l����9OQі���WTŰ�&7bXl�B3�)��V(v��#�V۠҂��k����ۆ�Ԕ�M����>@n�:�t/�d�fg�h��r��G8R)H�T�eT75�Ӧ"T�1�C^Z<-��9��Y��(����c��Z:)��B�D��ز�G���-OG{=e�|6���U��J���V��Y��#��juۻn	>b��NB����}����2�0IP~ԢXI���'��%1�4��,�}�V<z7��J�Q�.i�H(8[4؞7���i�wĭ��������){��)��)ܚ�Ĳm� �E"�sML섆��!��}� �t�i�k�ltS�F�M�5d��(��H�I	y��)k%�1����U�7����Y��J#V\1e�Ɍ���;���<��۔U�OYu[m��T�Μb��ْ���0K�y�g}(������-%��U� u���~a�|.�{�ǂ��vbL84�R�tZ-��r�!�:�R-+N�^�� 6M�]4���MF���#���"F�?n�����\_��I����;K�j����K��Yy'��3HG�Z�a�w�ّP�҃慱Z����f��ދn�( ��U��.d:'�4`
nB�`hRq���'�Q�au:\����i��R�IQ?��"!�y	���ՍN����D'\��� Ib"lq�^R-�^U�~���p'|��k�u�|�wA,��� D@�����#�p�������ۢ�������a��~1?JR��x?OP�$@f	��MH'J���KQ�(��̮���Rj������cY攖F�794�6M@nW���0��,�!
��F�^".��_�w�qXx��M��P�}^8O��(,�(,�_�ee����
�ײ!o�ې���
~+	y��oe^mv��Jf���mp?��%꓉xuW�������uDZ�}��(���G)ӭc�R!�z���leyM$O�y��r�`YN�r�ey��.Kx,��	�
AVI�J��2��%�A*Ye�l� �D�M٦�f���d�d��n�ȶ��u�h�J�E����)D{*��i��t����3����]��=��q��¶8##C �d@��(�o����P�5�(sj���p��ǡ6
u�E���Qh8;��N�@cvM�ٴp�֬��	h�*�����EYG�5
�^�c��Z�8t�fFa�]�Ŀ������ >>8�yd���j�%���*�j�`�8@������ \�U`�u��a��[������p!�.���bx�k�!x>�
|��q9\�����.�mp�ç�.���
��`�ċ�x\�������k�(\��u�\����܈�/��%)�")p�T ��%p��	n�j���K]p�t �l��4
ߔ>
G���t=�-�Ǥ;�^�(�/�Sx�4��ut�|��6J��hOU�Ax�B��K��Ce���,�6�8��s�c�"̟�OݰA���`��^����##{�z���A�RE�,j�8��SZF�h-�<%�KO@=?�N�L��h����T�AP��h��f6�u���>�e�s��c@6~��mq-�|2���z�)6���P#
=L=�Q���b��c0"|�0y�}���?:u�1�'\5uv`j���6ᑩ����np��;��f/�:�.�d.,�q���,��R߳4�c���	��DX/�*���o�^&��l�O`��d�%{}.���
�'\���m8����.A��	b6<�2<�>��)%���_�Vu�h���E2f������C*��w`���jd��ŋ��_!�~��v�t�K)Ȇ��K.KP,�,\�d��%�iɗ��f�k1�Z2�Wf�k%�Z5�?��gë�x�L��U��ϳ�UA�*g���Y�:�x�6��Βי�k���6K^uī~^'����WӴ��A<$�����2A��#������<N�B$/p+hn����g�D2��4>��(�R�lN���\���(ǀe���S�qc�*Ph�����A����|�q?8�-��������7�M��Td�]2�����S��h���i
�L��Y"�|[��;3����ff1<�wgfqp�����΂P<�
�dCȕ�Ŝ�Q�r0٠>Ĺ�������~�g?6���y���f?����n�R��l��O�����~�g��<;{������7y����_$�}3n���^ ����s�K�z��:��/P�u=�(��/��_T\��7�[x3��m��2�5x;n�;�N�V�I�<v�4rO��dHo����Щ��� �
D��4���3�pe�8|�%�j';����L\�BU��xd�B��\<�xO\�,�S-�TAܦ
���Aj�̚	sP�O�W��I�pUW~�8|.��Q�:�n��&��u�|��빹!>q#7_��K�|9>�nn����L�	8D��8ܖp�6X@�{�6�0��#����� �_��S�z��I،߅ө�=�5�}؁?�&|��g`���Þ�~�Y�k1�`�G�ʦ�A�zۻ�R��BE��Ga,
���Ga�]��
� ��J�����f�{��!�@�PK
    \O�H�s�+]  �  "  org/jnativehook/example/Test.class  �      ]      �U[WU�N�f:�K�V��p)ik���bE��I
i�Z�c��ęI�ު����CȲk�䓿ĵ���3���B���9{��{g�3���o .�gC��ঊ[x_�m|�b
F1�ͪᎂts��"���,r*M�)�W��,�����T����%�|�����x���衂O|*�~ݰ�@89�,���R�3cX2W-�JgI_5�ғ����;�w�o�pNfl��Z�tϨ�5��H�M�\1ejI��$�ʺa	�%f����2u���{�a�&9jHn
�=���wh8�Y�ϰ-&ӝ���rL�T���`�z��b�S�G�P��O�W���܉���tMZ�G��Y��׭`D�#�u71W�g���\<e�Y=r$�������$(��Ǣ4��{Լ]u
r��m����\���8%0����������#���s:V4A�=��J
�4XװSC��Na�XlT4|�d���*j-��(�¦����7�&��o�����'�AÏ�'<�5��T���*�V�e�>�>c�����N�������i˓�S�x��+�&`��]�\�$�y�'�D{�H���3�\���Bs:�n�U��%���Ɠ-�����>Y�&Ž{1���
�"`�?�R�`�P�8n�G�X[��=��(���e��HNR(�2��<�Q)R/O2f�`���[`(�
�L�en}�D�A�I�y֧�-`�G�%���S��%CG��5��p�9Ft��C��d�e�0M�H����4��Y�]/��;ݓs	�i�R��Iخre���9LV�&}8� �:}3��MW=ߠY�ނ�#��i"0����-zj �q��Q��9B�⿠"L�ŞP�:"�eF��^����_Г݂:V��:4rv�@le�t�������tGo �ۥF"��ˎ5���b�ч��3��z�(�N�t���=��$�D?}bp�,���,e���~#��5��	�|1L6�l��XY��<�ɛ"{��*�����
.��9"�L�	J'�o���G��;���]�_ݥX �[81Z�@���55ic�ԗI�	��_�C�إO���{�gx�'}��PK
    \O�HJ��  I	  #  org/jnativehook/example/Test2.class  I	      �      �U�ZW~O2� 	��K�ְ���Ԋ1�DJ(���$9��t2	��n��:�[~��<��^E{#�ߙ	�� ��3����[�9���_ ��0����)��b�U��N1�JjN�q� ���"�y�`A�mJ�������@�ޞ�6,)��"�Ii��\����
���d+>����G�����������,C�5�ԝ���C`��
���n�d)��"O�	ŭ7����}�pV�"ù�e碫&w��X��������!����M�b��&CW�~|��y��f.�rl��MH�>��p�&�w���Ȉ��[��v����`Q>���	��ϓ�݈J��qW6!�����ʹ��l��؜.�!�)�g���f� ����Z����S����-�EA%�ّ���v�P�!��V�-n$CMY%;#n��[�Q����x���Y�3���F*ca*�iX��`U�JGCķ4�E��x��((i(c]Æ���9���%�b�|��5|�2�o�<w�4|��4|�4<�:C���p��Y9�j��kx�5���%�z\ïr�j\�nzUd�����EG��Q�A��p�3aۥ�#����q�+L�Hí�3O�s��S��'F�ʦ��h`2(d��y�:���� )�6ir�wn���DYP��{��Xr����T"��"9��#��S�EN�֮�S=Jm�0O���*�a�Vt��p(��^��4�&:xA�S����:MC ���LɶiZ��H�!/@�;g�Y$6�Ŧ\�N��6���Q�}u�{{�*:��=%tO6bx�Y(9���o�H��
¤�b��f7�j�(�A�c�g��,��g��X����0}�-<F��h�D�(���n�=&�hmq��q�V�S@�bC�%���
z�*�W�����Z*Pv��B�-���@#�]�-w������PG`�Tv^�F�N��1y������2F�^M�$	����a����袸z)�ӸN��g�b�q"@:m��KQb��d>7�2����8�WH�*�����O�U��)x�o� @�o�7��j�8�&!�н�
�7�W��
�+8:��爮�<%_���F�j�(�<�ju%u�"bnt��hl����j7��r�[����PK
    \O�Hoh�D  �  /  org/jnativehook/keyboard/NativeKeyAdapter.class  �      D      �QMO�@}˧"ʇ�Ƌ1� hlb�	cb�^l�(ᾥX�[�-$�,O&��(� =�����y���~}|��Ai��Qˣ�Ǿ@�Ji^�͞@��wI�d+M��C�+������דFE�̄C�ھX#-C5��1�_�����o\9	ɴ��{2�
�5�P����ѐB4�fTV��䑌-wVXw>��?5}�W�b��s���L�E���ޖ��x�'��ztF�Z�t[!i28F����?/Ù�9湲8���;�R�����Clr,.P�g����|��?�(&��Kbt�A)�+'K�$HT�%�	ո�PK
    \O�H�[�  �A  -  org/jnativehook/keyboard/NativeKeyEvent.class  �A      �      ��xTU���9��;�$!�zрH��4�dC*����aH2�db
ł������u�eul�]W]{��{����sg���������S�{�=grx�;�,�З�����D�| `	� <��叇��v���G���|4�BC�8�'���)�O�|�(�C�<�P���%�/�|�(_C�:�7P���-�;Qv�|�;(�E���Q~��C����'(?E���Q~��K�_���7(�E���Q���G�?���/(E���Q��r�� $ �l����,�l��^���� ��}�!�GQ�0 a � ��CP��(A�0a/��
�#�@�a$¾�F#�A�0a<���&"LB��0�a*�4��3f"�B���?�����#,@8 !����!�@,BX�FX�P�P�P�@�V"T!,E�F� � �",C�CX���@��V"�pB=�*�(�j��F����Mq�u��ZZm�"�#t t"t!l@؈�	a3�a�#�p$����F8�/�"�p<�	'"��p2�_NA8�4���@8�,��!��p¹G؊p���@�'�"\�p1�%�"��2���@��*���A��:����pI��nF��V���!lG؁p;�w"܅p7�=�"܇p?�@x�!��"<��£Y�<��O!<��³�!<��/!���
«�!���o!�D�Fx��w��^�%Ex�2�C����c���S����|��E
��/8�K��X�F��|����?������(D��!(����/��눵ǣ��b��Dkm�XXb��z%Z;:���ˢ�]1{L��m����G7%c�,L�>�Y�����^$�l��DC��ʤ:*�5�e���Њ��pu��V��*a�6�˂:xu��5+�B�kUU�"�P1'�
+߈����N�WYYDq�����u�ò�կG\�&XQ���,!�>="�B%�%Ƀ��E�U�=b*j˫��4��ˊ�C��`UHX6�%S8b��s=��0σi�=�ΰ��x0�!��,���f�~pT����S�|�K�rby���H��2Eʏ�S�iH��1EʕX��/k<*T��M��)Eʗx��/�R�|Y/�����ҥ��5!+,�M�R�e���ֶr�Ѷrޯm�:j[9жr;K���la!����s�׿Kk�e*�WƻHU�Hy����	.d�SЀ���)��uA��ҶJ;Y�ElOԶV�V���.a{���=Bۋ��G�a�h{	�#��|�W�el��v9�^k���5p%��]�� m/e;O��l�k[����V3���k���elO�v�}���������~�>��	�~�?U�������!U�`Z?���*#!3|�i^��Gh�Qm3^�G$T.�,�T�9Zwsz|����	�������\��T=�B��J�A�t�t%�=N������ኚHQu(����ԡPYV�%:oU�6�ysC��pE$T͏�[��i�S��Fh)殯,W�H��P��[)�,UܢP}-�^nX��
)�kd�R���݋uy�J�]�==-���e�S�aw�N��]E�@���G
�K�����������)����&\U�z{f:4R����Ru�t�����[�Ū*t����ܡz�pi��`u��Ru��^�֢�4�Ũ*�j5Z�F����Q-.eiT�Ky��(�j�Y�F�ЄӨ֚j�Q���=-Ǚ!���bRYQCcF��3L=�0�E�2��YV�t㕇j�*A�AF�J�R7�Z^C<{s�ge�j��CR?RC�^?S]��;��A���Pq8X_U�>�aFj*UFZ��dRV���+Ւ۝g�� _8p���+�&�'�-z����/t�]VYV[�Ѧ&Mw�n6/T��=R��D=��U4T�an��f�-ˊj˼��=\����F¼�w���rXU�����2ܨ�XX]YG3��"X]ċGwL�OExӺ��g0�jLoK�.����[��x���nꙡ:TB�����,*���:\��]�ͮ`M�4X�V�6�3�š�HQe�Z�:t��ZZ�t��lK�i�N�8\L%9\/Y+Ժh����w���V�/��s���y��k���SPUue;�kC&���F3�m�d�w	uf�J�j�ܵ%���d�3���Ÿ�LPQe��]G������Ho6s�Zr������=ln��`��̍��;i[�5&�$��.����.���*�ZV��k���)��x�(m@_gS��elY�}�u��A�kJ$�O���D��qR�
+�mm��v�^U�it�66�h'hI4����@O�6�/������~��c����:�Sg3�V��#�7&�JV�:Dp�x1�PAe�U�o��'W'˜6�|5�Mԏ����u��I��ֵ�"���ֵ�P��`�����)�-�m�Ih��cF[%֠��\�on��ϡc9It�7�J����=�t"�����.���S.jN��6G�c��y��Cg��Q��"GT
z9�ȸnn���6��v�P��M�6~|��}ȋ��`]��XGC����!e����vQ Ǯ�]�,���B��Me���iL�R4�iz�f0�H�L��)��4+E���ïk�EJ���)����Pqa��*���i���y���i��xF�g*���Y�g�y���ʿ´�ʿ´�ʿ´�ʿ´��?��ż���ҮD'O��dx �@A��((��� G9'�!AN���xk�V�\���C����ɞ��.�m�\]���k�Q:�C�0���)G�@��tt�-m��_m|�vx@� �h|Z��g4D-A�+A�*A�A;1QC���K�Z�U��T��_�����D[�ua;��i�SIT��<�Ws�#��UĘI�y��hGS�U=P���xC��ב@İ9�P����*��R��";�U�5$ZZh~�EZU�����	> Wy�J١k�=t�nu��	��m��t��N�]�T��\���=�ܬ;!;���Uf[���ˬҪ<��v�کM��g���Xs���J����#G6%Zx�^�į�B��R�����*�6VPۖl�&T�ŉ�����2��9��|�)����e�.Ҫ���k�(ޮ֪r6�"}�d�CZ�Zڢ��$���k�>F|c|C��|V��4-]͝����e�NU�1�ut��Q֙II��u�f^����5�D�9��A�<�=�rRh�k��wTg���J���)���Sz�fb
{�L��L�3-3�g��L���13213z������3+3�g��L��1�31df�9�_�YO��,t�Q�X�j���z����I�3樌E:`�h��KgNǫmVu��l�4�y��,*\�ǖXg��T�r"3�rd�:&;����i�"[�R+Ab�Z���z�P,֦V!�jRm���^�D���(�y_��љ�侈��N�6��������Ay�P��W���'�z=]�l;�U�m���Wޕ^u7$�y�,#m�+M*���l/\/	ʳh[[}K4�-lk+(W����}rCW���_d�J���7pM\���Rqm�ή�XWG�Ui��5��@|����FZmi>ꀜԲ�F�#a*^/��z]1��^�h�H�EZrR�%��tr�9*y{ly�d$�N��G\ݐh�w��}�f�룝���VjX�6����J{ߎ�D;�_jP��t�ʭ�̀.�uN�R��A��Q/�⴩�7�c�~���>�sU�޹�U�{���:�Z�b�<�#]�����уX��ꕊikO�u�6������[Ӟ����+�v�Dޣx%V*3�&�^�*�2���3�[���N�jH�m�r)37�z�gq\�5����E�WٺR��y�Hm��'g������j*�k�����\,������M~����Ї��O7����zJ�e/����HO�e�����y9r�����)�⳸�����B�9E���y���������q*�������1NoE���CW>M�I�>�Tltc礚D�y}���N�<
���f��߳����� �o�LOH;ng�L����\����3j���*����(�f�H/��\_�1�=�mzN�#��=y�)s��ՙ�*�<�UA�����pK�b˲��`:(�-Rg[L�t�Uv��t�UZ�xJ��W!��-���e�u��_n�
�>�x��bp=�*��īw��`p#q��5�kn"���x����-�'n#>��v��;���@���Mě>��p�� >��-�G|4�1���X��#>���O4�$��+�)�J|����a��g�7�>�������������<��'����$����/2�b�K���__F|��W_i�U�W|�_G|���&������D|����j�m���N���ۉ�0�N������%������c����~���%~��ǉ�0�I�~����%~���_0�E�~���_%~��׉�0�M��I�m�����.�{�O���d��ğ�)�gN���_e�����-�wO���?�d��Ŀ�+�o�N�����A��0���G���g�M��'F��Yg�܋8����y�!v�'�kp?�� h� ��!j�0�ޛ�����#އx����2x4����3x<���#�h�$��O!.4x*�4���0x&�,�g�o���#�o��/4�����q����&^bp)q����W�I�i�$����_�����#6�����Hz�Kc �}"������4���'����F�c�k^K�dp�x��뉛n!n58A�f���ww�E����ě�L|���a��[>��h��!����g���'|"�I�L�W�O!>��ӈO7��3>��o�M|�������x�Kz�K��/��/��?��i�걅V�%��+�y	��g9V�t�8W)���n��~�m�o\?�6�����뇷Y�!}�.���x������;����Vֽ7Q	 /��T�%*�,���j�?�h��k�t��:k�X!�E�9�5_^&/�,e]�^+�J�Ke]Ea>���V�.GY��+�w�(�&��%wY�-��k�O��Ei������0z^�;o?o?����ۭ�T��3dq�s�-U�.V��}�K����5/�k^�׼��y��B^'����D%p��[-����[T�9:�W����7x��S�\�3n��d��dUB�*�����{t��ݑ���Hrώػ;r9r�8R�9r��y�8�;r��E޺'G��!�Ķ?q����m�-��ݑ{��H��%Йs����[_�����bU�X�NS6PsѲ��yC�)��U.����j���^�~��Ƭ�>B��z0���4���eMڋ�g�\u�вz���#��!=��%ݗ4��L�˩&�GUe9��H��$-"DZB:�t-���P�3H�����ELi��I+IHG�'c�Ja9�I�!�H:�t)���$E�?�hңH)�s"�Xz��I�Q=�I�g#��F��H!�2��UgZ�r�ɤ�E��@ZH:�t*�VR���~�Nz�*�^R�����"}�t6��HJ�9Ԗ�����KJmiQ��5 -���Z@��Iu�T�$�<�BRnO���{�b�i��g������m?������>��KH�l����}���>��������~�"�~ZJ��E}���:���uT?�j+���l{=�J�҃I'�8�XRjk���٤4���R]�e�M�<⤷��#���ʴ �y���R��L>ᓤ�I���.|��HR�[H�u��"�?GZ���H��;{����"��v�FF���(?�7I����/��!�|���G��H��P{8/�3�����~NO�����|�����$��E��oW���d�����|Ët��"��{\��|e��D��E����T�.��H���&#io��H��q�qy4�����9�r:���7�H��KQ�7��)ҫ�j��|�t+��"=�������4ҙ|و��q|���5��Dڟ�%��=&��mD:�/
���{E���*i5�P"��渽vX�I�������*�w�*���W:��t�;X�w��a�^J�v�wG(���t_w�����c�qJǻ���NT:ɝ�t�[�t�;M�tw�ҙ�,������q�*���W��=@i0�.L�EI�8醒nI�]�t'�p�]�tK�2��ܭPZ�V)]�V+��5Jk�[�t�'�I���{P�]�tN��$����*�F���ېt�n,�I�k�nSҍ'�uIw}�mN�-I�5�&�6U�n���Si��A�Fw����aJw�Pz��E�Q��J�q���X�8�ǻ'(=�=I���_��➪�4�t�g�g*=���ҳ�s����]�V�<���P�O���)�ؽD�^�^��
�J�W�W+�ƽV�u��J��ޠ�F7��&�f����*��ݦt��C���J�t�Rz�{��{������G��Jr���a�����)}�}B��SJ�v�Q���������辤�e�����)}�}C��[Jw��J�v�Q��������~�~��c�����)���B��WJ�v�Q�������������g�����y����wk���Ж��-_�������0_���/����Ǻb��!7_��V^��-7_�k�o�觭��b���A��/�hkh��������*�õ5"_죭��b_���Vl��Ř|1���q�b<}���!&��M열���<ݢהx���'���W<o/�#����=M�n�o��b�]&޶kĻ�J��(>���'v���>B|a'��O���������'�z�}��;K�a?(-�	i�/H�_�Y�k2�~S���2�~W�������o&�_���7r����ۑr��%G:���c�ar�S �s����Qr�3VNu&���$9�)����r�3K�s���|t���)�!g�\�,�a�\�:U�܉�Jg�\꬐g��u�e��Z�pb� �I��U�&��9ZƜ��Z�LwΓ��%�չZ�9I������f�y��<�yE�t�c�����W�D�'y�ߒg�Q��ϓg��s�r����?Y^�%/� /�/�W���U����*y��I��o�I�&y��hy��$�����?O��D��Z��O���;�C�����G��g���W��n���#���+���'�"Z�u��ߙ'w�@���p�� 'ˏp�����b�%Vɯq��W��I��m��$ã�.<	�	�灍���� &!�<|\|
��+�߁��Ɵah `D�� ��al`<�L��`R S�8������07p���f����OM�@{�uɯ����?2������E���ON�����y�> �_��I���Iu��6��Շ:��ͻ����tO�x:��y���t��x�t��E�{���:O�{z��+==��O=�y��ӵ�6y�t���=m�t���==\k��.�yU�oZ��=��t��՞z��z��z��fU� O<��OGz:�Ӊ�N���S�?x�����2O�=���O�=�ڳ�k�n�=�����ڳ�k�n�=����ͪ���YU���O�v�ͪR��w���iUz��[X}��������r�!3�Tޥ�j�:��U��o�wz��>���=���>֮�bb��&]��y`��R}@�C�5r|��L/�����dN�f2��M�T6����lZ�t�<Ѷ�F��t�1�g�ٌ�O���R������ޞ�ʇ"�]�� ��:^�WY��C�<>o���S(�c];=���[{�s��;�ܞ�����_����/�h��!��<ϭrJ<_�;��ڜ@��VfZqa�����(�Z>Պ�.�������qk<iM�����5���ËV	�d��Uk)�a-���U�ӊC���X��]�8x�:>�Ά�g�s����	_Y��֧��|g�
�	?� �*��71~#�1�'�T��}>��g�����h���^b�/O��#�������3|�V�q�o��ҷ���W���K��}Y�-���{7�R���>�Yc�򞬬,��֖���c&d�]�_@Hy��PK
    \O�H�9���   *  0  org/jnativehook/keyboard/NativeKeyListener.class  *      �       �O1n�@�ŀ� �� ⤴��� @�gX��/:���<�G!�vK�;�������w������]� �6Ly���p���0�,�9��_���$N�Z���*�?R���tGVkV,�~�m�ߜ�l����3TLU.�0���G2����w��<�J�G�D���qA�m�D��n5W��߫�h ��stz���wPK
    \O�Hӷ�]E  ��  3  org/jnativehook/lib/darwin/x86/libJNativeHook.dylib  ��      E      �}|T���l�	v���F]a� 1$�2� 	4h`�$����}�P�`�	�!*"����U��>�U �j�Qk�����6ꇏR@4�sf��;�H��~���$���ܙ3gΜ9sf�ܹ������^��D�@��1�e��(\���ie�,�M��?����춮r������36d��Z���5�y\�k+v������:ƞ���X��d�2�k��z�3�-��ݚ(`�,G�,G����-�.�PφK��d~��Q�rK��<����
�����͞����*������3+$���Ӗ�[0�t���miP�b��eW��Wɲ����l��ή4i���Cyk�<���<��x�C^�F@�֧2̣ցJ���՞���6�P��[���Y��f�9�G��ղaE��y��Z�U�E���1�~��	vͣ�Q[���fțM��C�sfs��q��0�XJ]�oM>��-.�3kZA�b�� �	��8іr��� �Eŏt:�U��z��[�,n�
k�ñ|��V1��ℾ4rո1x;sO-��,0t[�RW��g����2�.��*#K#�h�+�Ⱥ���"c��Hv ����Q9��~b�E9�m�����Y�MLtI�$�&B=ъv�k<r�j��Z;��V�8W����ZW:��]#����m�P7G��s����ʪV�G�hu� ����J#��顼���l��%�$γ,��:�u�3��p��g*�H7�|�"t�q9y{CpT�Z�5Em��<Z�#&�+k��+�ML�e��fWVN� �S#��>d��m�N�t�����Hu���r�"d3�dȣ{Ð)��P�ɒ��>0�\���w���߅��.�]�����Rֹsec��	w1�yL��F𻶈?�I�/6i��4�Iv��������i<����ýO�Ӿ�/��N������';;��T@;���ƣ8��������{H`�;�g����x�
��C|:Y����߇S���Z{:�cw]���� ��X{z4@��kO��9�1���]n����x;��6kO�#�ekO߂	��1O�#6�O�r����\�'\�|�a���\O<�'4~�*L�&0���
LZ_��s~�!-.|��[�h�n��p�.���L�5&����rN4u���zO�{�� �_�Iב\�L�X�p�x��M���^���,1߲x�;s���<�"��N&Yl�g�/�;�!{��a�`�̟�����M�J���Bp2 Y��%�ĥ&H*<7R�t.Ht��y�f�I��?��� _�I(5������yi�v�גi��C&��Ov6���z�AH�hy���K	���Z2C�Z���7@vM6М�<�������(�l���(�㟯Ey�
�M�m�P���h
��	U�x�y���fᄯX]Ѕ6b^7�B���e%�]��@�?A�9t�)�]��w�B�	���P�v�9 �X��X��:��D��S��	m����bS)���<�ug'j�k�9����ߵ�[ ��B!J!M����i���ӽ���N!��(��e$����V���@-1�g!�S N��]��߻�jN	ca� L::��Q��(�	�¼���s�ٯ���
3�?D��(���'�A�iLH3�ܥ� p@tF��].t/�.�.��l�.�� �g��s!�p�s�6�K{����Βz>�-��2*�;�����}�]���&�L�.;��b=4F�/���R���XUNcUh�+�:x��t��o%���O!��\�g�|<��8ϟ��h�����!>��v�J��D@`X�	R�$��|ky[�g3�lN�,/�� ��{
o�@��vw^N�@o0����@���
���6=�MVx��������9�qjō�F��;�Hf������4��rU0ST����Н�I��+2��^��4Av��H��T!���4)e�SQ���t��|�Ŀ�7/^���s_���e$w߇z�D������M�Q�Z��Y;��(�Wi�E���(��'!�ol4G�4"%����)qi�PV_���D����y��㤬�{�(�8)���ʍ�W��}�)��Wf�6�y�>����g}��QO\�[��ʑnmZ�����c������K_:���Q�ܓ���d�N\�^Y�]'��	v��D>	̓��1�C�e���)�Ƞ��`X�)�P�A��jR}D+�^Q�q�����7�[����䏻3VN�U�a���c�yI���$q����Ac���ٔc̟D(�E�Ȋ�DV�'���&�W�*n|ei�m0Mi�o��N���r.m�n�8Ō.(d��0.MZ~/Q���D����F-� -�I���	�2ח�C-���|B��	Y˜�,5Z�/(���%Z�4��V��s�d�����Jv hްH<	�����ڗ����$���Q	_�p��R�W���� ]�w���[��<�pu���yp�8L�n\�/}�E��Լ_k���QG�[f�;E5��9���)�Oɣ�)e��}]��ѷ<�G<�$f�+�Z�Mm�V�+^�M�n�B�JwwA�z���Q�ĕ��>��Nr�L����ŇY�}�%�8+����zVWφ}�A�Du�s�9GOi�(��u\h[r�b�І��>��|�,P5�>qL�v����x��g��|����<5gٱ^��~���{��Wx��L��x�"���/ͣ��3��U�yF���&����3&�g|7y�S��<��p����Ly��<��y�v�g*�I�y���L�&�t���gz8��n�̤<?�yf����&�ʳ��Cyr��.1�E7h�4jn�-�������U*g��o�oĈe�Tu�4�M4'������:��r�~�k2���	!���W*�Љ6�E)�S��i<��d�z�*t7��[Sy���gz��"dm�t-n�Wf�'M��N�F��Q2��=�_ʟO3nx^u�x�߄�����uZ��1X��
m
�n���H��U������n���H���σm|!u?��t����џ��}5������Dp\�e��awY�O%�,L���~��d��+d���tW�w�����@���<ˉ'_�L�Iyf-��F�^!/)ߩ�
������|��@YԞ �h�V��fY�E^��r�\�T������{6�k-_Ƶ�2.�L����*�+�P�lh�qЂF�p�%�4cI��sfx�=/x�x&Vu�d|���� �����<[�S��W�|q'���yBT G�Xk��F��|>h��E���g�!�+m��� <PDD�'��V1\��F��V�CH'CPW���ԧ���B"���া��D�^�L�N^)ƕ`ք�t3eND�d�l<ۓnޟ��;���u�Fdn�t�92i���]_�n��V7�̍ȾX�ͪ�{�M��H�,�������%����u�3������T��Y7�gz��cy��Y^������5�_�ͦȤ����O�n�t���y��u�w�'ݬ�!R7����������&2�IY7��@7���M����dݘN����H�L����͏#k𺤛�IGd����:ŏ�>�>��.�W����,��X�㠿��ɳ��N��.��JH�n�ϓ3��9��ߕ���+�����<�����������Y#̊O��{B��X�i�%��oZ�����6@-�)d�-ӧ�O���K����0[ａ��?��It �b d���ޏj�k�@�mf���f��0��HNyH�+�odv��^�)?�L���Gy�o#Sc�:��?�)8u�-в<�x�����@Kkd�T���<��љ��w#�0��@KBqD4�#��]M<>5@�^��%��@�&�i� a>�&r�Gt��8[R�No<5�s]�ejd5��(�fƊ2D����hY{�b�7�&��UZ�L$	JMe0�-��G��_���=�G������%a����%�j��4��F��V���h���`i��@�tHC��"�-�M���������En�-�hkF�׻(x?E�hA���_WR��'v̀r�>nx{��]��Q��P���,Bj�l�B����cB!b�>1�u%-UE�U9������NcDb������1\V],�h�<|�5�'
��$(a�F�{�߈�^�_xc��{$���W���̀���qa߁���3Қ�q�38oܷlY���14���%;�x~�n�FeL���� ��->��q�I㫦�hْz>������o�cC�C��p�
������V<���>�_�|�	݋e�t���L��wC`�r1��.�q3������4�	�?�������C"���d�D�I��s�
����틘i��d1���G�������h�M<�$�h� ���s�"�OP�՘lB�C�������<y~�΅�M�f�%�W��®��r= =F�١Y�~���:���=^������!o.~e���@��-��1L�=��,����I�4�U�)����7��~%�Yi�à�:���C�qr�u���Ϙ��u|��/�.�� ��v#�I�ؔ�%�4���k;�]}bw�������u��`|��8�Iܔ�P~H�^��>�5�lC�m��J�6���-T�sEgp�nC���Sp&�fw`,���:Q\���3����U{�NV��zT��A��}�>�)���wt\_��)P�.�}�i�L��K ���	�hz��Otp���u����^��J2��J��^�
��kO�Z?���W0���	9���`�:Z�ln\�6��p�c��nI�|���?��7����SOl}$_�5rO��Y���#����$��34���T���|1��R���9"��#��[�C�!��R>��͛��N��(��������%0�����x�|u�khk�� �|kv��;6"�������S��W��L����ߴխ�;�y�`�f�фj�k4��G�k��[��@��am�+ik�V����1w�:G�~#���}��1��8d
�U8tQ�X�z�D}�Vj���gZ�`��]ͯ���b��#���U�Zp.���ۓ��5�������d`|fߙ���<ľ$>9�Q�M�M��� ��8|X��^|�/V�w:8s �t0H.�ͪ� �<���3��]��7d�z��W��,�&u�^�m}t϶2.��R��:+(��k݂����|�������; |��<�N��Q���+@�{xsl��x�'��Ӛ֡߻O��ru�0��I�W���E�I��=�/(�:�*�"��o�}s�,w�_��8�:Ԍ�H�"7��4cMh�\�ug'Dm�)[�2���|Z�+ ~H��8���7�P�uX�*�Ak!=�
�.��'dP�q�b�˾����bu��cPU�!�v����&l�Ы_~����ot���a\zp8����Հz�v�+��o�5���z��0np�5��]�B��D������~��B��R�.�;�^w-%Y��vBi�e
����x&���&g��{��l_!�}�S<�����T/}�I�\c�����-3���f-UD�*?\d�h����lM����{��#^?��/��GF0��%�{$Qg@ׇ
xnDB��E1�w���ـŷJ�`�h?$�	�ll�	@��JM_��׌���[��Gp߇�?+�|c/����
�9��B�se�Ͷb!�]��x�����{7����[�t�W���cg*�wV�O`�^.�?����&}ۉ�w��M�#a3�i���BjN<k8�u>����Iz��]�e�m*�5v�7'�/�I|=��<;`z��f�_}ӫ@�Ǩ~���Q#%�
VNk=��)x�Kp֒3��0�����}3b��+��ȗ�X�A�V$�L�.�o�Tڈn������7,���i!����w�P��#�.QQ���A!}[�
�	��8'��k���k�*�ߥ���=���&�OO�>�|:����4br�2���^����n�L��R������U�y��;��������� �������w�(`�.*�+�^�6�Y���{��{P$?�_p��zRy�m}c���ۤ��Q\0݄,:���I��VJS�P�'hVw�G�(�J/�#����&�c�bN{�+T�|c��5��ت�OadB��J�Є~�Щ�*��c�H֪�c�䄎�1��Ɇ��1��*ɣ����X8���pY����韞`%���ܧVdF�f
�w�8#l<��1�0m�D�4��ud��q%a��T�����QlT�a�}v��$�3�tp<ό���U�4xw\2�0�*���%��2ݪ��ƥ9�4�C\�ϑf�B�ɠx4_`҃����KěMG[Â?�{�ܩ��Ԣ�V]�Q+`��ή�ۅ�@Y��d&;����v����90�4ae�⦔�J�<䀧���M0.���{5�TK(� �_�ps���LT��״*���uɂ_8��}�s�I�*���)���>�2����-��;n���� |}Q���;>7T�w>��.(�{�02�f�=[���]P���S�MÛW(N��{�������h��������[ZH��,�#�cc�4�{Ǩ��L����X�?Lc7����i�?��:�ۍi<�,�4$�����4��xm�+<'���i|H���~(7�1���|�m�祉��7W���J�Xx���K6W��WRe�U�K��1c�Ky=����5���e��?��0�mx�7R�2�v�ype�����U׬u|�����)�FL���f@�� o�ѫă_�U|�m,�UWa�k��	$���~�p�I�/b^��+W�ߵc���\�*�,��+�6�J��6�t~�m#ֿ�� �߉(�5�Dn�a��bAP�	p�ġ��w�������$⍪��H0u_v�Z��nl-�e�F"������BV����t��%@������^O�-�
T�0[���a3��K̧�GߓM����^�Ɔq�`��q;���s�B[*��yy�2��o,P&�l�n�4����`�`�	�����~�^'�u�nͭDh2Z������_�/P�G�x���wuQ���u�f^T��lO���ˎ���;6�ܽ�k
�=�ދK�~���ſxl\��������X��KM����<�I�W�� /�㐔3������SE���<��m��4�s��i�È�w��!���N�+(����5�y ��P���L���|��>��hL��Z|�7u$�~n���8���l	�������_�����%!7�����������C-iS�'k�1u��˸��հ�q۴v��|gD��'H�K"�0y��|CD���K�ƈd&O��5��<VJ�s���U֎���G$�)������˔zk����	�ⵒ|sD�̷XY�QH�F��|?D[{�K"���� a5�?j��$�S������R��|��M�'2�tC㵪1������	� �eq�����o�?�[P�`��d����`��O�����p�Jy��Z�}8s�Z��F0���Q�kQ�i�>O1=\�.K-�U.�m�ST���i90I��_=�2{)S>	Z/���I�^7&�E�6��K���(x�>�gg-�_˔-KYj���$��@Ki�8��v�9p��̭q/J������:=����/��v)����"y���d$s�L8���� �E<
���.[����+C����y�N3�#sB~���7p.���	Cf�*&�������#�����s��}����� ���Pī�\�Tƪ�0Ce��]�[��/F�Ph%3E^w1FnԶ�:Um)Ҕt`Χ��Q���'�d���*�է�{��y B6���8醗G��l�H��F?�6���V"|s7�E�3A!��Oke�|��IPM��>��*C~a�1�eK�T��H�w����H�} )l�F&��d�xz 4ҧzo3>Kpw�/�F*����w���T�RO�"壁��x��v�@�X��/ZNRz�@���-��#���|M�����_A9����$6e�@�D.TR&w�g���!I�� � ,&��)F��m���3�Ф��N:�ǹ�3��k�]�~��R�Эs��P���$�;�y�.��E/��c]/w,r����2ż��9:�	����HQ1|����� S�{��	��'�j(��l��k�d?l<�F|j(�sr�J>(���W�Y��}/��o�|4f?�)����H�]k��+�\x��▅3ɚ�4���D��Y���gH���M��U����n�p�8���ƣ����߼$����ac����濭�	;���ai��!Y��h�)�=��"��%�O/�!>�lB67ʹg��#'�#Eqb[K`����Aj���m�v���Y[�F���1�#F���Dl�5��a
ճz��oy}$��m�MT��&��I��p7������6�'�F2�wy`N�
�MÝ��ua[�0P�M����g�Pҏ/|�����䚟h�����'r�v���G��O���,0�l�^+r�m۳�k��J35��F�,��f�	�Ħ�4-�xZ�߸_���틳X��i���m����jW���G�C�]�SN��_D�;�?І�n'�U�����Ň�����^�9�_�_������ܩ�0dh|�H����4y�W���+�/_�0���
�>A�K�SH���:�M�����z"	���S�����G�^��/�+�R߿ؔW���U����P-�:� �ݸ���� �x�~����	z/�'}�����]��;�k��)����v�	GD�T�j�gQ%�@���O�[������������r�4�W;@����H+D8%a��_\6-����Vt�
^�w��t0�����R��T��p)�p�e����>\Q2��n�}���	��y��"�Y^��a�҆n�h?�<�v(q��/�(�s_�\uz��Z%��<�cR���#��V�󩏣wt}���	������/��h<s������εg�L}��G����xh?\�fA�� �G�~5?��o������4�7�7w����R��(�Go�H~�k�k���v�d��Љ�k&�Mƽ�xdWJ �6Bxd��O�xJ'��\���b�i)/��`	��ωp]w�!�"��=ʹW8C%�	N�������8/���܀����>.�͟9��f���<��|8�$��ɝ���$����^�p�_�x]�]C��8\�Oe��<.��.s^O��D�nc�"�!r�k��9C���W��z��wS/���et�~z�K���~��,����~3D��eĶ.�|�W��[ҋ���W��W��ے����A��H��׺h���w����{�������ի#��so?��p�CE�}���HR��$�~s��cC�������34�_Ճt%��
NI��S�N����P�NG�ƶ��!��I�t���$�N��D;���ˌ�v�E�h�_0�C�����P���M�7�m����jۤm����d�B_��ze-��n���������&o������y��{���|�<���`�r_��M�D��x�!Ͽ��LC��ChG�8���:�k*4�K+i�]�Zk�r�ݧE�y��Ң5v��?�]���r��C�}�"3��Rd΍�9�4\1�6)��[M��Z�W'$�ֆ3!-4N��&2��xf��2x=15�oZ���CT��Ӑ��nвiв-��6�G�Z���԰�E���;L�;�@����=��*Z�'�q[�L�#�`EQ�J���V�Iy�򧅃E�L�,A�P�ş��Ο��)=�S��'�Oш~�+�O'�V0X�Ӽ����0D�Y��Oߡ~ڏ��*A�ӽ��fJV���`R�觏�9�O���6�����V�pĕ������1M|�j$��{P�_]3H��]�&=ү�O���[^���'�;��o�uq��*~]ï��į��u=����F~�̯[�u�>Ư���v~�ɯ������"����~=̯���Q~}�_��������� �~¯'��+~=ůg��݇W-���5�_��ʯi��ίF~5�k�f�k6����8~�ȯy�Z����Z̯%�Zʯe�ZίK���_k��ί�����U���_���_���z~m�k6Z��ឌl�P?�c���:���ؘ��	�4����aCo
�7tP��ȡ��:�C���G���$pl�нG�%p4��S�h�j��Q�n8�Fh���@BS�f#p4��p��Ʉ�8Nh���|B�G#
�y��hJ������ѬB��+����B{�������B?8]��G��
0t���C+���U�h��%G��8�gh���HC����8lh���lC��7�G�h¡o�r9��ќC�:���ѴC�<�����C�	�=����C[���_�h��f�c'�.p�
�:�c�U�E�F�c��8v��d�cG	�8v��P�c�	].p�:�~�J8v���
�G�o�.�P�رBo
�W�����~�����vKݲ��v��5���?.6mU������t��n�2�F����+N� �x#����Y]��2�2ĳx���n��n�2���3ZWX��F��z��ƌ!�ˆ�a�����0��檷�+k�N�p.��	�vG�ž��i��1�)�qZ-U��;B��+�|��"xy,#&��QTW�qs�	�nd���z�s�g[k��ӜN�Sґ�NZ�z�r�����"�����M9�e�E-�?���$"sZ]V�
k[ �j�	E3���2����e+Bl���Vm�:]1��[WW8,�**c�u5�	��'��wTY	-v��TRj,N((?�w����وˬ���T��-X��m������xW��E=��j�G2VX�I8��)�
Kq_
��w<�|�[TEj�[��nV�p۪WC�dk?��\Vw��Qou�WG�Z0N��F�J����M�L<���G�˖A��b��{�B�u�)N�	��Vg���F��v��Y��_�n�2�g4��k�r����c�1sN��V�:�-�Vc��㪃�auO�[a������<66�YȔ��R��>Kj{5?'��-����[-n��bư�F�����rU{�Y�n�6r7�mf���3�ut�,�'��E�u�tԁ�F,�(h�H�i�7^�&1>z���V��Y�������y�%���-���g��,�Z%N���	�RdfT�nu�nh�ƶz;��s�"qȒ9d���1e5�Y�j��R��u��p��qث�Ye���.�9�媐*խ&\�:��gs���+՗r�K�%�EE#d�[;n�J��n[m�K�Z!�a�Y6(�ꮂ���ɍX�w�]���C-�j��,'ǈ3-��Yla���n��e�0��2ZW�QCP�&<�R��0Y���Z��gIRXu7N�2���Xi��pf7�o�;V�xU�0��v1V;�s�\��yUV�[�9L=Q:K}�]���;��.I��:�Qot9<�JkV�4��gN�
>#tf�)uFO��:��:^-���FGe���Vɜ�mc�5&fy͒	��)6��-fb�5���C+����W�ds���][>��b�k���E4��ֻ��e*�U���g�B��jYn�բ6�ݖc��4<�d�����&o���xJٔ��i���a2%L�HYg]iT���4��C�=�L��
��$R�,����U�~�{ꊱa,����}jA~�2��dv����bR��΁=ո<W��ݮ��+*��Z�y_wx�r'We*࿈.,t<ԨL�@>h�S�źk����f	��Z?L�2En<#��hsQߩR��'h�����E�>�RYS
d������2"Q��2���r.��%�:ܾ��u��j5����ݣ�Vg��c�ĝ6���1���6�CG��B��-��`
�3g��u9a����%����%��xb�]�xj�>��h����
O%�֫�As8��Tj��dݵt�1~Pu�W�d��nn�2�G��]Z�g�Oe���΂�Z�	��vԫ�T���zX]���_/ܗ&�fJ����yx����y�@��R%*�ʊ�aa߃&%WV�3�s�J�;+�1(��hc�-�'�y�8�Kp��%s��%Q�^�0�����*��{4�Z�6W
b�bx��HA�g<sy*�b����H��'K��Z`t�qW�<�
����mF)I��b�O�d���fG�ϗ\�P\O&D��V3(��"GTɱ�R9�YZ�E��e|d�Y�*!���T�,Cm����+q	E1�L�S�l�@ln�'�`�s*='�1. ��&9�8�F���,�plv>�C�7�<����9�{(.<D�d(��.#��)�[����`����c�R��,�8-�z�Np.v��\�-�8\�8��Vp���|G��-v�Ua%A��,v5k�O�,���f�"=���@N�^�c���#2����Y�Z�\�|�c���	3O�l˪�V0I�l\��S�P��h��SV���R�L��'����/�3\cW�Nv͌l ��d�Y*�.f��Rv-��e���H�?Uu�fW0���Ҁ�:����ї%�~,��R���pLN}�{��)PZofb�	�=�1�� %$BiIP�J
�@5���z��b#�8(q8H��r��(������z�tH��H����Md��ˇ��?r_���ưUl\�JvE�@��U1[�* �bc�`-��f�;^6�-b��naY�ʙ��6�ߍ,��M��̈́T+�f��o��l>��eSX	�a�b���f��	X'+d6VĖ�;�m��wA�B�)&�[�T��N8��nf��J嬓�U@������~�lF�%���!n.��(�	(ӱN6BɱŬ�����<	���?��b����O�cٟ,"X�f��O��tA����� �� n?��jxШ�~�%~�wK��X��eR� ��A0�@�u�?��<�6Ȏ݀׆��)tЂG=pO�� �h�Ϡ?��q�HCw�@�4���?ñ:[�gl'�� l���c��±T�?����~v^�D���AxB;�W!��8��B���X*#�L� @(�P��B��6Cx�N/B8�m� |�-��B:��� C(�P��� l���v�C8 �(��!!|�ff�!�	B6��
!�BX
�a�&m�@x�3�!�
�]�!��p�Qh�c�v��>��z�6�����e0�����aB��4�O��K��CQ��t/�2��xd��7ѽ�i�*����Ϟ|bԹ����9�\i/�]���w���߅��.�]���w����w���gI�g�"x� s�L0�� �i�$h"8�`6�1'�J�����o&��`5A;A'�U�"�D�^�m7�B�Q���A���!�N� �W	�I�]�<N�oO<I�,��zu�L%x9A#��3	�"8��d�g,!x#�r�k�t��`�f��	�Op3��9�g	�#��?�+��	~C��m^L�j�����4��.&h#�!��`���B�w<B�����OLr
؟��Mp
�������}$�#�� �k�/|��C�NP��/��!�Cp�"�	Z�\M�K�>�?$�s���G�5�$�W���� ~�vHp�56\Gp=�6�	n&���6��|��v�;	>C�y�/l'x��a��<J�m��|��1��		~B����"x� ~b�PKPG0���`*�4���M3f�&�Kp���,$XL��`)�2����"XC�N�����*�k6l"���z�m7����n&��}�<hW��M�8��j�0���`.����t_L��S�����4��}w^|"q��>{g�6�K<�ؠٙd0�Hة��6d� ���׶���6H�[zTמ؞�3�]�-�=�����h�6I8��W'j�G}�ވ+�Yp9џ1������1��Ѩ8�g`���h&�z�^#�^E�d����}q��9P�p��$O�$�1��OlM�+�}�D�4��t�G\�_!�+x<��kT5Z~|?�W��MV�+x<��$�;����=����#����G�༾C�J��P��Cj/���u#�;T�gIx��o��=�!��H�>QŻ�;~n���غ��U��.�+u�&���� 4�DB�����K�m�9ȹQ��Gq�\:����\�{��6�����dz������=�
�&�?�x��P=c���.iU<]�.#������ޞ�?Ř��W蟔����]���8�����?�
�c�c��F3vE�jt���s	�#��oOP�\���$U�=�Ga�����yc}��&ǩ��<Iv=�O�+��=��%Ƿ�	ɪ<	�+Y��'I6#���2Je�K�Upn��;N��Vҕ����)�G\�ϓ���@W���z�G�@3��'���<�M�y���@3�r����^ԧ��5�*�~tS�����?�+V�� C'�S/�S"�S"ɏ�R^�#}J�]��d�r��0��� ��Ʀ=�
}{�J���?�g�&�G\��&��6�N�B=��p{Ic�A˘��#�зI���\����W�_ڳ~�"z�{���yB��Do���4C����_��:��%��:aK�-�����#�8�W�W��<�p�C���Lx
�N��7�
��_��O���ᦇ����U��ޱv�t��>4���V�U�����g�Q�>��Y5�d�x�n%;Qpޏ��O'z�{�o�	�a�G\��)��賗3��#�/ى��~4߻���Do��%��Z�*&�{����=��~'�#�I܇b%�c}�D��J{��+5b/�}���c��ӈy�v�q|Q�?���C�F8v���c�ԧ��'�<q�_�lVL8��r±�-G��E+��f�џ� ��n±?!��;�c�+��� ��i±?��8��k��8�p쏅�c��p�6±?z��x����g_��x3�8��)�8��o�q�tM?��<�f�!�:�V�a�XI8���>��p��#�c_��p��t=� �x±��R���/$ǻZ�q��H8��V�qN�^ȉ��~C8�C{�pܗ�1����k�?<�^b�r��%�y���S��g�Z��9�%�U�ar�#��=�U� ��B��?�%d�}u�"�W���hp.4�?��Q��s���=�-L�x��	��[K8�͆��,ܻ��p�׷�p���W�q__���}c�}~��-��U��^����s�_�� �����}�7%�/�����x	�R¯���^#�wHx@�"�;%����'���~�*�!�$|���H�W·J���_�ߓ��%�],�G�$���U��$|��?)�/J�%�S	�F��t������n�p���1��I��%�]�ߒ�?���~٥*�+���`�~�8n�|�!��'p~��Ϥ���K�wK�~	C*�c	?%�4�V�gIx���)�%��4U?�MS��i�*Ϸ�|�Zǋ%|�e*�	�#��J�{��Q·����5,e;�	�J�}��<K0�~�	f�ƍ� �O�5k�y�� � ܫ�m�!�p�6h�s�}�� �E^<vy�� l��C�����s�y[!��{� �£���?��4�g <a��!���kļע���Vo�p+���j!�Aph�s�m�����<V@X	a��n�p�5�;!��n�B���0�s^���	��j�z�/ ��~�q�Shۉ?�E^h�����F:��*�
G�+�p"���m#��3��$�3��������[y��Lf�"J�]>?�(2Z|�'��5��� ��C9H���c�t��ba���Vj\�C���u^�De%����8q^�yUVɢ�@H�"���r;��q���O!]I}�P(�u����!�Y���3�t��O�2�Pf:K���E-e����'��K�����&�9��<��|a���ݺ��lq�-�5f�s��GPQX���sP��Լ�8�
����j��z���-��#ϧ6(����ܹ�-T|��dgg�ʍ>f�N����ӷ��� ���nݱ�VA�o����rI9�,�����1����������!"B|֬����U����̆��\c��g�#X��]���n��Qe5�fO�ш8W��ND*�VZT.zS]�H���D�@�'����;�+TWh��vx���*<J �(�*�CE�KԆI��.��1wy��9��s�c �]}�o�b��^^�q�G4�b=�Q"���e��㶮��+uP����nv�y�,6��{~��3��1 ��Z�m�'nj���RT��'�D_��ڃh;���t4M����Kl�9&�M8?��>:�����Gې�mC��4U�cD��������I��~5����{�T���%�?�WSc>�7�8M�,�y)B�V��^��0���p���3O���q)����h��O����vn�����k��W������ƿ�)�?֏��'�&"�u&=���1��9u�n<@l���q �{��bG���)i��z�^�N��y����{~Ȍ����ųC��q���>��U��V�Y`��b���ⅻ�*��8���sw�Yu�|���Ӹ�l��CfΟ^ 60�Ꞻ�m-q;��bk�2w���ZT�#l��;ha�7�6�ŎH%�	�����0��c��d:������VX���Q�h#��w��ϧ���ᣡ�TU��r�*�A�u�`�C�$����l�^q�����|���C��$D*��[�h�8���1�{�2�Ӳb�����h�q÷7Y�[�qf�`3��g;89��
� `�'�[*w�q���,��@+E3����Y�ݨ?D�ɽ*"A��.�#J]O�[�{�E0<A���2�f��KMTݺ'�6ݗ� �Y�^�Oʶ@̻"R���#�ʑ��S2���õ����a� ��Vi�V&���)QI���֣-��fUT�*�-�l[i�b>��.S�1 �G�O��$)^���a��R���4�$R��"�
�`��Ǒ�ʶ��v�	�!�87
�8��gE�*�U�rUv�jɬ�l�d�0J0����R��p��<�q��Y "#��U3��VK̿���"�T�#�"6ܱ�IjJ��)�0�R�+&���Ud4)~��/��{I*|D�FU)�]�r͝m�ӏ�˪��vQi����x����ӊ���I��ڌB鎊[+��W@�ts�V|n�w��0>Ř+�0"AwGů�ؤ(� �>b�q8�a,`V�p�c�	���t�a��PK
    \O�HW�w��H  8�  6  org/jnativehook/lib/darwin/x86_64/libJNativeHook.dylib  8�      �H      �	|TE�8�&�	�H&��p� 9��!�L�����dBCf����&Q�������]�ؕݯ
^	�ꢮ.�Ww'�#�r�8����7o�L\����>��UWwWuuuu��^�����~$I�XI���:�M�%�YJ��w.�1�d�.+�X&E�ڢ��S�q�?��k��eS�+����B�V�W+5(Q����Uz��fgp�&�k��_\?k��᲻��;\����ӯ|U���~M��\�`��p\�b�Q���xx8����kCx��"���7��W[��k�Q�}��`�&��e
�g��ָm����;q���C�K�E>E�e&E�����8�[l�����V��_��O.�u�����K��V+p%?�7s��f�l^_�tX]^w?�����ni��wb��y�5���~;ng0^�+�������^��.�]*~C"�U�(;��_痯	���G��kS�����6�?�*��������q~�4J~J��+=�0<�_/�w���*����3�,ZX\T"����p|��R�J���U|����fU�78]����6o�{�ӹ.�QW�Ums����4�"�E�1f�"�`�����*�G O�Iz7�� ��Bw��T�r!��r��_�I����ܖ�^+ ���3���_����y޽����ό��:fy��r�M�g�o�x��,u�n�{s�<t]��u�,��娫��9����uUvOf�H�Zaw{ �E�H�U��7B3@y%��y��@Ir=��n�P?|m�Jg}t�,�����L?>���.g�ڪLo`�S�i5�:&Zf��2�<Mݚ�*�'3'�@��Uҍ�;��o��n�<����Z�=��V�d�^�G������3����Y��,���~:����������������������a?S��5���`�T���k$I��x/���:���q�����KROb��S�'b6��y��Kr:�uҞܮ �����8�X0�I
 �3���v�"� AUS��?���i^w}Vc�?��o�=-�.	Wا����N�viR<�̍�s}�=�mNO��-c�/x}��`.@����g��7�x�����vakp���5��t�ň�T���":�4,�Vfnl�݉=0�b�F!��R�
Ӳ���J������-�������� �g�`�����6X�sK֐��L7��.YF(Qu�6������FR�`n��Ҵ�t���9�A�t��Z�"��<���]Hܚ0o�����Y�[���v�m��_��%~X����0߂h&���y��6L�b\��\�"����͍��K@�V��J�	Z�ⳮ�����V�1j�ܡo�M�Yd���,nI4���p�l���r�1�ܚ|G9ɽ�nlӮ��0�'`1��M,�~��J�լ9�hY�P�ּ(��EonɁL��Q��-K�Q�m۠�����c���#��c���q�-�[��f�oh²�l�n"Ea[΃�~s-��?IK[���w.J2�w��E)~�1ɯ5B�i ��=�z0V+�3l����.!�����9������8Q��e4�������9�UF,3���BY6(�{qx^^��1aeL�O˨�2z4a̺��ʬX����~Ϣ1��Jd;o��l��m����������΀ߋ�oa8��3�w �}'����?�׉���~��7�R�le��F�mK
2�̐m�X,`�K�;����-��ٯ)x;y�>s�{��x�Ȃ��oV��}����Z��{رY�E�l��5&��s�<K�q�y%��}0~%���� �[p�:������!l��}�.���J�A�孹�K�$�x��q�27�o�0�$'�-&G���Dw����Kob�-��m��H��`�a�$5A�� <�`�$-��G7����i<�&�S�'܌�~��E��M����Y��f~��έf�P��-�Mǋ�8��!,��"A���|@�'��*!a㄰s��C�����S�6^��<��P+K(�� Y��L¡,9�^�K`v�c�"�ѳ(�#TH���S��t�7�#3��zdZ��r�\��KK������L��l�ʘ:H(����p�P���c5�ܫY��0�b1������DI�9����U��8�����Br""�l<S�ۥQ�͵6�/�@��� IU Sg��s��T��*;>��mWYPMe;}Be��Q��(���OVb�֢Қ}Li���g�Z&����R�o�	%.�P��������,!Eu�2��LcK��r5&F��y<׈N٥e�	u��s�ܶ<SL��y����FS�
�P�/E{eEϦ`*:�K:GE�L�I�]��H�ǣ��Um�Z�Y��,jŏ�
ſ����OşKM����o덳���OD����ͱ��[WD
M�p��FSh�G(�;7E|���[���e�}�2WT�)�"�rC>�x�ڧ�#8{!)p��}�}@��dn-��]��5[ͧ_�5�qG��O��Y��EB��>�����C�<�r�R�Gi�4b}��j�~��ÚhC�֫D6^%�����f�^�[�����|5�g!C`���z�ȸuA���h��Q�"�dk^�.��wJ̚�J��+�Y��L��zi�뉴�r��Z�Kv��ȔѪ�Q�L9��R��6̔�Ou��xBC ��=�Z��:��|�<�N`Go0hz&p�" �xi���>��.�%m�ω��S�-3��Ǽ#غ,ض���[���!ܩ+v����7 �$$[��F��F@v�Ȧ3���d����"٩�D�+D�� d� �F���4 �Z$���]"[9 ��HV�Ȧ��� �d����e�S��'{��\Bd�r������į������Skdl�$�Ձ�4݈��e�l:lL;�>{.�|�+\�xsk�|�J�?�t�1PB�y_���GHR��F`v9�����`� D؊��V���v6Z�W�J�"�!��X��^	U¼�S��h����'���-�|��e�2��U�����F�~�c�Ȥ������s�v�̰����1�q�h���&c��d<D+�&#.�:��O �fATn
庙Q�lݏ�쫩Q�g��}���5�j��z	4�IRsǦM�j��f��x��N���v��v�[�XZ'j�;A`���*_�l#���)����T��
\׃�Fn7k^~hi�eteI=�s:zjB)=)!��34��,���`�j�V�b�M�Ҩ��M��־����n���p=�.L�Z�0i�+���J����'�d��m�k�����]�vў�dr�e�3���E48�@�{�q�Ӵ�A�(�L�g��pz�5�$R��������n�p۶o�a�$��JPS����A�(�����o��ě��[`���O�Y��K������S�9��I������h|�m7�|#LmRj�lj;�(GAɥ-�t[�$�f��Q�?l
��F�8����Py�����3�](�D�|��\Hz���~J�&j�=��ch)��0W��7�#=�-���7��z�-<M=l�=c=��*{g�\�B7���CIKd=h�#=�N���k���@��J=��[�Ì�=|6S��?�����3��L�V�\Y�Ѓ�%�CINYߟ$=|���2�9&Y�(���$�!����g��p�t�PSs�zx��ݜ/W�v�/KZJj����	�Ck��fT8��z�G��gO�.ȏ������y�z��~�zx��}�\��;�V���Pң�>=Nz�3R�1����v*��?�I�͍��[�j=��t������p3�w�\�ׄf���CI/�z��M��hWw_��56�ǹE.���=�y��-�B�8��A�-����[s_�$|�Bӆàz�2��?C��)�m��@����J����Ǳm�~�"I�'���h5w5��n�	K=}�	cc|iP�3ɪ�IlVv��0l5w`������p
���u,�j�6�fo��lA�h���V�~U�l:�1�M���"�*z���VqO=`�#v>b�q1���,l2�{� ��XbV�X!bP���+Bl`>1v�l�̖x=�}��Ei&��µ	���b�n��Wp=���>'Qs��}�өX�DQ�VHE�H��}�A͙3H3xڪ#���}ϫ�Ï�����繫���,;��mۀ?x�V�1��A`dW���6�	��jpK����	��0���7� �O��o��n�^֐l����±M��=v��	�"Ov�Qnk�/��"���B��ǽ��%�=:a��O(�����^Tn5�y��=�+I�.5Y�"-�� K��8��s��߮�\򓢋,ׇ2D)j\X�(����91J�rb�r'�La
�^)�ʅe��[�5�r��]t�mY?���=���զ��t�[���a�����;�~�W�`�/�?�/,��N�ܔ�B�k�b7eʃm3y�]�M���-@v����e���]�$A^�7��*T�ǜL~�$�%�ʹ����$4`�'s�H���:I)��&kA������Kk¸U�3�C��佗�O�^K����0�_Iٞ�t��r6��f�5�-�-��y_;J\F��ٛN��wvDÞ��ĵ)��c%���и���?3����E�����jzI��9x+��s�+�]�F	�#_Vŋ�}�T5�zѷ �Vw)�-3<�N ��3o�bҀ�g@C3��dցR�������a�/~�ܒ�{i�1���j��t��J̖Z��AoR�$թk�i �w�ş�Ҵ
[}"m�~���ҙ�Q��7�!_��
�;p��_�
X�ڳ-��������: qE��:��MJ��}s+��'	wg�0�C�C���L���r�(�y	���;�NS��[Iz��mo��B����g>]����斄7�c�Yz}9Z��wC���/��t����N!-���*J}Ma��"ʂ�w>H��x�]hL�����i�?�g�l9hG3{'��w+:_i#���y0*������ؗӁ��6��Ʈ�p��F_�	)0��rm�٧�Ƕ�Bx4j��Q�S�Q��5j�>��@{��bn����Ι#zG������7\�s%��ʼ�;�g~m�Ҳ�S��̹����+��͚�������~��3��4�����o` o��__�s,��d������l4��>?����{�eԽ�fie����y��s�{���9j���D�*�~�b,=�{�k�?f3�?P�K�?�rA�[��e9����Ioе ]�����P���8R�FFT�D�b���DT��
���
��(����Vd}������� dlHX��<�I�͐Ԑ�J��ImHXX�3XHw%������Չ�v)�:�;��1/�H��,��ԑ�hC,u2kߖ�5��A����� ����G���O�� �N@j5�'܄�-	��nfyo������Q}�A�Y��r��ԙ+H�t���n�Ǿm�(��yI��E`ɓO����n�%U���@+{��1P����$��r��S�����kZt)$���嬃_�}0�ۘߟ����%�c�~�5�e쟜D>O.��I�e��z�S%�^Bb�ڎ������@��dp���ŗ͍���7�Ӓ��<����io:މ����:��o�C�����cYi%�p6��o�������/�yq��|���_���� ���� �O�烯��5^ߜ͸����T�f3{I�'�o���5vm<���${��wq�~�^��D�ߚ?���	_��Zj��/C7��˰}v�
�|�Ğa>��x"�`�eD�qk�ᗱ?Մ�\p����0l�edd�Xp/���]�K�5�4섦\xM�!�z�W��CFd�:�k�6�c>~�?V��>L>~�N>5��G����
��	�W ��`��q0j�Z�ݓ`�_�-����<a<����t�@�bfc1y?�i�om�Q$��� ����
�g]O���Q�W�W�n�=y)�i�V�KnH�L�3�A��#�=��� �)�>�I��O��������㻖���v)���qm�]O�!��4'�iz���xLXE	+)!�����PH	�)!�ga�Յ�0��z��X�|+����!f�V`�P�1@��k���� \��W�Q޽��+d��
2�-+��I<A.�C��+0w�
�b�F:���)w�,j�wf��G�|��1/f�u�xa\JHQ�N�g#+�%F��$6J��F����z* ��m�,1�m��zf7��9��g\�AMϹ��{F6���7L�BӐ��ƃ�����cˉ�l�/��ݗ���2��ө��ӅD3�X��F��c/̏R�#f7׍���$�ڹ5<u
��%�'-���,irx>��ΒÓ�ĤsY�W����k�v�އ��A��?���k�I����<�?%�1���GW��/#�Y����e��lZF�cZ�
|�2��(6_r��M^ƌ?�.
�����ǝ3�m�?�yσO�5w�7_/'#z�^-���"����6"|u!�2���l�Y�#������>�20�w �~�,c�����Z W\up5���c�z�_�C�*�)�'^|2���m(\�]0x�w��� w/��R�{��k�'���+����ʶ�upeC�] �� \G���;�Ɗ��ǽY|���`�m_M8���uK��KYs�-e�'@s��Rs/]����W���)6�`)枽T4�ġ�a�}�i?�.��Û{����%���F�]K���YB~�Q�΍�5�X�<�v��{��z�}K��뛮���u3襾����;��/��-�� �4N�-��hz���-�=����b(��iT��iB��P�ZRs���a���ފK�4��"���'��-Ȇ��c�[�%Y.6�j�v��{��6���INaR����i!Ĵ��-e��k�ќ�{"�҂��2|�GSY.�8�=�����@.&H������|9U(��PeZ��1�x���B�r�Cd����y�=t�������b���1���r����LW�̬{1;���%y���{S�-T����dTS|�?����B��98	���PȨ6-&�k��k�w�����=��$�&�߮&σ{�Q)�Җ��]��O-	���6_4_lJ��t|��(�����פ��*�}��MP̬�o�֦SRg-��M��lis�:}1�:��Q�9@2yص�C�8[�	�Cgy����Rw��r���e�ş{��xl�\�"��M������L��?��z��@�z��C�m]$�UW��K�L*e�)�-��/�k��D�Z&ՕSEKM��'
���^䟕R������CdƜ�&3_�~I*�?a�x�?���:[�^rNZ���@��o�_=�y۹���RR������������T��@�R��n(e�)*�Usq������c��f�����E�tTN�����9�|sf��]������������(�hc�����[�S��e{/+�S��"�7� 5j����a!��B��[�&J,�%��O-���R���k-L�̘���LLWT��l��@���Qi����A'��?�PQ�ܿ,��d.+�I,�"�~<�ܸ������Ⱥ����|����ϻ	�NI�#���3ɡ-���Qu���_��~������ag[�^#�j���B���M�ԏ�̸�B�Y�}���
��h��kʇ��j���/�f�$�H�RH9������hԐ�o��@4�u^��r�!�N�h<�(���o��@�%��}?D z6F�+G�@t<D�a�r�� zF���+ Z�a�er�<���	�̒�q�i*;A�˥C	��u�16h��d�y	��F���迕��G�9�X��ν�2+nζ�>/&�fAi3*^�T�l�M��� t�N�}��iz��Q���i�����ψvv�h�k�KD�a��U�p���*���ϐ�o�_�w�1����_S���6老��ğA�d��-�����wӋ���$��"�iK��3. <�.�}��i�^;�7/�<�
>���oF��f���l�����&�/��4�y�\���_X���U ���1���n�	n���2�?/��|��ŷ�ߚ�j�|w�P�C�A,1HB;n�c��=*�]�F��H|r�o�9n�5�Z���?�i���բ��t+ۜ	e��*,2�ds�z���R��h�y'm�L���a
�I�3�fP������o2�d�1Lu9�pll]f�Hg"�>��T�-LM��v����k�xʻ����ϘN�i�N���ܛ@�L�mD�X|�(Ϗ��=}���]��\>$t�}R�$����,���h�ȢY6_�Mt7���	�JK�w�3��6Q����%g�Rdzk�"�нP��O��*�	,dQ>Yf�M�D9�9B5㦐j��G����j��Q���$�ԛf��#��|,���,:�b��c�~�y";���������7ݏ	VB�}�@	ếcW� ���Mż_`�lU�1éԌP�/'wy�7�}��Ӆ�m��b����xbm�eO2e8��z��1/�Ht�tA۽�׭%��H��V�8���3��b=�Q�^�䩱!�wC����B\�ᚫSw�Pb��S�{d6?K4���԰?#�Qt	s6~�8-y�p��[=�`{,���$�x�&�[*��a�7��	l�=-���$���s��6���^ˍ�H�VO]�cS�"�������Ʌb$��gܜ&�s�C�-y����^���)�"9�OD�*��^����������30L��W�����V:�������O�����9d�۬9(���<��&��6��9v%���IU��L̝u͡�mb��;��b�D�ϴ�{����@ix�)�/� �=&V�&v�D=bⅸy!װB�9P��T�~cx��i�њ�
�V'���܇����K�C@`m�#���G�:&�|V��ya9���4Q���W�`Ş���D|��^>�y-��>���OzV�;�5���y:�������x�A��*�������|�d���	(MT��rZ�z5f�@.&�+��i$�<	�����%�Ԛ�}�ArAQ�gE-�Dqʊ:)���-~�n½��"L�'���;^d;�'��dH��ϑ`0_���{�O�?�<�~ga����;��zɼ��ps�m����Ƭ/z��n}�x۷~�%��OO���s����I">�8���m<9K#�[��9u=i/Ƭ�e}#�2q2Hݫ4bx���<�؁���/y� ����)L9�������3�n�'���w�q��S��9�`�f��?%��f&�(�`��}sn�P���P�ݓ)q���S��L�g&�`wߢL������~`�P�X�����$Z6�q$�d>$AV�*�Ɲ�7z��H�c	���/�����ܓ�����`�xڑP_�;�Tg�������7xx��`�����{&�$D�����a���A�s%��%x���j�w�J�a0���z��_E�o�f�,*���a��1��6-k�Y�����M�u{l�WM��ܞx��O ���,>X�?��$�N��B��B�Ӡҳj�g�� c�ϚP�Ό����4�W�k��~�j�	�� 6��7��c)� �n�����A�VAܝp=�p~�t*�����^-��i�Ԓnd�|�R�]W��S\hnIH�,�-F-5.��LJ�etj�(Xi������oi�����W�����������Y��B	n�8�<#�~ôR�y��)����fu<5P��pV���>V���~1��x��4�H��f��K�t��"�r?Ono�x��q�D��b�fh����t8�=�OJ`�ʽ��B��,��^��0㹌�t�<먟��{q�7���}�R��s��O��x<�G���;s"����h��N�п'.L��������F���i��=�O�w�1��+}�������?��HW���^��������gC���x�����d�Ϟ��Ӳ��������_G���?;��)՗���\�SZ��_2}ߟ%��=K���,��'�,�.B�_pe��_t\�oG�{����9��^�LA�r�L+�=Oh'���7����nd�FX�O;tT��uh���O����`�ً15�̽f}��g�������a>��������wf�����&RO���#y�,[�F6��}\�BoWf
���6ms����.�J}���\-S]��T�3�چ�j�����K��8$��q|3�$��8!��>$N���nK��DH+l�k\wv�C�6�B���;#¬����w��]�-,�1�uFX3���ax3>j�0� oƗ���j�`��u�گ�כ�͈�L{PѹӘn�H���(_�;Lʉ�_ӹNRƂNz5B']ٿ=����4���p�o?Ӱ�� �oS�E��.�fR����@���:�U���&)����x�Ҝ
���5�����P�گ@���_q��s2w�OH]���zP��F�g��`��4>��
���ϻd����g�>s:��֨��Ă)0�XD�yt7�}�-t_D�2�/��2���{�/��*�_I��t��{5�k�^K��twн��.������o���t���[��@��ҽ��7�}�o���t���mt���w��.��M�_��Wt����t�����wt�N�G����@�t�ݟ��St�E�g���wӽ��/�}?��� �_��+t���-����&�w�>�p+�W����X��fފ�9,|��Yx3��,��p
_��a,���a���(l�p��m�;_��C,|����r�b�%~��K1���%����1���M����0�b�Y�f�\W�p�-,���|����,<�i,<�cY8�I,|.��,����Rx8�?e�w��`���u>��?�§� ���Ob�A��w�����?�pwc���c����`x���2��%�E,��g���Nga|��m`a|N�=��_�p<�����P�y����������a�#�_a��c�����,�[og��0�+�5��X�7����·a��­^��~/c�f�Yx+���u�faܯ�6���)^k�`�r���d:l�"��>�P����O)̳�9�����pVټvC��7�<ۀԙH���D�a�D��%�l��j�����^�5x7���iϯ�<DZ[_g-��:��歪��%�{M��K�;��6Gy��n��0fY��n��,�e4�>n²_,U�"�<)-��Q�Ի|^�r��RHS�}��5���N��b���V����Z��\O�2#*)��9���K��K��r��?����7ث�r���Y/.YP<�ؽ%ER���:��j��nO�u�͕N�����о��	���rN]謶���>�"Rjmn(�0��z��c�K1�d]�Y��^ƪ�QW��lʋX�.�祵v�#��`&�t8L�K�/CD��:��*��\k��J�No]�f����E$��[�v��n��0���Ҧ�QR��ns��&���u�,�s��ʲ ��⡾9E��X����G�Y!�g�6�����'tc�]R|=������UW���e,XTb�����5�*���p�A̷{��7j�n��W��Ƶ2�
�cUڪ�a�g*�>DO���V��봺�.��kuCWL�<���UU�=��#܍����r����	�%�L���O&�	�[��4�5`��׀y1�}j����������Q�۹�?��<�f��;l���g���V�2���ą�Z)nVT�awS7���u.��Ө"琩���_�9�AIj��I����k�C�����O�!3�Ѻ�)��PT�_Mx���:�^��t�]T_Au:uVd�oT4L樵#C�V�Pg�֭��c��VI#$3l"̬��@��*H��݀�I�"e�"���*rr8ӂ��)-��U:�yd�R;L%��M^��F�G�G�\n����Z�I3R�Y�~r��k�<���F��3�����衪Faf�v1�8�sx<@�Ӽj;�j�";L=Q:����]����3��WB8]��箲gFA�3��YI3Bw�d�7����;7�S�v���UU>��^��m��0���kU��U9�c�x�,�M�L%ZQU��>�p��u���4��H�L<���^��EC��.�T�2�U�9��X����R�m��n=j��o9��AC��$s��_8`��N`�M���bVH�deN�x1g�}�A�U|&���wA~�L��"����,����W�~���-�0�*���z�߶�n�:Y=0��yTLJ��;����'/�9�p2/϶�梾��y��<$S}�Y�l�Q�R��E�z,�[�>��cʛ�dǻk��Ĥl<��P��}�Z�M�Bf��!קe^����Ĳq]�SoQ��0�&��\�r.�}���[n_���*kM�z�G�J��VWo��g�E�6rϥ�6� ��6�C�چA��wԭ��a
ȳ���.7�6����tH���xD4�d��V��㖕��u�X᫂��>�44����*�#j��Z:
A����Y&��LS��ܹ��-��3��O�{�a΂z��A�'x��PXc�������.澬09��4E?�`3_��k�P�J5��'3�N�MȾMJYY!1��F��;��#�ic��SZ<%�h9��Kp�ъ��]"1D&oZ
kqFP-+��汞�V���'��D�H���l��ĊI���-�d�
wN0��'TC�Wy�fDIl>�~l'�%��4_�LFq}���w�@T�
Uɑ�
q�Y��E��	�2�(5S�JH�;n0U�mkP�S�o�-a$�7n�`�u0��z���9Q��e �a�&w�Q�s};&0X���9h����{<�������h��u��+�G��[J�K�����?,����� WYf�oт�\u¹D�*��p)�W����ق�
���+l�]��J�Y�l�i߫v)"/�S�����(S��}D]X"K�s3i~�I֒驢�N"��3Ow�mS��&�6	���)(.�4�o��&��:���(B�j��Q���8)(�'�J�i�4B:_)M���ti��!��2�1R���d�+eK�R��i����A�l�9(�)Q����Ru�kp�N	�}p��à���Q*]̿���b��X(M%h��I�/rM��d�_ ��JS��P� i��ܧ���M�f���A�D�%���~U�ieb!P̆9@=��Z�H�$�L��R7H��j�&�K���ji�d�^Z$��Y�b�2)�k��ٵJ2t-�rWHc/��K� ��5�2)!q���-�LR�-�k!\i�T*9�[BA�,�I%�:�:�*�����	�<i�T X���Y&]*].� ~%\Up���$W�k�+ .MJ���J ��u	�-8�x1���J�*�B2wY��v-Q���F�/a��K�{O���9,��%�BE8��_������px-��Z�upm�.���l�"�W�y���_�t�>�p%���~���	��ʠ�5�M�&�J��_AO��Ng	�w�c$mL̐a��)%�!1e#Y��fg4Ʒ��������.7�-[#Ŗi�*I�:�� )�#I�t�#�6��#%m8���4v�������n��� N�b�����I��/�4�H��\)�l��k�%rH�E���Y�1,��K1��Z-ȚcHB�c�IC��m�8���ië>��4W/�4��4I�ŷi�~�h�/K
�a��b-Oύ���<m��Q�Tn/��$S"�QU:/W����Ĥ�Ĕ�D�)1͔�ݨ�Y{K�1�e/���F���/HL+H�6%�4%�7�9�Uw����b��3�˹��J��r%�9�����|����ܧ|E��#�z.��?�	�7���{�:������U�@|8��n~�!�I_��K���t�ϐE������Ĕ����F�<P�u�3�yqa�cJ4�����aݻ~���B���2����~��}��]��Rxz:o�<�%&�|age��l���X)�'���T���Q�����s�g��Y�BQ�h��n�������(�xL�n���
\�<]%�S�y���OB��n��N��i<}�*�0�����??P���\�f�[b=���Q���?�_�����Ỹ��O������:�_�����ء�`@v ��/q}F�W�����ҭQ��H���'FI�����fU�@�|����v��ƛ��k�g������~~��)�����ٶ7X������}���U�W8Qa>�Wi�<���@���eo������/���>��_R�5x=����׿�5~�a/��s����8L�p&�E�q���Z�6px3�ws� �;8|�Ã���.?����Z�8�a��9����a���8���m��a;��q�������8��C���a�ph�0��9�9\��jnⰉ�6��v�ః�W8<��G�r�=��kɡ��t��������<��aR�����>����#���'�������#�O�G���O���}�;xz_��O���͵�*�<��#S�3�=��s΄������������������������sI�,'n�n㰍û9l�p;�;8��a�9<��a�8p���	q9�0��$S84p��a6�39����a��氖C��8l�p�m��a;��9���.;8<��!s��a��^Op���&q�¡��4�9��a>�f�8��p5���8��a��8l��n�9��!p���sx(��ߎ��0)��l�8tq���q��a���-�6rXv~��Цiд�Ѡu��kvĴ��{(f�]��P�!�!;ɐ��=�aP[�!��]1�����bb�cwh�b�b�س���l]��q?�&V#�2�Q�j9n.���m��p�R_�	Ǒ���o���*�|}����翇�w����W�Պ�u��P�{��C2K���/pQ�AU������ύ
\з���T���A�XN/pA��^��W�ٚp�G�������w��o׆����+�]U��(��',�/_������+q�O��_sz�z�<U���A!�$�P��W�w���*�G��R���p| }N�U�����L���W�r}\��p)�C}(q�<���7��-*z�oQ���Y�;T���������;���]%�'���8��e��%N�}2����.�U�����O��qz����j�����Z�/��,.\%��R��^�����(���Z%�=}���we���\�_U�G��iO�1z���R8�'���^��.��	�W���ߦ��nީc��U���tB��������(_�S��S9}��~��^�����ǅ��T�[�X}�P�'���2�'[%�@��0��qz�����P��f3����u�J���O��IE?�|�p1�'pz��n{f����>[E��^� �$���������o��	���q�xI���A�������7��/Sɟ��_�#}�?:�ѷ��W��W��{y�N߫�oN�ĩ�y/���o��W��0�RN/pAߦ�%N�p!Ý�^�k����&�_N(>�^�#}��vN/pY�*�W��7T0�AN/��m���qNߠ������_��;T�f��߂��A^>>����:>�_�W%�0���xޟ��x�'q���\���x��8^�q3�Wq���9^��8���ws���r|-ǟ渋�/r|���x�i���ǻG��e,}�>�]��3R��P���_4$��|���ü|���[e�J������~������oWѷ��;l2��O[8�)�^�������8��}���$U�U_��~��M�������Wɯ���qz��~��^�+��ǡ���s����esw�>��q1?�+�����q��c���c8.�i:ǅ��qᯖ"���"��OWs\�'?��ŝ���S��+��{�����k����pῒ8.��h��u!ǅ�*��_�����m��_7r\���q\��v�����	r�~��b}���b��Kd�X�s\�6!����\�M<]�7���?����߼�q��-�W3|����������b��p\̿Z8.��q\�Ϗq\���Y�:x�s� �?��!�k��<|�x.��~�t���Ņ����?9.�sZ8.���9.����t���#����79.���mq�Y}�>C�6�8>v8/��r8.�'���
N���W�t1�������z����i���q�n��x;�c�a�v��s|Ǘq|Ƿ�����.������b�Y���ȡsȧ���_��U���9*|�
�R�sT��R�7��{T��*|�
M���O��#��t>O��T��U�*���
S�Q�'T�>9�³Tx�
�%���m*���
W�W���1%����g��r^�¯W�1\���?��*�*�K�/Fj؟��/Q��P�KU�:����kF�����	���$=�J߯����_W�S����V�K	�Ǫp�
���*�6�]�����R���97\�sT��s��5Y��P�_��+U�~��߽���*�jr�FJ��k���a>��9lఝ��8\�o����߂ܤa�x�o.�i� ɭ6?�������N���Ƃϋ�Ѱ}�_��+[��\O��4\���>����������'����)�vϖ�o��ί��g�up��k\���U~��i_�.��~*���6Ϻ7�u5\����u\[�^��^��?���&��+��I����\��?��\�j�ߜ�^ÞW=>�#\g�ٿ>R����fU�78]���I=�*�����Bv�ݝY�7Ee]}��r-Q�9%�"b�O��Kã�Q\Q0�|T+���'�y~�0��K�����8��9�Q��������h��F9��G��"�r�O�8vbُ�� z�#Dx$�*�{�n�f9��c�"S�)��L��~#r�{��{#2��V"��8��H]+�k�sa��\\E?ф���V~�,?ȕ��U��V����X�#&�����ݰ�j�zmU�V�{��"xQX�+�(x�s���8�ӭ���^�б�?�h/>��Zf��3�1�?�;���偊� ������m���sz~:��0P�@د;v�U�$Tr��� ��2ӖB��38�d�Zm���^�j�#Y;�H��I�鴾,������p���a�P�>O`D7S嬶[�N����aq�*[=�!����Т�Ҡ7�G�CL��{֣���m�r��f�ϋma�����L)�P*⿢6LB��q��ϓ�������q��:^>��*�h�8IK�8]a��X�K%*�޳���}^�&^嬇���t
��f�9H��9=4"�#���"��9^^��s��g�)���D�$~F�Ds:�@w�,�d�V�g��eg41�I��x��{�1�h(�N�:C�Q0�mFq$ה�ǎ���'�����I��P�@u�3t�VdF�![�Ԉ������Ι���_�\�T��Q����q�!܋��j|`\��V���b�뇧����tJ�L��2�/����"�����<I=�	��C�iu�~�@d����N2b��s�϶�_�3�3Z�D������ϖ�/A���3}�,�\�G]�G]��+r1u�m2e6(|q����_X�G�s����Z�F��+�E������۽���2�[c�ׯ��*"�VK�(��
u��㊯��ˉ}�a��I�����1��d����o}���\���O1&ڑ����m���5UW/�GelH=���'Jv��F�p)�W�#��#K��"&���(	���K�xtoAYB��K}�2���FD��i��h�2z�m�}9E�o
16�>����x�� e���g��"Y��b�ĎofL����CX��W�%��?)�O]�s��{�"J`x��C�2�Ύ�W(1��Cq�ms�1)W�g�c�6��yWX��oe$T9<�|��d����P�|�0F��9�U���ؑ�<F�(RQ�]�C-�@����UyYI�¶E�Xh~I.S�d$��Q�ׯ0I������2���㠚Z�4�K^�Y~�l���0���qF�VvJ|	`j���ƶj�g3�_�Mu�P506H8/��'�T�i]�<;$��.b���H�*����n��Y��p��-��;i X8aeR�%S�f�fR¦"R�dM��\��=��"�9.)�0�zIA֬��dq�����5TIh�4��p�_}�E�4��^��^�+F0�;+�VY�[n�|��܎���̀q�b�t�8=۫��h�SDѲ�z���p �X�*��Ȇ�VO�t�%�9H��PK
    \O�HD��mW  �  /  org/jnativehook/lib/linux/arm/libJNativeHook.so  �      mW      �}{`SE�����ѐ\S�Z��EKI�@A��~X�ЊU�4��Vڦۤ<Vv� �.�
�Z�V�7jEDD�*������"����h�sg�܄������00=sf朙9sf�����?��GK���?#�d���c,��یdf�a*3#�;;�ER����L&i�!'in���=�7x��ĝ�k�2ܤP����Q�n2����@KN�l���e_<z_K��-�.��.&Yz^��6.�ȯ��2� �Ru�����.�T��U��,,/�Ɲ$�K�H`�|���OBw�����b���.��F�e��O��+�]����%�]%«��0O�7��2��$�.n�.���S�Ctqg��W���:�O�Q�81N���rO��~S,�K��1i������4
X¸������:Ay���p�[3ux����.���.\W�G�b#�.����%���&�ep����"������/��p�����g��)��;�g����'��_��Y'�c���ia�uӥ�>=�r���($p�I�Nv�N(�g]�������=t�
������y��a�ؑ@�66��o,&� ����`����߀�.�@t��ӿ�o}�&�g�Hy�6B��8��Q��Ɩ���� �%�_|&���#�~��H�C_N�"�7�����!9�<_#>g4�)�������.쩘�^��cr�(��,��ʍ��6��'$m�J=U-}C?/�<���s��1�<�m��m3���b����ى�t��?CcLy[cʛ�cWF��� �o&��~����obL~�-N�c%�?��1�n��1��ك��������˘xe!��c��v�
w6�ڣ?<���n��y?�7�B_���������;c�!�L]�v�Y��rQ�ρ�����ώQܶ���1�΍�o�0�0��O��5��F�{�7c��)��1��Z��/C�\]yL1��Ӿ��O�"���b�Ey7��;"�_�ɯ>f�C��h
�WD�]L�Kc�o���4���>}c���>$\��T���)���`�u�tiLyƛ�:"<�x#њ>^��h�L���1�?��0>	z{L�{�X��<1�m��ϛ�rH�=�v�����~+�o���x�S^����YW�g=�~sOn�h�3�}�ro����+;/2�W B���?§��'��uf�~��~�U<�p��̨�W{Aom��a��� �L`�qE<e�Zߌ�@�W[4aD���W�V��q�c<�s���[Y�{��gy&�t#*���/�*+�WT�j�U��?ۭ�;P��0�(�>�gV�����:8�SZ>�]����+*=��3*�gx�}���
�w�/���S����>����\W�V����3=<��q��ENԼc�5��W��w�f\uM]p�,_u�3}s����e"奾���U��>�h�O1��>_%O�	���\6�:_�>�p.�JKQy�v��uD�����jk���7���vD����[孬����,_m��?���K�$Z9GVj���rj�YU�<�`�[Z����Ds��,�[�;��:~�8�e՗WW��eL�P����,<5�(SGp��<PcW�����k���ʙ�+�.�u�u~�װ��4o�Lμ���_V㫦�Uz���@=�D3P7V�O��@`�xR��v.���[#�?��(Fh`nU���_�cœ}���2-�_m��X\8���QM�M$F������y}s���Q�T������� BX1�w��
���ڏ�o�/������!�L^^O�O��*�C��j�6<���+��i�VT$�N�i���#OU]e��SZYQ:�C��=j�괖:���WYCb�9M�TeJ;��<s�_�R�Y1�aA�D/b��.�
������h�U�(��Zo�\/+Fɭ8(�a55(��	�r��P+MU��8�q���|޲ +��C���3+�������Xa����QZ�*�HG�D�4��!=��E(Fڊ��t�`O�d0=�5\Aщ��vVEp�F(�r��W��[Z���OE�Q�@����$�6GM�JG	��?��a�=����_M� ⧯���4.0����� �o�	 ��k�� �tV��kf��О��3#cxG��`�_-�4'���+*����#�&���"�cVLCW$>T�5aEGc�+��{1���MkZ}�8�3>9�����"�"��j3�/��U�!j6��V�+����L�q�����a��2�/  �?n�O��A�a���f2�S���|��Ǣ(�#���܌Q9���q��q�Ɩ ���Q�0'{Pؚ�;���A9�e�aIn`[���i/񈀫�A��<�xC-cG	b�=����';���X��� lթU�Jf�~%8k6�0�+	f���E�	��f%8�;�K�O�Ea�/&X���X8,'���J����J�wX_4J�ؽN���#H�0��A�	��	�$N'�k�0�Bb.�
֎O�O0�3���#���H��X�0��	��<�!x.�C0�!�
��ڿ�`:�C0�!�5B�^��Lȇ`oȇ���� �Y��>����A�C��Ck���I��� ��~�X�%x!�a�b=G�b�S	^��	�a�5��'���m'�������&8��]�1��`>c��u7���C�}�v;H��G�r�)A�y����A�|F{�q�6�ƺ� ��v�ע�	NC�,E��¿Aڟ�t�?�
�?������r��)���O��O0��'D������|Z(���[���}Brs}Hi^�l=�Lh�J������ʒֵG6���5:�j��οD�_������:��_��O���t�|���?T�����t�t���Ο���u~Y�?�U�D�?�����?��w��;t�m:�f��οV�_����W��Kt�E:�<�?��W��e:�T��H����G��Cu��?K�O��{��I:�]�u�c_�����������t�:�6��ο^�_����W��+u�%:�"�����+u�2���_�����#u����O7��ZP�W2,k��5�ت�a�� &���CƼ�{1چ0����b݅p�jhc�E!��6�,���%VC{���c��J�ږ��>@��at��k,hhalah/�a��ޤև���!�����KC����l��V<%�fE�Z{IC����"ͭ:��14��& ���}[V�L~j?P�r1gC[�ki+�Mv���U�+�-
���O�Υ!;�ѵ��Z�d�w�{�\���B�pfc���3v�n����o\%��߄K�$�E<�
�xr۹�}����K�I�|r�&��4����]%�fVئ�x8hnL�2��G�ƣ�x���^����ɂxIΒ�,����B|�<oA�s����ǯ�V�}��h��XЏ�������|7i<`E�2	g�{�@��In�%��M���5D�K>�
�c��	?9*3�Eef��P��3�5:$�n�۲�%�L_����m�Q�o��Tb������i��̋��7��K���6;[���Zby-T&3t5��P֡�x� =�N?��s�e&B��nu��L)?
7;y���B�Z�eVW����n�s�
�ي}V��jx:�K�y\+kB_+A��k۔�˖�������쇩���4�����ꊐ3N��8�N��1�I�8�����B�V�Mu��ׅYℙua���/-ܲ�V��f�A:l�b����|jA{&��9�;B2�~+����r�{��й�js��������xKV�e��5K��d'��&i��\�C��2��C��SYA����h�-����}��ϧEG���o����u�ɿ��v=��?��o:��_@�{}���S�_����O!��j0��.��"�`9\	�|� �T��-ϑ��~5�ϧ��غs\��eM�1��k�zNzɚW�V�[�)X�����\�/-o�/���6[��k��'9(��gr��Qv��?����m�Gc��JZY���=V׿Vi�[:4���d�Q�5����5׵�t�O�D�+sf�b���������N�TІ�j�r���t�w��?�u�$:�A����k�Xt6ϳ#�K�=�J
Z�2P����_��Ay�W����0����%�l��"�C��a<ק[ޟ�����1~�Xw;dwd����m0�k��_B�1^�OtEc�-С?���1O-Q��<¼�Ԥc��y��Cy(�MȄ��Gkoeu��Qr�)h�+�����
���?^�*P�$�˂z�L}M_/��^61vG�u3��D����C�{G���X�#kn�d�u���$������:5\�-|Iw�xW�F���@Q7�H��dE(s��mN笨9����E5+4�o�"d3H�=�)x
��,�\�sB�%�2M2]����%[2%�����W�N��(������:c�Yr�,���$ׇJ2���J<�^.䛓_��%^��̈윹��{lF}�X/!��1r2�iw�����&d;X���+�g���+�|7K�{2�{�;gP|�:;�o䫗�A]�W�|��7՛BN���0�$��������=�y{���_�����3R���{����ƞ�z�!��h=]�W����C�&'MX��4E����	�=j���^�h�o~h?�ԓli]{����J������%���3o�ƅZ;P{$���!��K�vRy�4�^j̈n�֟�K�h�E��o�L�.��v)�]�}����NƏyff�\�֌_6���x�2ߞ���@Mz�>�\�j��@eR}�2=Z��D��B�yI���D���#�U��S���к��������W��t���E�ir'u֟nq��V�gyZľ(��N��4#��<䏌� =Pw{��m�]����m��ή��������I��E��t���E��S�.o�<=�_��S9���I���Ʀ�|�ʌ�&����4��.<AK}��{�1wx?+ܿ�`����J��?�~E}*ܟ�c�??%Z���x��%�oЍ�f�u���ֺ��m�76r�b�z��ps�h�b<.S�
����������-�˄�����
n�e|}�6�����:�����U�]w1ܨ�|�g�opuH70��j�ap��'����3�%��{  �.��mpG.�k*�8�f�>wΥ|��ϱ�����4����-��`��x���k�� w&������q|�v�h���g
�Ta`/������;�s�?�`
�!���>d��O2Oۣ*h9���v�kD+�h<�D{o�#���rwh��Y��aK��.�֢��b���֦���F]��Qi�c 2�����^T����?����jo��	��a;ٹ���{Zk%�"�=U���2���(�#Zmlr�����$�c�~�o�T�^�f�����k��0F���yf��2`����9�ΛC���~|�����M��xb��Z2��-��W7w�%��:4L�[c���P��Ү�,���h_���o�ع�d[K&�C�	��\x�䵖��]X�/m �}���N���� ���C k�n�����*]>�|�D>SA>Y�����'���t�x���
��v@�6�9i/��]-ɀIM��F���7�� ���N^ƣ��ߋ2R��D��d^��3�+�t��E���<�1�g�'���Z<i�}}��_�gx}�榡4&ie���<�!��iV��ZSx:��n����m���3�N�e���l*��u�z|#�qT�c���&Q�̀= Tu�
�x��c�:Jy�>z���-��N�s�v�}��@�y�w���c^)���}��vƼ��%�9������=��i4���p�3P��m��422��뢼V㯉��SɻIay7a̽���UJ^���2sY�ܬ�T�+��
z#�L������6��=�U�|��J��?�W�?Q>ݴs����G�y�ՀVϑnl^}Hv��F�s�<���Χq?ޘ�rt��+��`.�ܝ��к��霎�AV"��*珶o�o��YM	ͣ�4�a(X���aꪎ���́G�XI�/�c8���B��07&n6�Hf�N~&���gU(I��}���n	\:&*�8�kt��bdjs#{�άZ͕b�淄�v!�И>�:!���"������b���P��e͑3�?����v��+���.!?+YrQY]���JgQ�f�V��Vh��G�//��'s��t����Z��h���N�����J�΄$�+���o������ ���dN擜[���$!<���tq�[F��\qn���5�5�[[(W��V�!�dQ��Y���²j��.�X��ƛ�����5���2�V8;��~�W�kZ�����](g�-�nm�hv��Т3�C��K���6���c�5�j�Du�
�~f�6��'qf\4�>Tt�8��=qз�=��@Oe�Q��(��1��8^��v�zF4���@��ޖ(�U�e%x����x�ZyxM���է@?�DY�DY��+9��_O�����W��P����sO�>��EY${7������D�A�f��"�uih3�Ӊ0�X8�a��nA���7FfԇF��Ǆ���p?|}�(� �hs��q���{~j?p6ycRt������z�ω��}�z��s@�C�)��z:��5�>�uq��wv����S�ŕ�'����OO���o���$���S�'��>������H�u�x��fjw�e���4���H�h<�����}���t}�q���}(�Q�a�׬
�����D'��`~���¶�]�5��/v}x�`�WA��`Nv�Jen�J�%hX}<����V>�E;s�Uۓ��W�.?;[�����O���4�o{��_C4�6�ΰ�9+��k��o�lXAC7ȷ�ڵ^�%2�8�q�0� sY�H��y=d;��':��_�������sAC6ض��¶N����kS��D}�H��t+��e�s>��y�sG����[�����/��8����T��s>�9��׺;��}V�����;��)҄�i��ک�l��F
���mCw�j.a�a��aT-|�.�W ���i��Z`cOlt��-�=�� ?	���,� �x����=���Fؑs�r��F�7.�(��0���*���
h/����Vb�"��  =g��� �F�/#|��$�a�����/��@�z6�d��w�M��ݟ��F�tש	����������[
����q9��ݹXo�%Fw�T5|�����/Zx:�L�`L]h"�rs��q.�rY�O��-�nG[��$ے��쯭K�r�m���#}�-t���\߅h�N�L���M��.ih9��Z��]F���0��ZKؖ;ʶ��K���mFZ�h�"�ϋ�΀4��9��1��0��h��ߒ�n���+d`W���~U�.m�G�ևt��A���|�WY��7���0�O���1�HtNt�Ρ��-�o��g��8�F�c�,�0Q7�.��O�>�v���.��?��8��Lh�����U��܏t���!K���z�EnD]���ѽ�e	�7.�iQh��'mk�p�6���s*0����>��ϭ=@�����/S�Z��b�l�{W���h�7k�.H�\,X{F8���_Ge4���ɘ;(o;�rD��r�ӼB6=���҃l��T�f��#�5�m#�mjx��x���MA��n�<}��ڦ��(#��Tm�P�k����)��m�+�p�d	<�6�k?��[���H�Hנ�m���������&mmiT�jY?lkK]A�'���z��&i�a��L.sj#��an+��7���?S�䷷c�}E�s$׮P��t�]du���ۤ���R��l�[��E[�|���r�z�p�Z��Ϩ/��/�t������5��l@�Q��&ߍ�4ӏн�C��w��Sw"�;h�i�D���#�h$mϟ�1�@�5(r��H6A�����-�I(C���˽�5[��������z6{���'$�����-�⬀Gw����g�ټ7�J1?�^���{=�>�{�>6�e��pg��.��F�Ӱ�3�������Ovy:p�r�7�x��*�Y��!��m=����~7���M��~7̽�>dk@�\�$�$������=���q&�ګ[��+��=����Er-���J"���1�v=�/���"v=������7c����-;D몳`ah��|�L:`:Ш�ݲ�t��/h:�A����-��&����׉�B'(�&�Nl�щ&��Lyb-E:�>�m�.c�>0�4����/�u����֟����v��A�y���D��n�����]?��k"m�/���H���Xi����5���	��F�=`Y�I�ili�Q�m_l�b��Fbm��w/hsX�H��6����/�����(���W�E߼w=hvt��R�똬��w������S4��m@��#���m���b��
�%I}[�/��!]3���L:�'�]:d�/ɀ�0�зt��]~�+/Ջ��O�v��o�0����<�q8�C|�E���e6�w?�p���6������S{o����\�u��:Kr/�f�{-��<6��6�Kis��+�W���V�lB~.����PC}H�uز�ɘk�;5]k����H�R7�C��MjIr6�l��F��h��>��ɝ�$�΅������5n�+�N�;�X����������w��nqbd\8*�j��E�4�mʱ^�v�6*Mx~\�c��"�%
]�M���n������I����f�
��n
��q�%|
��Bu�g�#a/�N<T-�s0P犳̩p�k���}~��w��ze���¦f �C�P�	��s�I�!l�L�����ȁ}�b,�z���ф<��
w t�}�����5͐��>X�sc=4�����g�|���IL��n9\&�ٌ��9x�0���;�%�8\|�#�
�C�\���UZ��g螩	vZ9�*Vu}(<�O�=�R�[��z��E�ހ+�߻�m�Hoԭ%����te��_��yr8��ot���y��f�g|��Z`sм��%_�f���h��y���Fg5����9o#M��P�[<�Cwyj
Z��ٺvg���%�k����x"=K��O�[��u�ߗ�h���M[�Cw�"c�N��$�\���ԗ|Ob��ބ2�e�[Md׮ե�"�#"-�-+�
������0_�k�<�.���a��/��˝�#��?}�H�Y���6��7��k�L�ך�lٷr*o�$����3v
4�WbE���z l*t3���G��0/�����gZ`�%5���Fs�+$7�+4_"�pg�I5��A�Ns�h�nF�ԝ{oPoh�!k�%Н���28%MV6�����֚U!{�_��M�`�;U{����.ƿ�X������%lq�sghƽG�5`������M{�9:������*�%�>���?h����U_>�U���ş����g�K:�"zJ�)ҥ�K'�tc�����n��pCI�$��S8o9�l���_ؼΰS+g�~��Vԥ�����wx$���p��V�)��Z���
b}��]���������a۷�VI���7��T�g[�M˚ox}Ik��д�Un^��zsC�2	k�%�O�n�9Or�����7���K�A�\�>� D�6К�����:h�H!]���Fg��8�4�vH>��O��Ju�Uz���X򛸾ߐ}t�V3�΅��9ѯZnh^��ʉ��kA?#��i����G-N�\S[�J�|[�U�����Øql�3���<�뢶$��۲�0�v�=���9�m��&�.�߅��F��[��=4���~�b�OB��x����@ې��Fg�KC+S"��31��<�y~F�.,���Ҳ��o�Oϩ)�{vO�e��CcgW�j��%���j���]�#�%�BeI�)�AW;�w��#HOwh�1�_�ȯ�	�H~i"��\<�]�H~;���)�5��/��]㌖ݭj粫�$#�{��`ZlG'�B�ӡ��n(���vr�%����b̧p�v�oҽ3����[whcw!�S�Õ�y��#|�E������\��	������C�#���hv'=���52���ҹE��"'ߗ���u�Q����?�Mu������)��JMn#urۢ��g��wF�ے�����#ϗ.�z�f욡����_/��z��I���q�:<��ZD=�t�,B���z����i]=���������nţ����������D]�?���E�f��z����g�)�E��m�\��Ө[�H��:3,\����F�ٯ��ͨ'�7��מּR�IQW�i}�>н��.�3���.�<]Y7���e-�eN�m7���ӶNQ���H}?D�=��0�V>࿨sML��'�s�>�:wAy��X�s�m]w�i�p�s&G��)���=��́+��"��aK�Y��b����sLMX3����U�7D�0J���	!\��*����V�)�l�W����s�z��3�3W3�C�(_�Jkb��-���8͝�5��z,� >6�/7�fM�y�=���2x7���!:����Q;���b��`��t��ƚ�-J&��o�ܲ�ir�}~W�����#BkF n�F nD��~.lOa'�O��n�0Ƥ��nZ,	ԇ����q��w������N��`	�g��������NK�@ZSt��/_	�ۚ@w�W�i�����`�Px�����ʦ�}���=s!W �|<��1�ɽb�T���ȺҞ���s�0�3��v|�͌N�[6�����X�{rbC��7[��%�����V��A�z��z�V�2��稗*�/u�~�S��եۅt�t�(K���2t���A����2���Y���\.�?�r�m:�@�R)-=�
������ �(d@�F�h/��e:�Pa�¨Ʉ��	�٬���~.�:���?���c��͌5�,�]$�)/�Q�Q�tqϊ8
�w�
��i}�;���h��,h|mf���N4H��F��ZFw���xOi��P�H��1�djw��~�?՛5�s;+�4�A{���"��cC���� ��A]�{$�v������P<�>q���'��j��O*�(7��u5�l�<Z��p���<��}\�Uy����ϣ���mXZ-d�8T<����6�6\�ż��Š�{��y��N�����:,���\�|w�Y��W�]Dvc	����g&|Y��ka��,m]'������B�?��:���s�]��p�H�m{�M˟����~N��~ZwoF�mv��`.k~X��z��A��y��ȗ?k?p�x�`1���~p� �I_��'���XGGu�h�����#L�#���� ����S����"�S�s�:i���� v�׀�����>�]����~L��U�C{�E�f7ڎ�ih�&c�m�݋t�gq�s���п+��V�}��*�ć�j<O���_��1�˯�W�W�+�{�Fz��xI{�I��"�����zr	tsC+�ogyxO��M^�p�^���ϴ�;�&���zS(��F��見�chn![���聱���{��J�{i�����ɺ���>���-N����[�F���}ws���2��Hv�o^~�^���M��|�V�s��co���Q�w� �]+�t�/�Pz�H;��<�)-��ZΠ�7�s@SZ�żv�2�m"���i��i����~�Umv�xv�dFy�;���]�c��N�%��*���Mi��9.�?��=s\r��m��:7Cn
��Kx8�!���	?�3�4ɺgw(]8M��5MϜ�į��N�׋�p6 F�r��zQ�),�9c��ܯ�������?�v.���@���՝������|(�#�D.S��Q,�l(]X~$��'����Ʋ��hB��wH��D/:H��-ރ��s�1��|=3~������%�y�7a ee�u3�v�A�_��mCf���S:��� �s�z!�e�T�,��,5�
w��]}��{)��������2���h��u��p v�ȗ�F��{E�V0�_��Gk�\y9T��t���E�#i��W�H�"����a������i�?9�]�2��9F <��ҳ$"�z]��_����Ng���n+z�N���KA~�8S��>��.x�]�|]zf"/F�)�œh�����,
.���J�f���m�V��������ch��ftb�bN�)h��pͨ�@'�Tf���8ؔ�ݓ����hW;ݵw�4fR:�S���}ZE���"ޡ�|F�wh�X��5���l(ޡE��.>��߯C�=�����ޥUֳ>�_�1Z_��˪ي<.����{��t��P����2�1�>t���K�3����N,3K��v�~�2[4�Gf��I'�������	�dV����L�Շ�2;�޹�F��9��2�t Zf�N]f9�;2�A��'�YP�9�n��efF���dv��>t��ٞ��evt����O,�����v�2��Z�7d�uZz��$��:�_fO����l״��mBfdv&��@����2Scd����l��Gf2���	d�(������2�Dݟ��l��>�������ev-hnu�XfoYe'�Q�'3��ߐ�ɼ|��.�#��j|���z%�}��%v��m��o��/��5�;$�3�>	�_Hq�����t6�`ೀ�,���/����M�V^����42���w�7xg�R��C��Ɩ���m�\�tF�Wè�}�pR�����f����I�5ھW#dV2������n`�-�Cx��������?��Sk[oPopҾ���2�-N+D�44/�d�*	��E�_�p��_��!\�%��E�P����."�B�����p��_� �#\�%�XEx._��E�B��K�/0���~	�&> ��/��@�9~	�F���/��� ��!\�%�H"܍p��_�D���/�Ow4�b��ᰡ-C��5H�o$<�x�:����74�������q��_<I{��6|]{�3lΛ�k�a�ڝ��sa?�Úb��}��Bz�k����kgd�>��}ͧ/}ͧ��a����h]uY�<����25�W+�;>��_�?�x�J��D��	5��ˮoԧ��;>���O�0=����x��'2�#���҅���zY]��|U�ڹ��D�Jj�jrfj��*�������P����,s\~$��`mE���dEd����v����B1�r����c�/8n$��=�|�e�+|���X�?�7��P��2n��	�#�34���I%S�EF#��}+��q����	���%�Ӿ	3J$���\yr���O��YC%���ê�,9�}�	�F8�_���8�vU�?X1}.����@Ǉ��F�_�`�6=>���>��M<"-��=�W|{����*$|�s�Cw!�^Q�K3�i�B���:����XF@�:��!��Y�ʊ���k߫Q��m����V�ۦ�)�����P0~�8U���to�O߉|����B���=�7�t���(��3Xj����L��̶E�v�V�U�Wa�Բ�oe�����=4���I,EN��#����:�Ch,�����D�Q�(B��u���5�"��O��V'u��9�'��H�V�Z_��E��<����'R+�h�T�.�ǊJ*ITj}���gp棲:�_��Ψ�`m]i0���_��Cͳ�@\o������F���j�o�VN�T|��ʐ�V��e�^��2V���'�5����p�9.�)-��4^t��H\��ΦaNc�f�e��4�ADj�[@�����(]�������ص�+��������7��pE�O_J���"i�{ǥ���)�ﰝ��W(�AEu��syu�����������gv�i4�!��}������7������w艀�MO��t0���Ӵo'I,�XWfdݘL_ve�33;�Yؙ�ʒA}}�g�������>�*�S@�
�4P��:�=A�ԙ����A}��@��٠�j�ݠ������ P� P�z0����BP�E��ԗ�:��@=�#@=ԣ@=�c@=��@=ԗ�:�@=ԗ�� ԓ@=ԅ�.�堞�+@]�+A}��55VY����u	��׷ٳ����&�+X�+�X)����l.���7k_`d/��K�e;���)�hOC�o��f��)�إ��.CX�$��p�"��\Ʋ�j.e�:�E��F����X�i�k��36n���f��k���p��յs��f=����?�>q���T��O��~/��n��]'�L�����u5�T�k�J��n:�H�J������F����e����pup��f�����	��p��w��;�l-'�q�I���ML��͖�-��+���n�[
����H�����;�?�#s4����/�E_�z�Y�GOEQ�7@<!E?}���ۑߟ0t�A8���ן4E�?�U����j��H��9�j�p�� ��R�. %�xFc�̓�Տ���d�.i��ni�t�t�t�t��T"=(]+=$�Ik���#��G���$��N���qi��t��A�ZzRz���6I�i�'m�~/m�>4<#�QzV�'5IE�V� � �^���v�.�"%K;����"픜қ��-i��T 햊���j�?R���4Mj�.��$���H�Hi���KgI���/�ӤCR�tX)})����&IG�+��$���;�'�Tj��3�i�)�kH�0����Jk9�c�^�C����-=m8O�l �`�I/��;�ZTJ�J!C�C���!E:j8G��P%�d�F�˘+�m�"�c̔�5^(=h�*=dL���K����0��6�J��ݤ��i�f�i�q����R��Ȥ��������7��������Ɓ�{�Z�Cc����:��(I{�}���3�/�H����/��������Gc���q��G�b�N��K����5��G��u����>�N���ݮ�{\����p���\�!�#�^ף�VW�|���|�k�����|�k�|��	�A��!ד�î�򣮧��\���]O�O�6�O���O����v=+oq5�Ϻ���s=/osm�_tm���^�_q�(��zI���.��zY~������U�-���k�n���\o��v��ޔ�]o�-���V�.y���׻�>׿�O]��������僮�ȟ�>��p}(��H���cy�k��n~�t��Y�y��L)��M�武4�6S��S��ESO�K�^��L�˦��WL�_5]`�a�2�f�c~ݔm~��׼��2�ir��2�3�m�o�e�1�c`~�4��o� �nS��=�`���!�fS���4��jnn3�0�1�4�L�̟�F���Ƙ��ƚ?5�3�7�70]j>h�7f�`��4����2�!S���i��K�d����]�B�n�$y��H��|�|�y�|��
�~s����J�A�U�C����#�k�G���|F�cf���l�7K�z�,?a6��f�I�E�h��O��Mf�������l��1+����&�D�9�K~�얷�G���9�����K���v�(�es���y���y���|���y����"����N�%�����y���a�.�p���]�@���~�ns����R�}� �?���	��q�G�1����r�9[n1;�Vs��f�)�1'�!���'�ty����Ϝ!jN���ϒ����g˟�{ȟ�ϑ�0�+2�'6���4��W���9U�ڜ&c>C���U>jΒ�3_ o>S���)3��4��2������wZ�l�˲�x���5���<h�ϲ�x���,�,3>b���Q���c���u����[1��<j|��q�e��I��F�kƧ,�7Y�O[^7>g�����&�V�
�6�J��U�-7_��b�n�����6�+�ۍ�Z�i�aYm|�r��u˿�oX�;-�7-w߲�m�eYc|�r��]˽�[�3��o|����ղ��fyܸǲ��<a�Ĳ����q�e��S�S���M����-���Y�?�<c�����x���K�V�W��G,ی_[^0~cy����%�Q�v�w���wZ�L��jϸ��2�Xմ{�)i�Z�Y�L��zw��5iZ�M{��ϴ��;���+�kCڣ����k�6[�R�XKR���R��^��d�I}�zN���sS_�ZR�[���l���uW��ַRްzSߵvO}�zC��S?��N��z~�G�^�[3S��R���$�`]�r�zcʏ֛R~��HiNx1�%ᦌք���{��Gz(���/!=�ӄ.���3$83&�3>KH��<ah�	��%<�v8�e|��9�-iGzd|����MBNƷ	YGwڌ�]6�z�MV��L�=6�z�ͪ�gKP���lIꃶn�#��ꣶ��V��(e����mSR�ۮHy�V���veʓ��R6�L)Oۺ��m�Ӟ�����vu�6�Ԕlפ�h�6�e[j�+�n=w؞�x��d��W3ް=��Ӗ��i;K}��C}�v���vnʻ�~�m���l����mm����m2>����푌f�'-��2Zmg����cے��{~bKU����g[��ms�~[��l��<h+���mz��m���lj��6U�Җ�~e�����^_��=��U���6��Q[^��lJ��m���`;3�-W���]��v�zw����.���d�>ХWjS�G��]�I�ڥw�.���x�+]�SwtY��z�5�oty5��.ִw����������ܐ�A��R�u�;�c��j�}�������������i�}�)d���]�^��M��M���3�o:`�����g�M��?2}a��t��l:lo1}io5}eo3��1}m���b�־�tԾ����S�����;�r�à��0*k�r�ä��0+�9,����#Ay�aSrtQ�:�����CQu��4:��c�De���򸣛�ޑ�<�8]��8Cy�q��ё�<�8K���<�8[���lq��<�8Wy�q���P��)��Te�#M��HW^pd(/:z*/9z)���ˎ��+��W(;Y�k�>��l�G_e�å��p+o9�)o;�+�9�;�ʻ��ʿ��ݎ\�=�`�}��c�%J�#OiqSZÕ6�e�c�r�R>q�V�:�(�c�O�����ǥ�AG��c�r�Q�vLR�tLV�r*GE�׎˕oS�oW(G��w�+�;��.���n��{���G�W�O�_�u?�v?�q?�\�^�u?�\�~D����r��Q�s?�s�S��WF��+#�O(�����'�1��X�S�8�&e��i�R�f%߽E��~F��~V��ݤ��S&��W&��*��mJ���r����K���J��e�J�+�U�W���;���הkܯ+׺�P<�J��M��~K��~[)u�R�O|Gy �]���+%�V�&��<����H��G?P?TK�HY����xb��>�Ey"�Uِئ<��G٘R�J�Dٔ�Wy:q��9�SeK�~��ʳ����ϔ�?W�O�B�rR~�>��q����+e��������g�7�R���?�G���)��W�KlWP�t[�n�6Y�ҭPz��i��V�W{*+��zk�zh׏J��=Uu��
��]顝�H�8��|Ձ�`Ŭ����#����J_�v2�	�����ʲ���򬩬��PB:���s	O���;7~8�"�j����v�����w�����{靄��}�L{���4=c2}���8� (6E�)N�OkƎ���Y3m�GΏb��'��l�|Q�,�I�:�7��_�S�A��+#�K�̨�t�Ye�Y6g:*�;У���Y�]�AY��i�Yj��7�N���uZ����F�̜6F;�NPu�;�����#����6#`cqO3X��lv�����A��*��y|�Ac5��o_��N�l�|V�2r*ttj�o�	�^��z�5�\R��G���.xU䊊�2�� ;.��'J/���4��_y\����Ac'k
;��'���T�,�ͨ���J��xi�ǟL!��q���I�(�#���&����==�Dv��q6�;������莿=��Z��'����.qvMW�LG�-���Z�$��H1�d�G�l�hsҴ�,^R�H���������4��ѣ"rDی��%:^��ęNX�G�����ٰj�N�x�0�G:T�v�X��#� ��C�2�����o�s���3U %ե�P�p�Z:�<a��RFJ!ΙO���7�"@gˤ�P�Ju6�pZ�0�j㉦��@ �tx�����|"P�5E���$�u�(��F��jK}�qN������vɥ6;����^����O�鴴���*+��UH|�ڱ�ʹ�ą������B�t���W���V���Z�3'(��G�3rg%?�Rk,~�b���-�IL��_�P�3T#��:����^Î��W�`�_�~����z�����I��רHT��>֠��E�8������Ǘ<�G����|U������o��~��~���������o��~��~����ۘ�aAJ$��S�N�?x��w0~�4�l~��r6cg|DbҎa���C�t<s����Dg�wR?��{�N8��9k��#�9���w&\S2��3���&�����o<��g��2|�ƾ4��<*uxG��������1���H�$�d3b�5s��:���9ك���5�lW�ZS�����ݯ7f��"���V��xM�3��*%H6CW9I:]:Ә,�%u7�m�!�J,;0�*���<�+��Yv��j$�0X˲gT�e�����j}���{j*�,�8cٴ�β�A�����l_�gz�����x���޹<M�]i������Y����NXv�����d��M���k+��}��2="��q��>�q���r\뙌��eR��8�e�8gD}���ƭف'h�~^�����]4������yAi�8��|�?M��:p''|4�'r�1�w� �ǻ��<��Fvz~�t���\�r�><"&� �|r8��
�������������cc�E�o+��_|yt��ˣ����S���N��/��w^�|Et���p���c𣏄�z���,&�D�)GzEK�<&�[����ؕ��MWE��*:�����w^�rjt�Ʃ�񋮉�_{Mt��k��W_����_V��4:�hY4�8?����Sϑ�ӓ3���s/�4��E�e��s(o-����#pw����J>�N�AmZ�m������32��g
��Y��-p��1��W��׬��;�l�����*��7��6��o[)ߕ�w��6
�$������MÛ��I�^�I%�u�NS�����S�g�I:�F݀A���R�6��b���:?���������Ӣ����Y=�����o�������_t|s����s��s�����=8:>kHt�kHt<�0:�~at|��J��KX��?i_�A�2o�x�߮��4p�l`�ȯ9�<{tx������bҳ����52:~Ǩ�xutt|�����1��1�%�"�@�����Y2��(��?]�E��y�V'�xƼH"~�t����q��\D�n�r�;u��yK�? Ϯ'"�g=��OD�[��!�Q_����ϟ(&^.��o�.:�:3:�fft������������`��kD���[nc���?>����L�kb�+uCD�G�˧G]$?L�t~���~���3O?uv$��G��w|�>*��3����p�M>t6�I��9?��k�||[$q�c�>�P�eF޾��y}T����k��?�?�����_kE�c��#��(}c$�Y�ȋ�w���I�a{/ܞ�k#+o�yu��ML��:���#:����1���ie����ȏ���������y�x���F���I"k�-�H�S|�O�YǏt8'���4�]��U�Yr���4�P<��	DocKc�= �����㟎�5o���t���7��q����\ ���<��ؤ/o76���,���׷3��F���1��Z����E�wcʳ�����ѿ��?�9������E�s4�!1����DN}5������f�ޘ#��������mF�zL�Gfno��Kt��1xz>����0������z�`�4��� ����ј��,����߰p�c��ߏI����/��3���|���<���/��*�l�u��O+�_9ލ�C�.o���4Y��.�u�����܂~��K������~�&��(?5��/�">��o~�����	��+�	���)��c�&D��a๺�|��`�ƭ6���o����6��;"��ۢ�l����������6ACL�����q�Y���'&~_~���Ǖ����>��:}U�~�?��xn~n�g�x��������!A�|L�;]���<1�퍉���!���٣�O�G�������~�3�_Jc�g�#�yW����|}�,�_��A����i;߿������J���8��s;�/���vp{Q�r�������V�x]�rom��J�7ا���nN��u��Y>]KTY1�oim�"����l�w�gz5�E���
o��,���˘�3������v���A� �n�z����B��gb�g���Vy�+t�:�9r�М��h�(���(�_t�~��P��(�՟
S���T��3�jش`��$v��Q��7(����TykXE��	���o	#(.K�Q�(-=y�h���*�|3*��4O��3C�u�)�ko���{�ꪪ�"���'�(w�D�n`�~�Y��gZ���ZVWM�.���CdǇ�+707
��?�������xc��i�%u��#~GQ{(B���z�{6I{��'�����p�Ɔh*�闋�-�����es�'0���B]��/d���A$�UU橬���ڥ��ʠ�SS[1+��{�|��P�K;0�T��؁Wo�}zR�����_����*��dnJ��3���yF^9q؄q#b^�u
��l��M�5q���<c�/>,�s��х��<EÆ��D��}��܏�z+���1�㆏��C�������,���L���^��O�W4�S���G*�վ"у��@#���>�b�k�s��Ԡ��{��Y�Y�7�HI�шU�8���*r�8�=�Y�jԶ:8�SZ>3�TP_u�I%���ӎP:{M<��,�@v
�ȸ\�~9�/���!�{��&~_��ω��EB��mDe�N����RB�X�ڣ!ytU��ɞ�j��v@^� �QHz~�`D��K=��F�xy�`�bk�{r��cSXd>�dH^����=�'�<!ʑs* u���˫+��3;�8�<����+�����K���˼s��E��4��Q�����q�Q-.������w�E�?q���|z�3��O���*�q}i��]���e3��C��ǯh�+g��2ߜ�`T7׿��� ݋I�!��/�]�/�:_��Ұž������d�ʫi=���#޺�ɛ@y.%c������t�`O�4}z���0�f��OM�u��B;^x[,�?�������fUi����J-.�[]�:,����C�&��ը�c�����1D7�Gxt��Wt 9v.��JI�(3�[&��A�4&/#�^�9渶�0�b�\�|�D?E��w��s�T��6�u��?�t�Z�d��<��t�����tv�:�@�ҀP@�e*?� D,!�
�(%C�Y�:���� 11 �' f&�ԑ?����!,=)�^�l'����Ux��X��-��[��F�_��c�bγ���n��������\;��Jk��fޓ�!b�N��K�,K���v�ϻ�{�w�q��d�GӺ���&[u�L�����������Z��/��_�o�����_�|p��}>f����;}����9�!��̘��9�E��<�[ b=��d��C�E��c�L<��4XG�zQ��.�g��An;P�-歑�� z5Ë/a�p�a]�%l�wG�l��K����� �ƾ�����	���y�T��خ��s��?�����LET~��A�^�b\`���	�+���߃j���V�eؿ�5���7B�޷�W0<�'�G�D�X��,Wo�(�P�.Em�X^���[�Ɠ�eS��ۨx��P�h���X�2Ͼ3[�����W*�[T���L�:���PK
    \O�HcP��\  �  /  org/jnativehook/lib/linux/x86/libJNativeHook.so  �      �\      �|U�8>�L&i�LZ�P�j(-ek����-}����<��6%-��mZ@Q�E���Uv�]�(QPQ�Wy(OQ"�1TTĊ��Ϲw&��)�����������ι��s�=��ssg�ᔬT�e���?�l70�`�?���f̌��c�g"6�u��A�@C�Wn���U�N�0�� ����C�1����/��O1��Y8)�3A~<e�dC��|KҢl��p�`�P=�S�v�W�����ȬguC��"Ø0�_���蘪k�%�0s�!Bυ%�0\3�y�X�*�Y����Mx���6,H��2�)�K��p�N"���$8Y�S�8B:�� dB�RЏV\��`�0.@�l)/�9��	r!�)��!L��')�'+��H�T����K�E� t� �Tq]a&�rE�,�]z�Y�|�Ե)ww�|�����8v�����_;���]�/nN�~�È����ھ;)�3}���yߒ/�.ڜv˵��N�����_J�~f��`�?��U���Ĩ�4.[Y�Ρ{����|�nY���'3��=,��\��7����%���nz-�S�ŧ��_��^t���|[�?��x��7�ڟ�!�Gvǰ�6r^M�c��O���UsX�d��;R{�4*R���;a���,���m�?��xp-k��9���ߙ���e[��u\�����R��!���?��/�/U��-�?�;��� �>	��@_��Հ���e�@&�h�~~ }� ����T�pu ��ǚ!X�m����΀���������(o5�O�g���� �� ���7��_����� ����@?<��� ��Ћ���~b&&a=�
�A3���3@_��m�·C>&L���țs��cz1��;Hǫp�o �v��
��F�>2����RS8�d/�5��>�w����o�(��+��f�Ǵ#�����o��}
�4�@�)���FQ��p/�ו��	e
Ѿ�a� 埅����WE�_P>E�A.���3 �BP�2�>����X|FH�9pv�J�P�J(�CI?Q@o�_��0@Z%��ۭ��_���R��؞���!<�1̓R�D��`�L' ��
��,��[%�!�m�/����|��9[� ���>�y�B_"�+��1�9G|���_������p>��g��V�|�V@���~���N�U��jD���:&
�{ ����	n��T���%8�����z�mt�F�!(�ʻ[*�#,�{��?�u
�����*+
j���΂�������@�d�.(�W�g��8��9���++�9����4/xNAќBdPX^z?���
�%���{S^:=���^]8�0��2�J�x9�\Z��kg�/��^��TTU�V8K
�3��ºZgiyAy��3
� �W3e���d{���rnZy������zFAYE�����Y@��U��L	��1�\��eʜ"{���������ZgJ����a�}�����b	3�>78ެ����4��-�a��S\���BP���e�"e���� ��ZrՕ��U͛�Z�,,O����f�s�<���I��B�]V�����"�QYQg�v�T���*�
�$D��Қ�Bg���n��B����QPX=�Ɵ�3gn��+g�:jLF�؊	啅��P��YP,QPU2y�ˉq�D®�^Xm�����`��Y��-�$dԞ��r��f��v����eرz����Y:�^YR\8��϶UV���%�n)rQ_A1@�%��JQe���Y�fS3w�2�������I��$���fՖ;K��K�f`���r�_PUY�Z�FD00���*8X,�A�}�b/,�& ��*�YY�ԒF��B_)p��A�L��騕��R(kta&�ٝ�R�a�HtV�S��y�%�B�Q�����ρ�.��[@�f��j�h���.N�G$VU�Έ���9�s�L����51�~�
֔q�QZ�&_¢B���W�
̩�,�Y�D�R�1A&b	Ad�w�c����s�}Q?���BH?YZSY4lXA���gU��;��k�5Pl]�s.!��t,����+~aQ���6�T����8*ˋ��GLj"�	D,��F��WA5a�!u!M���$9�s��#�&��̛0��^=��!�M���3ӫ�Lb
9������@����9bo��Z���BJ?����G��`&i:��ҙWZQ\9��'H���]���X����6+MI�=DN���^��gյ`~�%hz<ڈD��\1;�$�ګk�e-�� vJ��gØ�M��P��
e�PN*��+,(�^SC�#�TQ̤ee�L*������⽺-���rQ������'��BG�\͏�_�㘗�ԙ�z��Q�t4�����
	#�jf�;��|�MZ&�</��8K�W��+�y=�0�^��axP�J�an��)���x8�}1��1��*ư�ٍ1�u�a���0�1�0G1�kr�a�p�is�
��`k�3��>ư69���a:1Nb��Ú�p�a�0���1����>
c���1�����qÚcX�X0��ac� kb�a9�I�7�AQ��F�1�5V�zX�`
�F�aa��q
�L�Zd�w�:c���c��1�sb���1,��ak�z�{2Lư`��yc�0��a��1L���1�Q�Ÿ7��0�vY�����:hg�GC;c|=�3�Q��Âi#ư6m�� ��팱�cX���&hg����Ú�c����1�5�	����1���am|�Xhg��A;c���80P�S-,�8�a!���fh�o����������ָQ�B܌1,0c0��mư��1��,π��x�?��\F`��0�]gt�L0�G���e�k�(��mN����S&�:W�n�v��������q���؎c@..�����@;���F��XI`�yt�^H`�t�v:Z�+H��zc��w:�<���Q�-�a#0zSn}w$I���a!0��;�!l&0�r`�:����*�#k���^Bw����Ƣ���w�-��Ƣ� �'0�;��Eq,#�'0�;V��Es�#�'0��8�H�	��:v����О	�'0��8J�O�y#�'0V��!�'p�gI�	�Ust�������Y�?�[H�#|��%�p��A��~��?�	���?�-^L��z/#�p�W��Gx�W��G�F�դ�N �:��[���?�f���G8����f���?�g/"���?�?���'�'�a����>Jڟԟ���'�'�1����>Aڟԟ�����>Cڟԟ�gI����iRw��'�'�E����ƦtxH�	�!|�ԟ�ش�NR�_6 ����cƦv�>@���n#06�#��B،�B�)8�n!p¸}�QO`4�P���;����MŁ۵6F؆p��t�[�;��i���ƢG|�p|g8O(��A\��ҳ	(��U�xmt��Ð�js��8{ �͓)��v6��ڹ�S�������g��E¿��l�j�b<|ۚx��f�K�	����異�؇�D�]�B���BG[ƊP��� ��9yDH�A�̔1M.��9'&,�y� )�D����e�ͳ�,+B��"���un���]���ݵ`�|���⎊QԶ�eBӗ�=_�#��^'m^�<�]y��W'_���ZAG�()[<�������u�������!�[;UM[�v���>��p��!�=N=m�l�̩�|�����M�K�WQߊ]����]mT�p���P<[.�6h^�Ҽ���]X�T�o�agk��kHS��M$K��k�o��ꓞ����b�f{���nov�c|��캄�ܱ��ϵ����@�;��+�{���6�x�;��O�-�v�o:�!<���<c��c�1#08p�Pƒh��~����6�c�9ݼ�y[\��f�-�]SrLd�[;i����@woH�r��1R��DK��$Z�r]R5�05�'��p]R�p�u�����@cpk��bu2=G��[�BVX�h���u^O���N�@B��Q����W�6r-��%�vm`!:E!��ق�D	S�t�@N��~D�x%^&�6�(�3Q��1�"��v�@H��x��n5P��y����{�/bs~Jl��v�`���
�&7�sE�]
:��硇k%'�n�w$����_I�?ɉ� �ӟ��U���I6^�{?��\�
��I>�
�J�uWA2BI2��6�@nn��C�{޿������ ��q�y1ݼi��vT��Xr�����k��jN�+�״�m�̃b�Or�x1���{�'�O-G�a`w��0`e��wq8�2��{�ȓFH�.��S��L ֑t��������X�PE�����[[p��>�l%���O8�M*���,���z�;��=��=ʳ�g��?�g0Ȓ����Na�M���ij����giV���4.w�؂ӁfwdE2�ʙ��IE�"S [Ԥ��L��i�DC�����^����1aM*S�T(�@l`d�qgŘݫHw͉�jb�|��k�����1J����l(烧'k��s\����郻I��Kw���`Mm3�i��(x.��mv?'�s`�<�sw�s�Q�[� �������G��6MIn <?���q�Y�s����@�P,��y��a��]]۠���.�����ͻNѼQؼ��;нj��¥�iND�MW1M6Dq���ֱ咷_5���������s�Ѻ�5s�9����+���h[��Z}h�/i���R�Pr��v��)�ܾ����ej��a�gd�g��y��
����j�t�3ߡ��2�D	�^	�$�����UMs��;P�:(��\p�F��{F���&v7G��Ԍ���;����`v�!�W��%�ܨh�H���l�8���
�r�q����B��+[)]�&	�!~֝Ѝ�S��_?}Y=t>T�n�v��w�U��z�ʢ<'�E��*H�;ꧠvEJ
���vň��d=Ev���Iw[y=�ӓ��f��������i����Jn��f&+[��oP)'���jN\N)]�损}��ܳ����}8@��5�C������)@YK���zV<}���� u���5�=P�2At��A�I�����0� �~�Ȅ�e�O��.�fw�Ӳ�#����]J7���}
��:oQ�62U�F}�[w��7n�Vy8Xd�B��	��g�u�;�:�-I�0���J\��g��i5Q����.���j�)�J�K���ֶ�Ry%w�.8Oե��5Yp�+�k��Xr�P�ޥb)&�������kO�R�$u�O�/Jp>]r���`?T����Jy���[2�}-��vᾱ�݉�q�����ڜ6欴=L������=Wg���B(ٽ�5�_�����/���-]:��<�x`���#ϴ��H�����R�#�<�N'�q�=!�D�Y�MW�jOh��k��ȏN	3XO"�8�"�k7�S�;�"�����'ݕ4�
�?i�;Ҳ�T�N��y��'���B�̳�9�'�-�*bb�(�Ȓ��-�X�	���I�*�7�L�[�.O���N�
���֕1P�<��ԿE� KӮ�_/��挮����a6Z�o�~�ā��"�!�C�XR!�t�oA��z���Х��w:��.҉�/"R{��#�C4�^�)(x�#���^���w ���O���~?�.����w��{灸B��/��c��_\����1�K_��#֋���.��y�was<��2�����=�_���R�Xٯ�l���!ny;A�WF)iA~�Nu�M�NM� ����A����O��ENߨ!�T��xϤ��|�>K6����,��s�Iܹ��#�7Qt-o��[���
�1��گp_����0,�'�o�q
�H
�t�(����J*��oR�!�e�GNH��y+��ܙ�ǋ��u4A��#�FS�����
��RQ�!���Ug1��I?�Ԩr��@���3tC�����(������ݴ*Yd�Xn_��ԓaٚ�F��ݤ"��Gh~�VIa�[������I��ͮ�,s�L���)'�m eû����.�Lx���[��S[/��6ϻ�i�l����&2\��M:9SC(��N����\�uw���P%n���م�J���6��z�H+d�ӚfLN����a�b(i�P�}0��M��*쎮A��p�zj�%M�A<f�D�i�� d=TҴ �$/��M���W�;�$,���S��F@v��m���>� ��=B[��w�ڦ/ir[ �i�F{���4{�����i��!�,���
XӲ�)���g�g%u��z�[�(��iϋ�i�����7/w@4B�im+�jJޑ7.[V��������T��,�v����ft�^��qxA���r�U`��Ê��]f�aP���y��Fa�mA���@�ӣQZPx���b��Ǽ����0�O��迭iU�+��p���"�|*���TH�l���1QT�ER��뒦�ȑ�
V�9OK�R��O�?Q֫�5�'�Z���¨�N5�Oa�*b��~��;Mkd���Г�y���j]'γ����I�hj8���e��h����z��� �JBO҆�����P��W���)p����u�=��X(��@$!�w��BL����D�δ�`��8�qFԃH���𢲛~���g���&&��*��hjPk�ܰ�[�.�����bp%�V�55|����q�����8�y6Ӱ�i6& ��~m�CeWٗ[H]��9���B���&Lk�c̒�pc)�'@��7��sĲ���Sy��&��ף���UR��W`�	��^T�Ewb_*y�=�<��NC$��,�_ Kdɝ�(b�t�1�vc���7J�F6�����6�TĆ�(���{8[�v�D4�F��y11TCZ&����nRҙi��:�V�H���� U�9������~��+���-����$^K���2@stH������:b�����9y���*�A�9��P��N���(}�2_��W�|��$��z�j���sP:I��9�IE��A��T�:F��HSʃ�w���P�@>��a�<����[@�Q���g��j�ue��~nUy�yZ�D`p@W�s���e,����w�Q�L�9ƿ74�弛��[�1{�~*��v���2� �*�X����6P7����I��1Qь*_3���a��-�?��|VοV����e3���lh3��[I��?�|�qa�t\��Y��oTh��w8X�y��;p�ဓ��{5�p�B#Ҡ"[Q ��'H8+"C��������LkA�djA��	�Pcud�h��V���p��c���tDp�6����0��б�	\"�M�=�q�q�Gi����5�u��ѻ[Ӆ�(ֿ��g�b?F�y�*u���ryh���z���<Y�"<<MǸ_l�E[	�l��l���c_��H�Oh���.�e3�v�2g����������lqO�z}2�$�om���^$��Vt(�';Ҽ�kp��Â��U���`٧{�U:��ɼz� �W�D���$?C�ʳ���4�$t)��6�pU� 3�J�ԥ����wZKM- ,E�Ζ����ɘŠ���|�Q.����&���n
�*�81�>�J�����v�����QЉ�`���S��2S�`��/@�Ņ�OVx�>�����%*pu�T��Љ������7��GG�O�����8�۫������4�ޡD3���!h:S��|h�����u����r4�����H����]$��~o�L��1�����8_#g>��� �_���ڱ�3��d�GΡC�4�?��4�'h�E:�K�#�d0�a��Vr:Qr�0�9F]`�n1Lj9,�4臮�? �7�^��s�+�����<�`�Xm�}N<�yoӶ���	�8lyn>L7c���l���#��0�<r7������35;���ܸ25�aE��H
�a���-�lD�,�+9f ��
1�{��`���1�_��'x��mH�\�M��ӗ���HY�mj�@v�7J���[�2�3t�u�� ���!����ܡ�� ����ʬ�,��_qwc�h��cϓ��l�Z���\��w�fa��y���5(tp���ˊ覂 jd@�:J����C�6(g<7SY)N���Ry�ǻ-��*�Z��l���T�aa�w�^��=���1Oz��zF.�*g��3�9��	3Ir��Ż���<��S�'�<��J��:���QΏ%����?"HC����	��QD���ܮ����Ƶ,[��y.��6��γb9���_���l��L΂;�w�������ͨɄ(�V���hin�[LN؍��1�3�S�&���fW���O;LZ���u���ł�|ד1��KM�jz�ll�Vgjs��w�Nʫ�EjD���=@r�#�iI����D4 vi�5g�P(� -��/�;�B���"ہ�N���^�c����u����O�`A�1E525�}��"Lk��Gl3�I㚶��h���`j�3C�[�1����	���;`ZcӘ�X�B��g>Ѽ�9"[��n�h9��6ð�>n]���5����jOC̑�&CL�	�Of�1��Ә���M���@	��	����#���}�c&��m�]�c�2�� I�4�{N���{f�����;魃���М�0�?<�f��ixd��(mKcz�ͮc�I��!��)Wq�����+���V�_y��Z�im�#m2�U��Nl/�"<=��6s��G��WgA]vs�1W�ԺQM��h��r'�9e=���ּ�m�(�6�u�Hv��y��#t/��:���i�隌�QⰭv�GZ�p�;���x���JlJ&��sXx�9�yOY3��J�Y$}�s������MZB|zq��X(#t��Oa}�κ.ԥ4�s]�Zw�á�VR�0��n���B=8��N���GUþy���6���>��tֈ*P�;ٴ�{T1���>�Eu��:x�	d���~z����93q�b�c���@<����@��p�����n��͒v�����@;rp�����>��75�Ě.8D(������y����|[Ɔ����4o����t���hQ����İE]�c�E�9���~�g�M�Y�W.��Kq9��R��[A�K��N��k�WwW\%�Ʀ�OJz�!��zN�5h�|>�������E���9*`����yV�M�C��o��8PH'r���p�J������3J1	���&%h���{�y_�����7�O�,mjw��
y	�U���wP�_Y^�>"o�����ޝ�qW!/�0�����m�w�R^�����"��':�m���$����1�}�CKd��p�D�Yx��(+��w�����x�uD�?=���\V�uK|}�;���؏R~���^^~2��ۇU�� Va(x�,w+Vc'ψwx6쑤�kejXO�Fo��16�dv)|��aC�-w���|S�c|3W±m6���Z�sP�{ʆ�͆\�5�s�Y�~��t�i�����V] w0�bxH�T�4��PΕ4�߉�	������:��a���M�Gv�d<� M���/\�5�1��}�߮�qXG�H�Ѩ/�yO�[���ͣ[~��F��ZƳa7�Y�f8���ɺ.�CL�������ի�@@��T��5ʘ2ֆ���H^��d3�46����k+��YR��4��Jܪh��#��9�W�Ϻٱ�»_��t35���ok35nÃ�_hM���P�Qh0�S�9�(��<�����.[��;�z1�^��~G��^����|`�}'_���H���hlH�
�}-.����t���s�3mI�0m��u'�]�@!O�e�ʰr��t6��u!�Ԁϖ�.hM�ȅ���t]�M��E�y�*\����)?�'���x��¯=���7�M�F�d;}:�ID5JdU���[�z�6\r��5
��i��q(4��|G
�1\_�̙��S�A�a�
��Ni��h�AQH�=HFXG�����/�YR9���O�(#p;��OB��f	�]e�;�Q�-���i�.�lqs��`2�
�*̃��9�F��'��܌����k�>�G@ϒY�/^�)ٮ�\Ι8�J�	���zV��X�8o$�ɳxuD�{��l��	e��(�9�z�H�+�No��|<7�YE�]uXG��� �>v�*�X��|�.�!F���D�S^<�y0=@\��;9�H$KM��@��;����}��p��-?xD��մc�[�DK.}��<{��M�w�|d^"@wk'Gw���[Eq�W�N�7���++�
������(��U������ut?'j��������������q\[�ir6I��$����T�?��S�F����_��V����\/�yJ��)��!��P�G�#j��M�?�����	r~_��*��&���1$�)������o!�H�?\��W��	$�����B�O$�wJ���|��Ǒ��R�9�"�'��o��O��{Fm'�_NlϨ���l��d�ͮ���ӗC�o�MN����L�������i8��=j������v��t�{��&"����y����v�;��s�֢�d�[�+�7�s=��qG?,�V^8��<f�O�FQ~��ZY�n����O�Faǘ��.���;(�<��M8��21��U�<[dY���ҡ Y�=T�=�����V����c,Ŀ�g��o��_�d);Q�{��}��R��9"e~�Jʷ�RVx���[� �����J9}�WJ���?&��VY��YY�6�X�?�9 �n�V��뽂ވ�mO��4~�,h�W�zp��^����	�L��c}�
��2b�u��<@;��'��K�~���f�]簧�#�Ri�z>�5��׋�J4�\�6UB۹^F��������_��	�`�����V���$�`%�^��%	s(�q��8U���+a��y1��bJ���|)AtbU�����5�.�Pˑ�����xI_�LO��V�u��� |5A^Ǎ�<��AMߖ���%yޤx���ޛ�??Z�l�a:�{�|�cg����IϺ�z2�Ru�U�!4׬'�I�Qɞ�ۦ�-��*��`j���5g;nw���ͱJE�T�����������o�Zy�K���$\�.��^zr�CG�Ǖ4��cM>>���u�x/A0�#��&��s���H������Wi�'w���25�O�D-cM����2���w��� �8`֨�3�{�|���ηs>�;߮�A���n��͔q6�L�c�����&���Nz+���U�mc�����}߽��Wr�πxVS�6�p�J\�צ�M8����q̫[J�N�v&�P��'�ߜ�M�U?��钶jA�A.��N74�15�%�� �3���5�J[�W��f�r�����#5��,,��ut��������STm���7p��H�:իa
DR���A� R��φ�4y����˟Z�c��b|��a�W+毇�0�R�Iv��_�����$,tS\0I<�f�1�kw�=����CѮt�H��y�TfvD����hf��_���|o!���Rn7Tq�~��fg{�i��P�7�N�Nϊ�ʧd����WMyoq��i�N�Mk�6�D��Ӣm5����6����ߕ��|T�%����H��Q���6\���ꐨ�L��Q����tO%��z�U;NKd��\�:#Q}��;*�k֥�	o��;׵�es��L��n����.���+s��3o\�����h�]����9\Ɗ�W�2���P_���2� =���W�S�\����Ѐ��N�ߣ���_�?؈� _ߟW�)Ɨ�B��B�'ſ�������]Q��>���)�7���0��k��+�Ȼ��F�{��S�&z�{��WY=#^�^]�oU������}�.#�H����[�}귎�u�-m�UY=��(=.#˗;�Y]Z1����|����x��^c���3q
<��;3Fe f܀|ixF2�]Y\ZRj����222�cy/v�Ř^z_�7 I�uVK4}�1^��F'U�BM ����2:蠲�<q��Fa�u����+��+�}��/����Ғ��<���5�צ�e�/^�P���J/��Uz�?(]��nIi��!oN�]X]�PH����0:S�L�
�^`����r{��Yi.GE��E���񇛑A<2��A��(&�=�wB	?�uR�E^���Q�,bp�Ԟ�p��˖��#��֮_+��#�!����
����\A�6��]�P�`��{� ���5�ɱ��7gT���˚'��7;��1������k���jK�vF��0�7������љi�E����4���5s�(N���1f�+�G�~(�+�x��@�s�}�YvN�"��(Klߪx�_�4�J�ck�Q�wLev�e�(x�5 �|s8�{q�WLW,�`�!F��j;� &^b(��h)�����t@ݱ��Z�5�B'I�5��=���|AIy%(����^��_V���Y�^�w�j�`���l>����|��2$�: ��J����L�pV��[��u��r���>iF�2�HE��l|�Yz];����Nbh}fE��
�Î���������)�.�T�̪�1��/�� �D�3[  �7A�,���f�"��fRXBڴ2<T����߹���/d�a)>���+�ҷ'�+g����������5��p��`4W�1���ͅ��3���*��������a.	�
��OɎ[Yv�FGC����|����f��������^Y��J����͉ 8A>1�vr�$-z�N���3**�훱��<`�|�:~�������3��tT6�@����GW���b{]3�.4tH�߷@��}�ck��(5�EE����cH�i�	cq�g�[����\�ti��oU�(���Ⱦ�j~���~��������ţ0a]�q��+�� �J�!��@�5Xw_���� ���Hw�_�7K.W���m�7W��LO��d���g9���j��.a�b���ؗ�i���Tv9[̮`粯���������#�*v$�&{7���̮ew�ֳ����me��F�~v��j3����Ƕ�9�vV��`��;Y���ؽl$������
�6�=�&���4�=��e���
�#������c'��Y5�%;�=�jYkdO�ײg���oY{�g�c����t�Gv��Ndf+�_���Kl+���W�c��bؗTv��Fv�j0���?�FˮWY�V�M�F�����ݩұ�̠�(�E9��j
��*�=�
aT�a;U7���f��T��/����Թ�u�T}'����\ͮP����y����v��'۪��nT�`7�G�[ԙl��aw���}�^�~���Au
{H�ž��~��f?Q;�O�e�15�~���=���~����N��~�������Y]���.e/�g�qw���T�8�eg�,�X���R�{ˋ��e�"�K���܋���K��q�+ܗ�W��,�q�-+���׹,op�-������2˛�˖5�r�Z��:�5�z�u�n���{Ӳ�[k�ĭ�l�Z-[�M�6n�e+�ղ�k�l�vZڹݖ�^�N�-�.n�e7��e��e/���wȲ�{��6w����e?��� ��� w�r����.���0w��w�r��X��:,G�S��Ӗ�3����-s�Z>�~�|�=c��{ֲBc�[5��[47�[5}�m�h~��/߮��whb���~�.M~�&�ߣ����̿���ߧȿ����&�߯��?���5V��f���6��f0���v��f�����f(��f��f8L���I�Ќ�k���d�KM
R���I�=�t�C���Ҍ�Ok2�3�,�k�h���[�X���������糹���"~�������|.�"��-�������$n9?�[�O�^�r���J�W��y���V�,���7y��繵��[���|���s�|(��7p�y���6~���p�x+��O������vn'����o�v�)�~(��ƽ����wro�#�w��������� ?�;�'p���a~$����p�󃸣|���}���}ħs�O��S>��������0�>�;���N�ܗ�5�I>�����y�X����N��r���3����|��-#w���������7s?�}�s|4�#ߗ;���~�{p��@�g��ߛ����.��~�p�������=���~A��z��I�X�'��������i��~I�\�\����F�k�k̯kW��о�^�}U�Z���M�^�m�z�v�z��m�z�[�ڕ�V�;��'�۴O��k�۵U���M�S��z��������h��ޫ}Z����>�귵ϩ���K�_�o��B�A���C�E�������K�G�K��k_T�.S�}I���u��7�ǵ��'���_j�T�ԮQ�]��hש;��է�ԧ���3ڍ꯵���h7���nQ�ն���nU�ݮ�A�M}Nۮ�Q�C}^�S��v��S�[��v��y�ھ/���tL�b���]��Ku��u��]�[��%��/��]�{��
�s}_���﫺�}_�-�R���F]q�&ݴ��:{��-�m���[u7Do���C��ޭ�G����p�wt����F�]�����\��D��9�S]���tq���T��uO���Z�\�=��Wݓ}.��9�3��'c�	�9b�9b��2D�	���	�9{:$,�L�!�됈�oBF�~���ِ־߅0�߇l��CȦ��B�b��=28������!����j�z�y��3/�k�K�Z�R����>ļL�7���0���i~U����>ּR?�����>o�'�Y���Z���M}~�5��}��'�Y���i��0o��Ys����}��S�����g�~j�=��>{�=���o�}[�6��[������G��5�G����`>����� ������o���~E�����O�kb?���L�j�1������c�п{\�*��~S�z��I}��+�˱�������Q�N�o�wF_��k}I�o��~g���������}�?�{�?����G}e���Y�~ҏ�שO���^�wAM�_���\�5����|I�yQ�fi��̲и�B�G����l]�=t@t{�����fohd��п�}'tq��зb���=zs��PW���8�苡��?3�63�|n8���pHs�����K�{���#���k<�����S�5�i�>�|m�D��Sͷ��4g�4�>�|o�B�����G×�󆓚�_i:�φ��)��FVx����b#',1j��F^xѨ�u�K��e�^XnV�+F��Q^3����0�uc��������SXm��4^#�1��{댑�z���uB��za�1J�d�A�l�Q�b�Ih3����>�6c����Wh7�;���Nc?a�����'�1�o�2�"�3�6�Ax�/�7�*0Z��F�p�8Hx�x�p�8Xx�x�p�8Dx�x�p�8T��8L��8\��x�p̘ |nL�0�����d�Kc�pҘ*|eL<�t�Ø!�2�N3�3�,�k�h��&|g'|o�~0��s�����\�'c��i�~6N����A�E�m���`��v�Ra��E��2a��%a��ea�u�p�u�0���p��U�n�k�=֕B��u!���0ҺJH����o
)�5B�u��f]'�[���(k��i�(dY7	����1�-�Xk�`�n�Y�	����xk��c�!L��r���<�n!ߺG�h�+L��%L���X�#L��
��iփB���0���Pd=,,Ox)���r�������W�?^�Hx-�cae�'���
o�&�
?&��\x3�aM�qam�	a]�������p��1�C�~J�~Z�~Fh�Z����-�[a���p��;a��{�a��#�sB��Ga����l�I���S8��p6���s�(�d^�s�yc�lvS����s���Z|y!p�����3w�Ԙ �D],˰���	K�F�\��L/F��eY$P_����@�7 ��@}P���PGu_���X�����:� ��@}P�? u<P�
���� �����@=�� �@=����@=��껁��N �D�	�I@��)@�
�i@��@=
�3�:�G���6���@=�s�zP�uP��D��ԓ��h�~Wz,S �Ӏ�j��6[��� �K-�_�z����e�>u��y���D	��������a/3T��i�c�a:�	�hc!��8��!��p�Ǌ�xH�+b�Bl���&E�j	B��S �a���B��p?���2N���� �J;g}�Ѹ�Xw����*U����oT��U�������R��oP�I�L�~1�a�5~��^Epyl�P�<�AI+@�J�VE81�}������;�� ̾���k��O?
���I�w�����Xz�2�d<0�'x �����&�y��_4�goZ4�������F�����ח�B_�v�]��p�w@�����6�m�~������`a�믈������������������B��A��Z,�b�%�?C�3�
|�����_�/g+nt�ϴύ�;��do��<�;������W��B�t�9޷C�fw�T�I��By)3�w�ٜEw+�J��<�[���+���Q��*�R�����5Z�S�/��B��	�3Ċ�%�-�'�:�wK_ƪ�������I�S,�$s��h
�j����ӌ�.��u�r�l�OO��3]����FCaMP��b{])$��ӍtsaUU�|�o,u�S][rTV�k*k����A�m�#��%8�����K5�z�������%����q��F��ӌL̔��`^�ͯ�&���V�vgmu0*���u9��<���Э�W)7a�'8����.	��jo�tS���EbhV24����7�����ʛ4�5�o���a@�����BX�������N���H{�	������O��S�@����wx�l�@8
a��B`�$�f	�A���o�_��C����A� M�]@M%I��<�4�{Ư�^��v��kc;+mc�7�|�4�K����^N�������Z��Ny���%�?W1��^=W:��8V��_ȡ3gɧ0|�<��	��b�r���$�l!g���K"#�|���H�)��]�)\�g�x
��y��[ZC�,�ڨ��Q��CP?�9_����@7�r�݉'��<%�eQ�,��8��P�-�����ے�<LQ ��^}'~���>叢�/��(�z0̳gA|�?2=l�*�Y�} �g�Eq��!�q��Ϣ�F�W@|�������yϊ�@�j�	G='�9?�? �/Q��e}�q?�4�7B���UQ�5�㯋�c�ܿ�Q<�@�ua�>�x(�+V��Y�W�bz8��&�A��STA<p�(n�x��~����=��� g���?�A=O�v�>��gm�z�y�D��ސ�M["o;�]�w���A>�� ���q#�DH���l���c�7p~��i�����g����K�L�Nns�uw�<(&�ܝ !�1QďD0���Q�(U'	a�D!¥�	CG	#���!y���"d%
�t�2N�$�H2�I��Dr�/$'	�#	N�`����, S����:��x�eV��%]/D$n�w
��]�.q��%�&AjR@jZ�X����\P�~��c�/y.I0�	q)��d�b8��9~������(�c�:Qsq%Bd��(�Ӆ�$r1F��$�jH�	��%�9L�0��Y�S��O���!.G�(X����`#%]�%��d��D�S����B(��1@*å#D�"B1��Ԧ����22dJE�3���ज़���MJh�^��IB\F��� >"�AcqLH�2��!6�*$��iBz"s��4!?Q��(L��R��?d�lcSB+#��r��H�/F�f�(=Y�o��|��|�BB���xYy��P���W���B��0���rb����?��e��Ͽ:�!�= $L�]�\�>�C��2O�-�I�¼TH�����Z��������e��	'��ӤQ#�a\�3���8/�]��kwCZq�(~��������laD&�RȘ�"�R��!?I��$LK���H�<Q��|������=�|Ȩ�����r�0�d��cSz��`800�����IBV1Y�I����!��	��t�I���0ǆf�����f���REeSL#�d2��GZ�a���(���ӎBZ�"�)g ��f)ƒ�#��)��O#�y*�.>	r;��|����c>ڙK=F��څ� b j��.�4'E�a`�\f*�F��
(ۼ@�R���iQ�vg�<Q��y�c��v�e��:�.�n�x���0�M�4RX�>��E��A�6�\d
ŉ�#M(O��%����� C��4���ܣjտ�)y�d���mu
���8R�+��	SR�i#���ﱩj�)#��'�hHMԓ�Й�$̓���J!_�J:<`��
 ,_��By���qz!g���"LI&��i1�i$t�1�_r�##T5W���ʏUTf�9�B~�0%��<�BU/RD��l�x^y�u���N��E��� ���	0�x8�\ai�4�9t��N��\d���^.Y��b+���l\�:�M��K����&��X=a��J�/C5��,��c�9��/E|h�;ϙ(k-����/�>+)䌖�	�mTw֟��B��n�3�|mK�S�i�Bq�<Z��1\��lP_!�'i؇1Q��;sfX�^|^�T�̰<=��8�H"G
Q�t� e$_)#͛!yWt9�CY�/�"'�$\�/�{��v����B�H�Vc}<V�z���l�m;8��3�d0�'��(��i�K��t�6���?R��$�pI8����0�ȍ=Y�:��8��9���L&8�8��2����w���R�2�H�dq�*��ǀ�E�X�qb�Y��t�Wq�ڻ+_e�w���&��"���X,�s��5�+!�+�o�G���k`�(��oa�B����?��B5I1j2d�xx���y�����V�#w�_{�s��L!��$�i�H�0e��(إ���Ƅl��>��0��� � �hB�Ef�e�d�8�9d��(���B�5Q���4M�IQ�c��"şd�^�y%����B�KUȖ釖(�a�xN��ì�X����q��E��� eH��L�xsK�3�cz�x����!��
�QɻP�؀��2��J�� ���-�ϖ��Fl�7	����f�%K��d�+�,!��L��BU(M�҂n䍑���d�	��rڡ��E�����M�M��Z(j4��ѡ�g���D����d���7	J���h���$	��?�l IH��$ӻ�L!#z
���,'	GtP�)��3R.�>��,/	i�T"y�0YN'��(0��TT���J�wj�� ��#�i�,XI�[�B$���D�^�>[&����Ba`ZG�n&I�fRp�4R�zh��-�\�"%�k��$=���V����^_��$�%�k��t��q�a=��(��ޮ�'O�޶o�1I����	^�,���=��C��6aO����
u�U���_��o��|/'X��:H�`�k�>_��%c=c&)�����d�fFj�����5�>��z���nm�*�W��r23�6�F�]*E�и9B\t8�ZN�L�)ﲑ�r��9��R~k)��7�2^N�P���_Jb�R��O�t-P��(�oH��$���WJEe�kJ���:(������Ǣ�_�"�F]�}�`�O.�´r�6�h2�K�<E4F����3p��<S��Da^�PϦl��;Ax��Uu��6Np$��/�H �$Ky(`�0�@Q^�J����3Y�3R���p���(��*�I��h)Ir�
ũ2�L��e˛dr���&U���)8��{A��TK��AS�.f�#dȪ�Ul��Ti�#�d�c����&}F7�����W3��)2��������������O��������㗥�V��K�R�C�I�\W�0?^+# ���P�	�H�>Q���>U������J'��������k�5q���d�k�.�b��"o%�p�#�yb�^���o�;������ ,���NG ��p��^�A!B.�u�Cx
�Rk �p�I�!��=�~�@H���B������;!�p�y��@��!R!�B(�Pa>�� ,���NG ��pk�^�A!B.�u�Cx
�Rk �p�I�!�7 =�~�@H��p�al��_,��zLKJn�K�W8++̓���f���[��J����4�&3L|��Y���;�i쐯fT��;
kL|��
@�����HG���ȫ��#��*w2�xڗ�ǣ�L|	 �UY\�,d�펂���Y�Gq�b⋜��5P�ʊ�Iх�J���J'�GyS>�k ��r�,�g�~ؿ�f�E$'�*c��0��?(LWGȰ����(L_0�kI������L�!����y[W*Ò e2l��?%�F��]�部+ߑa�7za�ҷ�^8����p��/�R��0�8��iE�p/F�S�7b0�|'	 �z1�by��P�[ �6H��3x_��V|�7[|0~�ء��_g ���E�
x�_���Y�c
�Z5+���T�������~�Oԇ������0�������ԧ#�B�o<B�:������q�:~ ��j�t9�cSF)��>g����X��f�����Yw�ꃟ�KP�jV���� �Lޢ�{ |���7��#|p�mw��>XE~?��)�ox��3�ӆw���i���#�
}eb���"��;�������T <�7"\�0GC)�4�Y
���t�
�����F��N����� � � � p���<@��L ��`54�Z�p�)�7\_K��#�Z_���Q�>�2N������p�Z�� -���A�WN���# �C7|T7�aN��� ��(�~
�i
����3�����˸燎_��'���X�^��U����a�S�-X�} ��C<!+�g%����r#��;���Fb�%��B�\���W��W�1]-�'�}���Vp�?�p=����y J����I�����l �X1	�6n��)` c< W���=�@�] �
>�0x�o���o��?�!�����ևa�K��8_�à�.�-�3P��a8�P����}ߖ��`y�	1�/�2��s���� ^��J�������|�&�7�`~e }C �o���������� nE���/��`J2m<�YM�#y��8�m�L��_ W(`������Մ�QD���MB��<�A1��d~V%��N6Nvv&&����rvf6;ٙ�a�w�*^DP/9(�s� ��)�b$J�H���,�`nz�x��ݯkf��@�������OU�TM������S尼sF��dg(��ob��6��#�;��D�0�S��)���3�a�
����=' _/���C��A���� ����A�7�B��M�#^��p܂)���Q�/1~����'�g�/^~L���ϻ�-��{|��/�}k����0���6�f��@�4�݃���<��[��g7X{F��>8_Ҟ���#�u�x���>���vq٠��;��@!�oF�-n����g��5��,_~n������1���#���{���;��ү��A?R�˸#<�t��kc4?�5��^j�#�g���W��|������O�,�����?����
���-;��ַ�*�ϟ��A?Q� }&o��Ü�گ�6a~�uq��x�6給[�V��W��crj~z�9'��,�V�����T&��Rb(��Iuܣ�iuԹYu̩���:&�1	eN��u(o(��^�2WE[�n�Q.+����k�о�Ut���gԙQk�*����2�SM�`q�%��̪�0;�����r�F�9�����ZW�\�\��M��ɒu�^�х�T/vNՍ�P��ԑ�v��j/��M�X��x<�	&�!�
C�\E(�W�2Y��qhY���ʶ���wŔgs�fS����\*i�<�3����(���!!�:���4ehH�PƦlM���4�V.1�,2���Ĕ����f����Ԣ���×�cmϑݹ�B,���Cr_� %���H�BP� �V��{@�����Q��N����/UF�K�26vx_UV�GJ��z�;�5ٯ��EaV�
rm8��iY�������#�2KA�'(��	Y�N�F�w��i;v���)x��rכs���]� �s�n��!��u
W����E�H�Ͼ���W)�j��M�F��}�>!A���!`t��3���z�b(v�S���o�CF��L7jK�cP�h�ELԺa8�3]�Ty����Zvs�֩)G��.�{���ūBBI��#)�(L)�Q��"[-�1G�OI�+,B�O�;������#aM�m�>�C)�5��p�6������&��v��*v�2��9�%�QO,)�
9V�m�`7/
"!(e�.ap�~n,DG���&�֐�=��Or<ց�\&on�3��\ly���dEĥ��,�:D��z>��Ug�:��9��8CI+��k��|�%)�*�o4�8O��r��Аt�ڧC~�b��玎 ���{�!�,���aTi��5{NG]�/�u����%��]q�'�����+D�)�������D�F��;\GI#z�8�8���ʰ�c�(0x�1"�Y%ֹ��>�����C����6�7�@��+�y��?��G34��uڳ-��[�K�6�]�ט�*�C�B&�u8A���-8w��$#�DO�4;Y�t���1�I�FRП�`�n��a7�h�f�6��3N�9�w�mhQ�w�����޺s���Aܧ´�A;S�w�]B��uܿ��ǽz�p�hp�w�����&��o���;T/�wa�E����4"�2��>��"Z/~�O� ݃�c���(،���}3L������tu*����#��Ln~�G�aZak�[������6��R�?��u=L�����W��i�!]��_at���������bt���i�^��D���}��"�
�ӽ��p?��*t2:�'�z!��t�L�ף��
a���+�?���_���t��)C�2襻��p�<9�[��w��G:ܟ��<}C��[�H�+o���7��
t7:�{�^�li�ޯqE�/����S�_�?PK
    \O�H2��TZ  h�  2  org/jnativehook/lib/linux/x86_64/libJNativeHook.so  h�      Z      �	|SE�?|ors���MQ�ChYJ��}ii)(�E�R�*�HS�b)k}�����n���Rֲ/� n(�eO �Q�?gfnr�6��������󾁛��;sΜsf��ܹ7�O�eV�<'�� ��8J'1|�Ao�zqZ����$e5\���K�S�3�o��0HQ�&�t6�G�ϧb|Y�/���SR@���yʑ'@��-J�y�*0�Q�'�ƾ�O8KG����w��'�rTD6.��'�WGF�����$UE�^�q����͹pU�\HXRi�=I;�Ő��eg!<�=X�Ņ/�RU�-��
O��=���WX�&��At���,�����(3�8R����,G:C�G��#�p��ct�cX:���y���,6����D���|K�����3�\v��- *Ӛ�+�R�O���"VG	�>t�ϰ�ζL���nշ3�Z/�0�.�����Å��k�wL���s�Og~��}OJ�W���L�����~{�N-�������{�>;����X7���^S�xy��i����s�e3�t���+���L��S۱��E�a�w���\6���x^<ӡ������'����+��x:�������r���{���?ZV� ��Ř9Z�j�#���٧�������\���8��ݑ�M�^��󵼭M�S������u�?q;�6폝�r�M����j��[sr���HA�/����|��4�'��+A��!H�MA��T7��?
�B}��Ƴ�ȹ3��)A�؃��xkj�"�R��R����qC�����_�����1�4�`��||m?�R>!��'��i��� ~	"'�k�}�"gV�z���eҾ����'H�oiǲ ��\��	"�J��s�]B��d��<g�[K�S(mg�DV�"��NV�9�yZp�W����G3�#WQ\^���)��_��$6Ѯfx�@q�l?T3?�QN�`�����L�L��j�������H����k����h���|$Ï2�,d������g�y^oA��r�j�&g2[l���KL�����s��zr�Lf~�
�����y�_gx*�C�?�g��s�>�o_3� [<�a�#L�7����j-�o���LN�k6��x�]o���E�a���m}!�1�n����(=��� ����.5�4��٢,KKӫ̮־w39mY�Kl���e?0|���[��k�x&'3�����I���|6'3�u6�����**�R��L�� �i�[�"֎(-�S;��`6��3�ex=�ܾx�tG��r�gv���8Vo'J?���o�Y��/3���g2?a��L~-s�x�?��������?��ɬ����)�?��Ჳ��g�9r��l.�����e�C�e����g�ۦ�9l���S
K�mcs��h^�9ٹ�sP@Na��@��=��K)�)+��q�S�
�m�������xڃ�Z,�sG�/#��eg�,+.�;�s�M�ʙ��]�((�.,�:��xjv�6;�Pq��4�V気�RX2%���+�O�~�8�Q0�6��dz6����m�b.��AN�p�6;�V�(()R&���ܑ6�V�hT`�mΔ�{+9�6��rE%�e6Vh8���b�M��
iY��p��)�r���9� E�-c��Kf5e�7sp�#�0�n/�s���=��eS��MvoQNaaI.�()�i�;Ɩ��3Jrs�,D�Ԃ��G�4l��Exd�89�Ӳs�S��%P=��)�5�LС#ҳG�+.,��㈇�l��<VEv�t��sP��+���3�%� � :*����J�O)`ܔ���k�͡�2i64���js8
�l%�y9s��Ѷ�{�`�d��[Z8��/��t@��%��ܒ<[���Mٜ"%R��S���B���� DԘ]T^�(��-,ȝ���s������Ғ2�2�D��Ԛ� �l6w���P�Sl9y�$>P�;JJ�r�H`)���i�B� �5}
z%�� ��S���c4\Ɏ��9`��R�/����3΃8QĞc��M����l��],F$����H?�.��vp��&&�����T����!�R�˸,V�*=��V�plII��/�t"=�	���h=�p
6�Xl_�O�-?P��e%��{g��{�}���b'��2[qT;��1�0fRk��6.���k+���*e;���i%�yR�tA�DX0��n+3a�!���L|4�G��.o�y�H/K��~�F���sh?�cW� �L��l�
cK��^�5Z|p�t_ �"����b��S��ea\Qc�]Rⸯ�8�d�E`��^��`���s��J�T:Bd�:�lžqf//�n�7[���`q���}>gʃ#�p�Q�4�f/ÐM� ����SZ ��h�S��ƥ+mS@ʶ�a(�ΞRVF�# �qC2��dwK��=떐�=�7�^��85���v��k�
RƟ����q�^5�>�ۯ���������Xy���p)�-�Vq��BO�����:�$) ���iE�u�L^�ֲ닗�ԗhڋ�G+�+�jU��}�e�{��4��}
|����K�r�P�W(�a
|��K��*�~
�e>P�/T�)
|��U����N��(�z^���(�
����+�Lޠ��
ܥ�S�%�]�_W�cx�r���r4��r$�)pA����>I/��?�������
\��3��>H��)��
<I�OS���I�
|������t*x�_��'(�Z�W�/+�P�P��)��
|�_��
|��������(p�?�����+�pޠ��)p�W�C^R�
���S�s+|xo�S��x�W��T�
ܤ�G)�8�B���2^�R��
<I�+�EZxK���[)�,~������4���Kxk>[��Q�
<_�/P�V^���*��=
|�7)��
��_������x��W�ʭ�=
\y����Q��x�oP���K�wP�����u>R�s+}x��)��
<\�wV��
��7)�.
<N�+�!�x����*�$nQ�V�M�g*�{x�W�w����4���_���l���o�<��Vk��1q֪z��5L���v��I<Y��/��xO�!M4q7x��i\��z�8��	�i�z��	�i�r�	�>ҸTs��-�q�uW�U�Qmw)��G�H�dB?�4N]�LB?�4NM�$B?�4NIn3��H�T�6�!�q�q�z
�8��9Bߏ4N!�K���t8���C�nF�'� �� ���w�	����~BwD:��O�(�[�	�
黈����Hb?��H�$�Z�t+b?���nb?�� ݚ�O�H�!��8�m�����{�� }i�����nG�'�6�����^�t4���+��!��}�c���~���~B��tb?��G:��O觑�'��I�;�	�0ҝ����#ݙ�O臐�B�'����������I�#m&�z(�b?�!ݍ�O�>H�K�'t7���	��Db?����A�'t+�{�	}ҽ����#ݛ�Oh�}�����i���	}�~�~B�E�?���Ǒ@�'�wH$��$�t�����N&�z҃���^�t
���+�N%��}�ӈ��~���~B���b?��G�J�'��H��	�$�C���~�a�~Bۑ� �=�R��l����?L�k�����9ʳV�)x
bcu_k��������Jb�v�=���E�)��u 9w�~��0��"A��T����jC@5�p	Z����&�	�$.h�QK}���k�=�؝C��A!ÇP(Ͳ7�Ro�f��j�:5?>k�F��W ��Ѻ/��
@Dt������:�{�s�	� �e���(�i�'3��p�5L�Y�[����ץ�0m���2�ӐO�Oڞ���=���R��B�;R�[ȿ����d��h�wY?��a�LXF��U��� �Oyke�{�D:O9 �������
�Oڥ9 �sc}�+��ʁ\y��A(I���WT���(�sp�?��K��<�<.yl�s�1V�MqD���r^�	�/!7��w��PU�qA�V���@o�:����i.ݹ��+A�ͨN<4Z�Z��ܙ�<f�O�`����P(�S[}��U�s�q�{ zfy�ЯЪ�?�����"p[�3�2��'��G�I�.����<M*[�1�?y�K�p�<8qR�ɓ�L��.����|����s��@��H���t�^k�{oaσQ��+Ù��gVGOc|jL�1>#f�1~lL�1���l�'���Kc����$�SOt^L��cV���֤Ƙv18C���$/5&�e�q0wV�ݫmQ��;F�c��Xt|�5G86�f9��c�K�+F z�L}��W����=�W��3�����L���z�3��KL�?ӫ�i�U?�6��%��s�
�%tgK��I�k�ǎs^c��b�;�Ψ^��G����-��0k���x�=�=_Z�;i%V�O�4r��G���ǎ��v%-�W��sW��x���qcҝ�x{�֓i��?�B�~r�Sɞ�Ro-���KO��!�L���2p���%#����0?ay�I��QN����ɸ��̓j�0�����L)��8�A�d-�@c�dΈ�u�p��u�h~�7(��1'�Ҥ��o�҃�-8J]qБ2�c�+�t�3�)��9Y�L�b2�� b �p��2������L�ϴ�EYϼW��X��1v��;�j��i+�1G{%ݏ7��޸��������ZK������>��e��J=�;��V�-?��(��MB��4��I��i$_�(��K�Ϧ��[7iOPz\׸_p�x�1֤���q�j�q�V�����Se���Y�UV���4�82�9�duN�s/����o��~�X#��7j�g��=�������Q~#�&k���Ϥ�N}̿����MO��ԍ+�T�Fz�.�z�d�q+�����k�l�+Q��+D���r;���܉��Ŵ@��z�N!z�j�@��A�5�[�4�ʠ �0��74��h�A���.\��6�گ=���:�C?
7����h�iӔ`�ꈗI��ޅ�-����g��V�*�����+C-��d����@���s:-�>9�c���w�3�t���7�g�3���j�@����-x��Z}�����?����Ya!gw��)�|iF?�����߅A��S���M"�ߝ�_u��C���/��wk����h~l��F�j6/��/���9����6�*{�W�snۯ*o����?���9�2��/��I���/H��A�s���3��4�@�� ��?�w]\_�}c�����m|��M�B=�����uJ�:�o��Hb�y0��?��T����?���XY����''�������������D� ��ԟ���v��Y�;$�8bm��JϘY��{HYk���ȟ�i/�h{�i�����n/�-��Y�͟�I��C�d�䈁��I/��[�;�kAF�����U�����Zr�I�q�?^�������eW<�b�,�I:�Lj8�{A�%K?���:�R�C�2��+o��z5�B��:�Ys��Z������sM������Z�h�.ոvXxFu
���ۻ�BP7
��dm�g���(`�į�������t��c�?��'�P���u��H-^�ip���ʬP���\�M�u��H5��w��A��%p�p�x�k������j<vg9�qdݟ�AY�-�V���z{�w���C8����p��y�]���B�s�>M<��i_=�9�$����y��X,{	�G;݇qy����ؔ���9��Dv�4������V���pmRW�u�e���g�<��yeW���N��+UkZ�̿]?i�}��u;P��C�c��۲�ɿ��ߒ�_��������?����F�/˿˿��/�c/�1����~0f��ΰ��W�"SY�%q�����C����`{<n�y�\}U^�̊�{qs�:l���Mv ����'ɅH;Vz���+=���+=��������\ �n~�ִx\i.����iҷ�v�[uȃ,0EtDP�ʩ�\ug�	�.�";��
�ǰH�qr�95��dg/X}'i���Oa_wt��A!��=1�/L'O�=��7����ǧd��v�剈>x��@�C��O~F��r�����^g#jF�&st�Ծ�=b��ͳ0���Z�~U���@�C Ӷ�0 g8�w���q֚�/ #LV��1�k�"���(l�������9��w�R��"�mrt�k�=֭7Z=k��������\y]�u�
����G�?�?����{MElMm�	=u��g�E׍�l�����dT�Li�5BLr�u�q�N�Zq]m�7]GΠ�Q�:���L4V�0�D���_u�X�zҚ�@[��;#��3ͣ1��9X�ix�$�2L��t��^���/���e��Ze�>ߙxPNM�N6�M�i,V�h�Os\���x*@:o�?���b;e��p�G4�� Hj���Z{w�%2qj~�I������U@�3�|_�|�K5n1��:q2v\�΄	�U?��s�dS�ѽ�`x�/@	Y����8�k����4���_��=�qP���� ���W�qMj_��{�o`d��b|j�H����
OZ�m���Y���%'�������Ou�I^��֜��w����y�d�+�y�/Q��^~ݿ���r��	��U,ґ�#��&;�U�R�����5s�=H�\R�0�.y���3T_�����wTC�8ӧ�}�i2j���ET��Y�M�-|��Чcx�5��֩��8��@
�mW2������'� ��� z�}�#gm��f���8�JO�^�y��`G��D8S���p����s�&pS=��'�7�92��<k�6�x�h�&R��+�>zp$|�̞f\��NO� ��C���dV��w&80㲖5t�?�|�G���P��ʰE��w~e�c��pY�7� T��GM2�g\��x���qަ�8p4ZT�!�k��%e���o��k�,V:��̂S5��
sk"���t{������1���w�x�sPc&�&ƴ顈n�8w�l�S���?"�sn)�����������Dm~j�ăvl��:�Z'��R�S�W�io^�::l4[(F�Hl�
��E;�8��N�0��,�cS·��x��e��;L�ĵ��7��OwA�h�7����6��h=�4����ޢ���ehMTK�����V
$�l��v�0�3��5�$3��kP܃�ƪ��E���Z��]v�/���[l�3����|�f�,��>��B2Y�_��W%o&Ϫ�#kg�&�hKT�>�p>��J|4
��j�Ϡn6�ϓg����<�L&]g�c�oul�ńq�ń���?���S�Ľ?�z��*%�=Q�u��R������-ŋ�.��H7�L�kXVJ��y'_�K�;����^�-Uz9���s�8W��=��V�*�ib)�Sc)��!����b)��}u�U���fx(�ީ��rO��G {o7>{.�q�B�<Y�s��v@���i;��Mۨ%�S�<p�&��y�`���5?��$�w���$��s̋�%����P���D�Ȫ��K�x��s?z������x�Q���AA��'9^_�x=B#��*���R�$h��%�y+�Z����w�tc���ZĶb������^�o	=ۖ��bE�N��mowҞ�-�Kx�^�RL����4��b_�ϥ��x'_`��/J�0����5��GF����a1�2�EXw��|���2:u������:�P�w�t�
,� �o����G�����)�1���xQ~�E�����{�'��
���x-	��pj	|����i(��	'#�Hx��P��=�#�S�b���p�~��&:ҵEޑ�{!�zG��B:�_;��$o�*h����r�����&�Lë��6�buj��Z^HV�o���Z�%��=C���n�i�fEdp��@z�ι���'����/r�N��]�z�s�;�F�Rh9MW�y��u��;b0��΁�_+�R�O����~�m�ٔG���M�>�|��Um�3��Ӌ�I�͡Գ�-U9]�R��p�}�m��y�R�ӽ-5�H�9��R��iK]������tʋ��n��Nx���#-ĨҮ
���+��Ƈ���!g�d(~�o(^3��.���E�`��ow�oTs"�J� 0�����V�C��{�󺂌�zf�ǧ�L@�C��+�*ˑ|<^�MɍW1�瑜DrM@V"��Ekq$�: mHV�\$�#�r�7��@r>i�Q�fd��-��p��ު�W�-��r������J��
�_C1[�ڱ�� ���r���+qdIg��5�*������h����7���΁��c�q*��/�lD����z�\h5�l��Ϋ)�:��8,���S��">�{��}�����0���
��|�&�P���q3*�ky�Q�pk�X���;<�y�R��
�f����f���N���遈�j�LCHFLr=s_�W�.�Q�Rݝ8T�y�V�[�ƪ�d>��Ց=T�M
WZCj"�%J�!%�%Z4U��u[u(������Xn+��Ȁ��~�~u�u���	�C�.���ô�<��n-�v��#W�}_Bo���o`�%�����n~[����k֤�f�ޭܩLoK=\���ccZ�b/?h�ν�}���z���
/���|���i��I!�v^^�t�;���*GR��XGt�u�!N�N�/?���waĚ��%ݿ$x[�c	~�ܞ����1g���%ku��|y��-><C�VیW1.�Ks�f";⺟I�8���ø1�=���@6׿�"���k��%�I0��fܘ
����I&��^��Ψ%��؉E���Pwj*�j�7o�R'����?/rhB:*�M�����9n�]$�RcvD���=�=�v���?��ͳ���� �x�X��&}⃝س�d�m썟�p]kZv-{���,�)��T��<]VՓ�2MI�5��2j®'����+��%A$&b,@�ZӼ��5a�kx�Q�v��r<a�N�U���ʴf�h5��=.��*�ì�:��U�u\6����/��S�k��W~�qM�Ƹ�_�,&�4�e��W���V�0.U�1V^�Q1����[�Z�C���}ϓ�ȅ�+����,��F�j��=�5��T�~�3�U�yr*p\RŁ
�E����̡qB3j�B���d�]X�hMgRHX��?�Ѵ��P�S�3k��왹֚!p���	V�u6+>��;&$��?�cٛQ��;�i�NZ_��O��Ѷ�j����{��6����ͬSe���$y ������&U��s�r��{��ιj)}ԴC=�`�@���K�Em����k�f��D��j��?{�uMs��e�nl\�Q�J�}��ӏ���{z��ɹ�6k�nԃ&į7:���
���N�Р0���sܻ�`6��oO������F�pu&���8��O��j��^���5��.}F�!gُ���%:﷧2n�+�N3�l �!����KCGR4׏�I�q�g�� �1ӹf���5��+Tx)��@���huk;�:��*�'��Bm5��I�=�x~?�l��r=�ē{B��h%���jo%Ki%�i%��+������E�p	W�1�iKy~���8�܊�;��E����6\6���O����}��^آ�5h>�BnDN W��BZU�l�W�}x�I+(�$�Y��)�C����WI�.߂��A��~�P�.�=�� Ƴ�<�@�w��>������P�i�іz�}�~a��s�'�=���(�$��d�?�o�����d��d�*�p��V�1�Tp56P?]c��T�������1�~������m8�L_�O��8��{q@�G01���~��q�'���J�@���gC�l�w��9��oB�)��3�O�s���X����������8y$^�!�:]������{��'��uZ��fʙT����ƤYNR[�8A�.-�-׳��{��s�b	��s]���N�X ����pc��3({�~�=o�=���HaX79�Cի�Y��γ�c֚�$����j��x4>>0T�Vn��A���oY+��S����	G]����RL�'ɿ�;gܲ���|'.��C��l`K$ߺh�r��48#yW��qobA�r3�X�{.�{����au���i (��_��?��
:-�ܝ��h�v�ZyS��c|�p�e�����Hiku�ØK��^�Kd���;����we�t��U�p��*�<��+w	�7EG,���<J$���`?+�6�:�K���QyC7+�nj}Ѱ�^�U�߈\�On �Xk�z���4��iǹM\�x����1V"�lgO��+�v&��K]��*�ܛ\��� ��$��R��8�Y��y���vSˎ`�vpղ
\�ݤ���Q_�&�ߐ^q�Ļ�f�q㑦ߝ�՝�{�ͨI���ʡRM�x��6ni�2�U_��y��hX;n�A슁*��q���ҟ�T��5�������8��T1�ýG�AU����=`��=T��'����!<��^�ٴ~������jp)zȵ9r��KTU�� E�B�ƪ�,G��1ٛ_�X[n�cX�^����K���v��u'�X[ޜf��]? ��5r�F4"�슝J 4_��.ܢ5������z��f���b�e�?ء0���=��;�>O-�ZA��}�*�q��:+�Zu�b��i�������G���(�}�<�q�D��k&��O��'N"�M�����,�A�wҹ�\&��M��#�z����g�Nl���HR��4]Ht�{�j1�j*����P�uP�����hZ��=� ��ޡ'!�<O���������Gw�ɇ�s�+��&����#�\���y� ��?��5�/'�4�G3��2��.SF�߫����;i��Y<�q���ߢ�%ʿ���W���$<�_Kx���0�0�		��B��(���_y�_^�Ǖ}��h<�/�9�}�*��/d��|��D��m�}��Zz�i�V�k��n�v��ݪ܏!�+�>ᛮ�{�;��>F���x���Տx4����f�c��?C�L�*�ӈ'����x2��+q	�a� ����"�B�R��j��9n��u�y�b�7�cc����V�ac&��1�����M�bpu��m��i|'f!G�H��1�M#��� q�U������&Ńk�����ጞQfA��#�{�s��a��?��F
���� �E(����K$�x��(�N4��E�̀4�Kir�������__Z��g�#]��z���C:կUw���5y�������[<X��ӂZ�;�u����Fg\�6�e�-"�~b���S�Ė�P�!?��,Oǈ��te8��=N��y�����#A�~�>{S{�G?"��=��Y��س�ܞ�6R{<�lO�_��������&�=K�cXҋأ���o��MĞ�����}�����/���`O�;�=����o���ӊ�}{�̞{����+�$�_�o}��&�rB�=�d{^�g�FbϘ����\��G%��z�_��t�oϣ��9J�*Co�|IDGٞ���<���S�%�=S�X��s��.���6m�´��ߏ9���`OA"�geW���k+�͡��\����s=y��p/�J5#�x�Y��R��k����|E�i����J�\���q]�\�)���zޟ+�r�PԵ�����C���\_��7vE�"\)׎n�h��dF(��:�F���#C<��-��_Op��n*�k7�%�k>�/��W��W~/-���i�W���_#XO�^�����,���:��O-���	h,��_�޴��.X�^���7|�q~�b��ϴ������XV���P|�7�[<.;�8S`�f-��L&��������P����=���sd����ˍU�q�\�)�uS>�S���층L��o��#�_��Su�8����ZRI5JI�����S�S3Vk���*��#?�=�D�F^�Gf�ƴ�	�wn�9�Zs�j���6h��\D��p�Tfr��z�|Uo��<S�ż��^X;,�U ,��E2�IƪO �_��;B��>��9���������P�!%\ۡ#T%R�k;�j�NܨIA�q��1Ǳ���B��Ȉ����u_R��$] �n�?�gL�4V�r�A�圕.�!"���l�4\!��6�AK�[���T�y�Ƿ���c�+%_�㬢4pu�nW�*<ߕt�H���;�IEx�]@+�����u�iE=iE�*��D���#�$�J��^��WSd��IM)C��@��q��ă�6�bo���S7�L�m�y�7�`�z">���U�
���f�1uS��K􉢾~}�r����r]�f�W7�2M�L�Y|��{F����}*�j
��{�n�sS�p�[�B����q�]0 ��C���	l���#�p8���7w�ь��6x����W@�p�W�|��Mx5Ug����>4��W��eR�l��+x�]���&"��V�s�������u�1�?�x��*��gՕ��1n��d|{[�.��0J���	9����p��$�t�LӛO�GV�%񷦻��̱�6��$���9f݆�U(��-9��iA806L������rNf��6�$BI8n��y��ae���|Ա����I�f�ݿ�KUV�礪�j7��j���6�`���{~�ז���e��p�H���+U��+����T�%�p�ol���e����;�B��{)����R(i"��!�W�����n�]�B�|�e�oy�~P2��7��Wח�o�CG��v��(����ڻ�--���.�OZe���<�[�?���>%��	��'�tW���%(ӼT��_��{�HW|�Hב厑��mE%�9�!q���1{A�Ծ��~�^���n+��g��8E9�b���Cӡd\|:�,#=�������e whzzz
��J������z_)�"�N˱3�t�C��?���%����%@e��oa�8����0�H.Fi���[VF�8ثL|��/Z��%���9�<�Ε2��B�p������"���E6]��k�Bvפw��mycȬ{1�P�L���q>Q���^��>�s

my&G���i3���y��PH
I*$�v)&�}��@���]J���dP3�c*"�.�ׯ����>�����	"O~kO��o��+G^�ӵ�[{����=�i���h�Ɛ�S������5��|l�ibl��>���9�yrk�wØ0:ڙ�b������*'wFy���#�M���9�6{e�7>��y<I��X���Ʉc1.8� �����4�!�x����)�j*��2�A̔�^߃z�F�&�}�e9��3�[����;��	q0����뇞Ud�J!������D9���*��R���6�yˑ�d���Iּ�Ɏ�
�!��Tq�̔� �l����F��L%C�K�q�m!��v���Q$�d��5W�J�j���-��|�F�� ���P�����O�)��>�e����p�r8�M��BLR� _��nb�=��w��I1����Y�T�'QSInn������s`��qE%8gr�����>��{8��@Zy�X��%H���x�س����e����Մ������[^����,��cb�r��ZRd�[�\[�N�l�=�dqN����l*%�ʔ-`�1M)�
]���N������R���y0�D�<��&^��;W�ʂAD^d�P�W����YjΟ���RR�h�����}NJ����x��/0��(i�?��ajq	N'&�/~�4:����oC"MPn���M,�
���I�am3�l3�����^=��޹��[��/RV���,_:�^�ƍK��	ο���\l��Q�p(���L�DЯ�LO�����4�x;�->nq�E�l��?�F�	��a����Yz��.���(�k�Mu~�5�ʮ���W����ٻ�n矿�β���DS�7z������>o��X�6�̿������K�������|�����?�/��W�~%D��į��k���Z~�����������o��7�?�6��[�G�z~,��W�;���.^���a�>>��Ϸ����?�S�C��+>�?�g�������?�O��q�	^͟���y-���Y�%������K|3�2��_��U~�����K������{�oUo���T1����@Ֆ_��ίPu�רb�:��ߠ��ߨJ�w���.���Je��+
����S�P��*���j�_W���P�T���Խ�����w�q�"u_�}���(~�:�_���_���ר����w����F�T~�z(�E=��Ws�nu�_݂?����N��3�/�=�o�v��4���!�A��g�]������N�e�`��z8���'C]���.�o���Lo
*�[B��m�`~G���
7͋�+���7͋���K�w���?���
'�
��	g�˄�������[��;�U�"���b�j�}���Z�C�:a��NXa^/�2oV�7
k͛�:�fa�y���\/l1o���	;�ۅ]���Na�y���y��߼G�ԼW�̼O8`�D8d�/|e�T8l�L8b> 5~4.4�	��_��_
'�_	��_.�7��|X8k�V8g�N8o>"�d�^�h�A��|T���G�5�RM��As��Es��U�Nܦ��k���q�&Vܥi/��t�h�Ľ�xq��������_�Y�T�E�L� �tj����xH�M�Bs�������&Q�Z�C�F�S<��%~��-~��#6h��c�d�f�xB�"�Ԥ��4i�i�`�f���XE�&]<�*���k2ğ4����E�H�&S��%^ь�Go�c���Q�;�X�]q��H/�'�',��%��}�~�q��T|@�H|PX&f���V�*a��V���(�E��F���VX'�:1DX/�b��Q6���E4
��a�h��a�8X�!vv���.1U�-�+�ӄ�b/a��[�D�#��
��������q�pP(|.��I�b��8H�JL�{߈݄�b��8L�N�)����p�1]8*~�
b�pL��̈́b{��\8%F���x��c�)�[
��V�y�n�'��pAl#\�
��{��bW�h~�	��Q�U1Z�&�~�����b'�7�.�'�.v��[b�#v���W��]�~[�T��}Z���}�{�gԋ�Ϫ�h?P����#m�z�6´B�T�R��z��#���e���}�5�Z�Z�~�:��:�'��������[�ϩ�i�Wo��S�C�/�N��]�ջ�/��h_V�վ�ާ}U��������ԟj_W�}C}@��A�B���7Շ�o��Ծ��J���k�"�7��ԇ����j���iW��kW�OhW�Oj?V�ҮV�֮Q�ѮU����nm���v���v���v��'�&��f�E��%m���v���v��g�6�/��ڝ�k�]�_���׵{�7�{�o��F���}[�ž�3E��k�H��}O�f�b���Kt�D��[�����Ku�G�{#�#���e����uK�7��6�&Gm�٢��:E��Gmյ�ڦk�S��ڣ��W�����v���;�ˉ�Z�*�;ݓQGt�Q���~�u�:����..�NuM�<SW��w�s���=����Bv�y>�xHH̉����!��S!�WHL�;$4�lHd칐���!a�?�4���/�b���K!�/�p�WB6F��)���ֱWCbb��t��5�s��U�z��-����^0��ט��kM��:�{��b�޴D�����N�G���e�X�r��v+�cۭԏk�J?�����ڭ�g�[���n���v���v�w�6��7�;Fo�Ol�C�@���I�v�l�W�n������[c?կ��L�I���؃�H�����C�֦/�mL_�۶�Z����^ӷ�6���~����A�&���@���b��c��?�=��0��~U�I���Sz��i}����X�~e�[�1���u�s�����s����oAokIo�pYo2]ѷ3�����/��:\՗���/j��~P�����7�R����7�w��]��􇾕閾����~ܢ���и�%���C�q�Bߍ��#T�+4���?���B߉:�I����C;F���.�ɨ�Cߊ�=����25���\s<��D���a_jN�}�9���L�7W�a�;�[�ٰ�4�h·}��)�ͅ����a?j.�5h.��\	;��9�旰���a�4��Nk~;�����sk~;�y��KoT����A��5h�EQzϠ�t�C���A/}`��¤�#�$-3��pi�����p���p�������!�1�����"�:CKi�����p����Z�dh#m6�����&i�����%m7DK;1�NC����^�m� �1�I{��>CG�C'i���������!A:`�*4���鐡���^�KCw�+C�����􍡧t��K���[���G��0Pj0$I���q� �!E:iH�NҤӆ����e�JnC�t�0T:g&�7dH?�K���e�(�a���a��a�t�0N�f/�j�O�nȒn&HoJ�[R7��ҽ�w��w�D�"���=��e��˲D�my_�c�@�kY*��|(��|$�,�Z�KI�R�e�4ȲJJ�|,�ZVKi�5�`�Zi�e�d��I���P�i�e��a�$�l�FX�H#-�R�e�4ʲMm�.����ZvJ�,�����}�=R�e�4��O���4Ѳ_z��4����倔m9(M�|.�XIS,_H��/��;��4�Zz��7��KK�}+}��;�fG�e;��7�AZ�쨴�ُҪf��͎I����4;!�mvRZ��T�촴��iC3����[��쬴��9iK��R}�����.Hۚ]��,�����l��	���\�/�<�Ui��Tc�Uz�r]:��t��oҍfi��;��6�9��t�~������?]��}�uWx�������W�+��5U�p	�.����ܝpל�p�ȵ��]pI	�-��p�ܭ��p��{����;
���;�c��=pw �8�����	�;w�N ��mnpw�{��;p'w��	ܽ��7p������� ��I��܃�;�S�;���w:p�a���Á{p��L�ܣ�{p��q�=���,�� ���D�F|$��p$�ܓ�{�jc�-�]�V�u|o���4�~~������.�8vr�s����n����K��r=�}\/�R�!�Z8.]���t8#˄t����ʚ����܃�$��7�KS���}�c"��1	��p�=��p<�,8�<�9 }���x�rv=ޮ�������M��I������*���2��0Ka�zE���B|�o!9�ք,|o)��H�w���2^G�sO�wP�bд���w�`���~�{X�L8f�Na�T���i
�G�x���F����ERǳp�3xOÁ��ß�9ᨆ�98�	2��Z������wƿ�Gf����7���X��:�xnG8p���#9&(�mS}�����=�'=F������X����������3nW0�G���ѷ]�o�(�ٕF	�0�(�(��G/����M���ݜ=�VXj�s�-	�ms�h�3�G�K};�%��br*��_'�v���i�3�m�oRX���7e��K���Vh�r�4!`��O�l�6U^�ժ̟Bn��ɆkB���=y\qΔB����|K�6ہ‏��+�] ���O���ܦ��&���g�M�R��ۦ���&�ORh�i+4͢�ȝ����Ln��@nj䔕����g�Y p��<݄7唖ʷ���V#�~���ŠOI����ܞ^h|޿`c���W2�<�c��{;`�q�}��,���wA�m�C
2QA&�ye���}A���x��ns�ۋAP����vJ��~���E�� ?���L���g��J�nchR
4��[�7��Se��/��7��5�ߵ�+0��7�T(�����n\ݦg�������]~�����7�����O��C����X�v��m���x��x����z��0���m�������3�G/�Q����v�<�>@�������[c�D��۷������oV�6����
�-���gJI9���<�t�L��֨r�}{�B��>�Cށ��H~z���.���⪅<�����\2�NF����	��R��,?Jq��i��Ə^�^n�r
=�~�C����8��
�,g&�Ge��g��n495�\y�
y�#�oLI�́O�u��PS��%E��q����ǘ p<l���.}H �B��߭��s�������Vy<����^���)�g1�<����x"U7���BZ)�V��ZHK��x��@�/@�ʽ����[&����	 �$H/A�i�a"�b|�5��&A���)��@�� �G���e0vA�LH#Q�� �� �H@�������Լ
����� ]i)�Ik@H ]��Z�U�����ٔ�:�R�&���n=���>C@��[ ���Aj�1��Fs��ã9~v8w�V����@k8tOP[9)|�9�:KW�lշ�1��=�7�?�� m���$��C5H�|V�&�j�AR�3�T�<_L�zUj�II���R�ɜ,��LP8I��P�։�j�=�m�H��	I����G&��E�L����d)�R=D2���Rd���W�$��7&sT�g��|u�d�T#��d����An���T)\��3�����ɩA;�Q�J��XS�*�g襸dɔ,�584O�� �^x9�(�[ �!A�f��-U�T?���9nP�:L9�夅R{N��x��yC1�p��w��~E��d��ɬ�#�*%�I�4)3M�J�&g:MO�If����z�II�H���?HO �6$�a%924OI��Ho{�1m��<La��>��/��>���I5J�u��0��a�_�h��TA�zҝ���GO��Ӕ��_�K�ZQ�� �8��(o�ߣ���w+�p��_� /5�vy�E�:]2=��l>��Jq����ԓFO�ktu/e%K�s�;S�� eY��#)5�WR*�7B��D��I(��m|�]�"���O�A��}�4�'5�;A����T��ףzt+��<��y�G.��_��/��y�p�n��7{�at��1��_~A��!��0������ ���C��|�K�����z<��B���������k�#~q��_�G��O�/�eK���� E��P^����'�~���	�61�?�?����y�4,E����0���>
��*$��9o���@74B�nH(��9p���r�ίA�,�;��og_���nh�TE;[���p|��`��P}�~;X��~�o�q����eJ���ك�
�~i2�ű���ڏ!~��? M5J/�?i��d/1,���[s��o�o�O�~��A�8�����}B9R�{���������L����ߞt�B�Z�4hQ�?ԯ��������O��}�ǅ����N�0��T����w��pX��qM��T�T�f;��I��ӥRuK�L񛌹��?Y�t1������� �� �u���4<��FL`KF�?4�T�K�Ǖ[�4��ȿz�C:��*�0<�HS�����ȋ�,p��d�w\N�S1�����z���],=|�?ދ&�ǅLPH@}�<T���0Z��%F7g�7-����O�������gi>Kg�t>K_d�"��a�.�~���,��R1��-Xڞ�=X:���Y��ҙ,���Y���kX���_��4K��T�e���=K{�t0Kǳ4��3Y:��/�tKװtK�f�i�^c�؞����,����,��|��d�|����E,]��],����Yz��bV?K۳�K�t<K�Y:���Y�"K�tKw��k��f�5��q4�Xi"i� JlĦ���}����1��;JJL�z'�k*�$�;�Jl]�	=��S����9r�@��t�|6��<aZN�4.!oN1���Ns�֑�yv[adg��.�-�ܼ�򁀼��G�`���o�)�eO˳�(ʑ�c��̡��C�v�FNQA.T]� _�*qJY��[RT���aM~��C9���*o�����8��x�k�q�����z�?���g�xgn�s�qM��y�㒚��·��%N�NS��;�������o�e6���d���R��5�7�Ο�x�w���-��&�a�=�r��+J$�����a��%�øp�ؒw�(��N��B�0��A&�Z*_�������d�s�ɑ�ɬ�ì���(dxÙ�'ħ1\L�Z&_�`�g�������Lfr���ꘜ�rv1|O����z���$��AƟe k�+2��?�P��OR�0[���i����g�� ����29r�$1����s$�3ކ�2��pyx1�a.��e������J5�����U�W0\[K���$����a���w3<|���_1�c��.��'Y�����<.�1� ���&G���_`qL^���
�G(x���^E۷!����q��Ta�w�������[��8@�o�^`�,�o�z���k$kU>_)?_�O�/�|�B�1�������ar��B-�M���ʇw���5Lj��X��ٔ���R�qY>ۄ���?��>���/���:����/g�y��=�m�>S(mg�y��H�R(��xJ�{��B���a�X����H�7��Ǳ��'ӧ0���Ap�Cl�*��kr�Z���v,��3L�𱔖�o)����(�!0�����29�ky_`Z��3��UA�W������_��V��=��d�7�Ϭ ^"� 29�(��#~���W-6-�+����/A�,�=D�Ħ��G"�K�<�[���6��3Ls��`��&��
�[��i9���	Z*� g\��Z6~Y;Nf�|&�p���X��l�vg�GA�o���ԏ����~�ᙬݽ�lt�܋��=�V���w��B��:�_�t�Q�.�e"�<E�g��=�qA�ۃ�O19(���o1���GA��39�Y\��E
R�D�Z\B���N!A�c<#��/�o�uj~���z��q�R���3��u"�F�Ɛ���AV��M�+,>�"�:+�t?����C$��Yc����g��Ã��LN-3h<��M�5?���������V����~�	xT�9����0�'�8#�{o�i���oX(���0�5�+X?��94ȼ)�a����'>���,yù_��Q�_�[�S8�+,��=�<?�f粳��26}����fK" ��Ź@Y̖��z�$�-#���Ye���r�ѷ�S��,�Q�HQ��$o�%.ye[�M�R�%;+�RT1l��Y$�
�ډ��ȁg��K*\�p���	\�3PG�����L�1��֬�gzzzf�۟>k��#��L/��h�TG �p�2|k�0���E�I.5eK�\���|�@�#5(˒��۪��r!��ĭ�<D N�5������-�x�Mσ���ƚW\_��� �[D�Lγlv����-���t6]�`m�;���ﴷ;O�噶��fQV%diu^dry�\���y&��J�!9�x���������`W��v��បB�����?��qog�/5�To����cZ���ǳn��p��+�ն�淼�n�2�CÄ�Gr�^�2��x����BU=/β��r��P�ivM#͆�V���@r�v��7�ez��d�_�6���*�\�{ƭV��s
E�p�
��"a�*i�J5Ⱦjmw���#��,S�jK�n��&i|-"�|D۴�av4Y�QsOJ���F�4(�hqK�'C�jQ.v�7�h���!A2C�܃�8�E��L�K?�nL7Q���y6��bF�zf�p�&Nd��L}Ξ�T��C��p�®�b��3���!����y�����yc����6�:?]���B�Rj����҉�(<|-F�Õ
@����|x��8;� ��<�BCI�H��Tg��t�Д�㵁u G��I�M��e�}Rv��i��Ĝ�Ӣ�u����B6G�S���Bo��"[���e:�ȴ[���۳��Q��Ǯ����q�c���?��Jɘaw�Aޛ���@p��e2���j2���ڿ,Uk8�.Y=�<Z3�W�_�[�9�ʾ�2���
y�B>4�&֍q/�|����l>K��_ó�l~�ث�d*�N�M!~�~��6���Go����yl}�Q*�
����"R�":;Ug��<����c�-�:siW__��sd�.�!]�\l�YK�殩������/x������ߦ�N���s}���/Hۿ�|OyT�W���������]�;�(�J��!O�nĴ�>�eI���\�?s��ѧ�-ɮ(�CT��O���(�K�p9�4����)S>�$�@�F?6v��/IR��.�����S~��+�p����]_�>�ק�S�O�I�����'�������$?����2�ϙ>�INY����1}ʓ�����s@n��E�Oo��2���R`n��)�޽��Kc?�S~�������5x�ѧ<Wh��1�=�]߱�)������I~��m��+W41�?1}��]}�e����ٴE��3xn������5���}�g�J�������^�����2s����ex%�#�����JC��D������PK
    \O�H���pf  	3 /  org/jnativehook/lib/windows/x86/JNativeHook.dll  	3     pf      �}|SE���M!@!QZ��E��h�I���-�@��RڔVӇm�kQ�iW���ʺ�.****�E

.�[�[�]S�n������{��ܴ������?�{s�9�9s���f��zM�B��	�F�'�\�Si�з����>l�$��æ��V++�*T�)��+���ve��\YZ�̞2MYVQdO8���+#o!��~dw��H�`����y�$�z��H�	IW�z��PF����QK��R	��%ˇ�^Z	y�BT�n�TJH^l׏�
	I� w~t$]�Kq��x�j�!�P��G��8P,�����P�L�nL�b��� X�HK��*3S�W#E����D歆T6��YyTG�okDt3SJ�!�늬��_���.�H��D�s:(J����6E���($�n��� ��.�Y>�g��XB�TU���JB<M��g(!��u�����mh�NY3mQ�F��9M3 k�w�JUwЕ�'-e�ƺ���~�<���O���uUp)Z���;K�i쐿6$ʮktƙ�8�����}C����5��Ǽ�9�& V�k E6�T��
�kt�؜��*��2x,�K>�|�}��Kʰ\|�CE�����������D�,	3�c�t��+=q*��X�?�
�4<z)Qa�9a!��FYpwF9P����^���b�ѳ�i]ˁ^+ƪp�KM'��{�������z�*��r��2�cܝ��Ƀ�������7�]��ΙXa�u=��e.�ۆBW_ͷm��sȳ��O������;%���,S�<sUR$;���'����{���Nt���Pm�>���ֶY9'q��b�����٣�%L@�1�eF8�S\�(��E;�P��BZ3�,{����d��g��cPC~��w'z|s�ɿ�	�cZ�0�����P���������8o�J�{��;�]\���M��V�u��߬��5Pv���1i]�[X��:�`�Z������̳�d�2���h*��b�n�~X��z�"�\U	 �`����%p��! H��`1٪XNW �{D�!���s���������>���:	��r�8�_�T^��,��(��PȜ>x���G���AϮ��K�ݶ�p]�0y�w�@��V	L��Z�n)<�Mo�>-Ɣ�hO��&��r�f��ئcQ[����*�x�,��r$@�<�N���Awt��?�w,���]sL&��K���=��a�*���ь��%z�]X�@S�z@����R�����[yݙ(�c<�)�|��h`9�9��G���\��P�()�GQ]f�P�1T��(���Ӏ �$��Ra\sRR�nUKUS�R�e�tT�w�4"'�"sU���*��l?��xrU�(NkW
���y�B�´��eC@O�� �*v�bH��b�Z��c '�|$�C��K%�M�6��A!�^�c�~5�̊�^��:�����Xz�����Z���+���oJF�id*.^7�)�j�3pi@�L����U��ˌuև7�Sr�4���	�-�����c
M#x��d��Fw#T�l>����_^�50�i�o=X�n.e8�?�s�3�)����K�c_�~�
�g�B��xg��x�>#��w�E����]X� �m�t����;/�4��k��뼂z�;��q� ����!F(��X�|4�����������ݹ蓩�m"�=j"��4��+l"���v��4�hy�&�zڎ���X·����BwX��8`$Ӷ��߿ra���Q�F��~���~O����[,�o�������,������3ϻ��{��<%�]K����4ۙy-���2���N��=���1*2���.�j�'�Ӯk]X۶<�J"��tA��n���vb�z���~��H�:	��Y x'x	�E��o�
��o��w1���k�c������1�:5�z+TΠuk-A��B#��b��]��m-���%F^�Jۻ�Lp�
�q/Qd��5k�Xk��,�O�#�7���x\�{D��{D�8�ɴYO���+��o�)��2�e4�P<u�w��':�R5~�&�r9
5��Z�����f�D[�H+��S*���o3'��C��$s�0FP������^���JY�Sf4q����έ!��k���n*����9�?uwp�`�G�W�T�iRy��4�9Ep���������*
[NZ/:�ms
��4����g��J\P��Vj�*�8lT3�t��vӶ�l���;{(mt/���"iW\�����v��J+饴�+�v�EHm?m\�i J,��c��hE���b�M���$9����/���Fs.��{�>z6���Vn!��þ;/�)��/Q��&���Y�O�������VL/�?抪�~ٕU�����#�sl�~��_LۉSB���TIrr�D�!A�IǼ0��a�,�!�P0T�4$��}r ��~�h�6�Վ���$���ǡm����s-éR����\�`&�ӻ���v�NF�;��&AM�ДC��=��[ዪmg�}��o�T�7߆���T���vQ�g��?V��K��q�/�é���W^ �ct0R
�!i ��NW�,��=�,>,��"�2�ՠ�A�M�j:���E�v|��C�(hk����ڦ5i��)c��X�	�b.�(z�B�Ķ��q��|K�>|��纨��eL��2W�s��!�Dbm��:�\UR���ڝ����cQ��"]-�"	�x�f��[��=k�������{���	�;�,��$�7�7Ǡvp�!�4Ǡ��$�#`�Jz�H���qn����lԕ���	*h:W9;�|��|X�� �W��A�u(���m���&�B˄�.������F9<l�)���)gmxrEEH�%҂r��J=�Ju~OJ�6r9�aӁ���%����F�n��ß�z�������c�2���s=%u{g�HyvQK.�`׏p�wm�|�JY��L�*�:�皮�zU��Y�1.GIU�;���ia�`kki�1Sm0��f��3m�:Ӷ`��;0�6>��3mf�B3m�3m�:Ӧ`��4�&>�Ʈ3mfʥ�6�Vt�iE0��h�|�]g���ef��gj�:Sc0��4S#�ɽ;A�8�	��r�*[��u��0�qʻ��/���(6���TŢ�����E����������A)��2��w+�ܓ��>�^�q�!�p�W~A��Ss �s龩`-��l��N�U�qbp�q$<{!�7���6�:�F�oDvb��Q ;�B�aN� 8]x�тe��Щ1��w����j2���ŧ��Sk0s�ч��Yk�%�$\^��L��)�)�qúG�����z�"&~���\��Fy�EFׄp��w`2�+�g]��^���B�c%�!�AOW)<�2O�BK�=՗f�6���uL$�-�HЎ�H�	�%b�S
�J��[Oq�N����yNT	���+!�9��9υ�wU/��9�_
qjIXE�X5�X\E	q�"�Z���X	"�ԍ�C+���>��J_�Ȣ�Dy�[}D�-*�V�������]+	���2֓���ŵ=}b@�ÚgE:<��pճ�߿?���|�aE�4ِ�b�����jȾ������B9G�v��}���� �.��%φ�۞�|},�|� �w�D�g�
�W^_�>�^"m�%����"~j�<?I?_����h�3]8�!�ƈ$�+*iZ��Ķ�qt���@mm#��y�di$[�{^���;;Ojf
O���W^�''�����b�E����������=���p��9���ВNGƊ�bWEQ-&����Z�h����Z�&�Ev<y�T�92N�yq��%��<��T��bm^�k�y�|�G��u7����.��'�$hm�Q=mX[��+kC=m�NOm3���ֱN��S���5ǃ�/���aD�{`m�=ԏ+t���b,�Ͷ�nv��tô"�Za?O�6�7�%әA��1\?Ώ�D-뺷�0^����r^�F�a�6�1u��ZdFH���w���v�3���\���D��`zڢT�;�:�������T�1.57�Egv����b�n��9Ŷ9��Êms9��m�A�[�����&�>�����jo��b@~��9*:���AΧ�mC9�B�]��e�W������GȲ��py0ee=.F���,�%�@=J�'A͘��:j�(w�(��X��3�*����fw�E�%&P�� PV- 
i��5o��#l8�z:ΛG#o��\UD����&���:��퍆�ɥ���GL�Q���:��z�������z~X�Z�5�}��z\����Y���H%\��^pks�Y2�X4�����7P�e#�>�X6Y��[��<1�OcZ:�.�a����Q��7�(����
�x)��t2����%�ؓu-ESpO�S�� ��>��p�w����d�x��Z"�V���X��ln�QO;4���!(�{����OR��Kh+��/g꤮�JIbӤY8��$ܜ1|�B��*�fQ�m[.���+�fN��OC��z�ĸ�	���*<�թ�kF
������{8�d�ފ+�7_H/����X��ere�=���cB�2w�|X������+����
˻���k������OX��X����S�>nJ���bW)zX��y��Vq�ML������X(&��v6�Е�<f�d�G"k�8^_~́-qH�qV>��Rz���ux� �GQ��f<#g/psi�_g93�[���g

����M�2�.�8ۦ��P��'�}���n�2�� ���y��&z�R��ɥNy���8ps��-a|-{>l��k[�f˵�)�
�˪ː�S��u��^��蕣5�S}�wI܍R���Z�^m���c�	��=�|��w�A^�;t�@U��} ���Z��<@sm�q��f.|=��E��+�3>.*��ch�Ґ��Md��F�������yL���*5hoe�jc5Oʮ��~�s;흏ph+7��r��m+#�I{�]�L6�[���@)3���b�M?��?͓�r�j:���6�}��Berv�C9[F�'`�6�������P��v2 ���$�3�N����$��6.Y,�FȔ����Sht�j�4CNO_(�����=�Ҫ���)�-^���g�L�u���D2���Α5����� a��a����Z�btFS_y��%��{���\�a!�h��<V� 4y�nl�4�E|�\���,\#+̨��7�Wγ��Qa���P�����"�;���r*����і��1e~��v���EV씰bU/�K[���� ��l��I��B�ʡ�R��s�o�Y�M#[Uf`�p��Oi���
����,��/��'�!$���Dgl�"�sNl ���js�ir�㒹F[˱�ɱ�t8���������\[���RSH���ӃP�!��O��ޑX)\|�͒��%�����8�)�t��9�	%՝r}T�d���C�I���8p[��
ϰ*�=��c�(��D<�B��w'y��i
��뾇�c��_�¼�Agﵦ]����gp\w�um{��?���RS���������"/����G��]�:z([�t���S���z1L8n���f�����P/`+c���(��-Q8Q�<���^�������ڌ��}�{O�|�R���Z�K�k\�C�U!�}X�^#�E��-��$��8b�>.�
 �Pv'��k�nq��� �Id�h��N�I�n��ʔ�Ma&�,c�!R��2ʷ�T�V�
������[}bV���ٹ�m�d�{gL�|��p?��2�_T�5��S�.Ղs���0�'�Ě���:��C�@��N�!�%��K��m�y�{t�J:�?�1a	����"d�m��`{�v��뾕���)^�Le$��dt��J>�n�y����C/i�_�:\#��Ŧ��ow��&*���S��F:��u�jy��A�x#<qVb$�}�7V��M��=O�yo����Kn{�"�����y�~���,u/S�H俲ߨh#ʆ |��殝_�$-u߂�o"G�-�@��O]�����7��Iڞ�#�͒�W�/�RNI[�%Q4'N^w;���Ij�m�c��*N0Q��|h�u�ևbk�[�u�_i(k
�i���F����gAdhM��Lxt"����oe� �J�I�+\���8gB�cV�_��1
��+�)����T����ڹ8��2#Q$�[�6щ����T�EG�w��Ý��k����V0#ysW��8rص󛡒��:���z��@��<~�˱Pñp����>�뎞��7��w�����ޭ�L�^�K=���/+8����о~�8�(�:C!߲�u1[���ᬦQ��w�p���5W�&��|k\���wJ��$Q��͜�4is����@�F��S��'�
E@>χ�˿&C�si�S{%�{s;$os�N�}�;Jvjo�S�+;�WJo���������¥v����n����W��)�Η�z	��4�h��-��W����� 5$�w��؃�(Y��.��a*pw_�bOV,�$p�I���Y,�K�x��������i��Ux*�dI�;���qy|'E� ��ݘ����_m�Yd�J�χP3 U��-��U�d���F�!�oY�����~h�u~g�e�T�B�U�B�U�"+f�o��H��?
!yXy��'hǸH��9���/��[���x��Q���3��H޽���l��R0?���c��f�-xlnyb��$i��e��H��g����b��-�>'��(��
����b��W�)�2T��S��u7�uC���9FD��Ԍ-���~ױq�:�,U����#jz�ů��fPAw�h��GH �@ ��s��ӽ�8��Ó�-7���R`�#�tB�6h�m�0~ ���n�V�ɡ|���tڞ|����H��������f���p�#����m�� �(�	n���߂,���zPK��ݾhh����O�|=���,��}p`��Z�E��x,_Մ������taRz��������`נ�8���ݝ� |M�:�G�O=1{C�����7d�}p<�N�2�p��jh!�P��ҏ؞u�8�%��m�KH[̺U|&n����q0���C0\T��g�J���q�
��t��D����ŠuR�C����(qݣ8��/�}��4=�G��H�&�[l�h(z�\	H�7���~�n���#��N�k��D�N�}6t��HMՓH'��:�����Ck�x�#^��ҿ���ǵ�����6@�_Gܗ� ���D�0B��FAM�i�龇Q޷��ME+̱1|C�;8����&	�eD�\�'}q���/�7�wC^j������^j�V=|?܊��p/0}�۹L;^���ut8w���O��Q����Όf�A���Ǎ��C��ch�sh����{=L_�����G�OrY�I~���}�mY��:���b��O�I׮>^F�<�?�>Ɖ����itK`�Cp~�ZC��?N�W�����2�3!�|\43��`<>��P �	��� �c@Ip9F	���� @�0 }�%���Ӎ�DA_�������쫴}K��{T��B�K����Se�Mb�����$�;ï!mQB|Y����ʶ7C�G��
��h��.i���c{�ݫh�f����L0���\�\>>�	�-_Hߪ�A{��]�#�~�[����ˉ��[�T�)ֳ�ߗ�Lסsd���%���'�I�K�ysٮXVά�T��T���TN�U*��
ʡ��qs�Ηy�z�[���!��H��!�)��.?��+N��`�[K_��B��L.d=șd��.���N	_yRͽ�ġ��b�+O�F~���sV��!6�k��R(������l���i�l��m	ޮ�����Yz{-��#���o��k��w����SȻ5�[ョ�YW���ބ#4�5�Z1�
�uG���� _s��:��b�|�y����ʑ���!_}�9�p�]`���q�� 4��O�rg�؉X��[c�p"��. ��{C�[8Ӂy�+,�"<�X�9��g		"K��7���nN;	��:�aOy�\B7x��[F�B}�p��~��`9J��.�U'h"�C�i�n���͕G
�]Gc�dȷfϵ
�q�$ThkPhv��v��]rEҳE�dy]*T6��?���`�}v�O�=\7!��n�,K�v�A���	g?mo_��(4j���<�������qɥ�7&��Қ��.o��R�m,��/8m�47�~�
tf^A�}{6�q'�
���q�����E��ϣ��D~���H�kޭ	�?)����ߎ�\�?�c����-����������H���!b����(?����!�ڞ�l���o���;�[�T��t@�456�C��o�}�ιIU�fߡ�0*�흪a.��f'��Q?T�܏;��+�8�r?ny��ބ+z�җ�q/��q�|���M4oot1���5�P
�����t-n��ц�d]��0��G_�p����s�(�9�e��f�i�N\78z'�cd̈���l����!�����'�r�ik����Yä�o�П@�ҶG��8uD�`�Pb�
%D��&��j����wG�8C�o_�����s�kN��w"..�����.vJr�g���c`�QΙ���N��S����]2<���P?�e��gaW�o$#���aT�0F�_i��#�y�`� ?�)?ًn���[�KD���y\�VnN��=������yqBY���sϕ\���������a��Zx�V᧻�(B�p�P��'9��9�ш0R�����^�!C�X��CPs�/J8�L�_{�Y!�G]͡��P7#�_e5p�9��"��B_��p�Őݎ�}��&�x�0[���:]�N(��h'���ut�r���nז�7١F6�j�#+
O�8$��U��9�#+��(=�������hy�*���R��O���`��Xp����%w���,t���� �2����Qqs��\5���-�E�kS(MY����H�����Ŷ���?z�ً�tp� 'T�2�-�/�M�t�
6�7s۳��6�;S�Ei��s��w�U�ɪ_�U��́˥����~21<g�$���M�\�ۏm�O�%nI�앯�Zʶ�"�a��;��7N7�K8�^�dfiS�kJ���1�貢�oY�,+��=�x]Am+�e�C8������(W QF�DҷB%q	�>��I�K��֏%����%z-:(��a��I4�B���$�!�%Jz�ǒ��y��H��0�:����|��0��$26�X�}�K�˨�D��l��s�KT�!���(^"��K�?�%j�%�nua}q�{�~���z*7k��N`��P"n�'{?��&H㛡�i�[�תg3{��bFX��o�f��d;ϫ�3��1p�e{���l/b��@�o�lO�e�������g�c����͊�N�gS��5��GX�e�s�b�`_��ހ��#wn�*>�Pf�c�S�����~�#9f��e�2��3�-�"yz��s�|w��|��a�Ea�M@����ia�+���w�:C�!>�VE}������18�K�71$
H�\��)�^�����7o�����z:�y�\^6]Ԡ��T�,��|����>�ket�*��%���aq���ƽ�>݂�0��VKC��������C?t��S6\Q��]`�T�evPi�*ܴ�[��>Kĭ����kz�@\	�?��w�Cw\����_aPH99���Qw��X�Z�X�T�C�X�~k=�<��a��
W�v%��*�C�h����I�t���:�x�b�����l�P�
�G���{�Vf�w�I}��q+���B��?���NG"�]|Ո���q�dA4\��='�&��n4�3X�k��D	nj���c�����&|��w����k>Y�%q[�@�ROS��>q����	!ۏ��@���	@�F���!�m������&�+kU,��g������d��g%4Cµ�<�ĥ9q�q:��v�x����ڴ�i�߈?/�	oM�b�p�ҡ�i:5Gh��*�DO��Kb��E��w$5�di(�'%��1ҕwJ�c��0���y����u� �r��T�l�1�B����X�D�'��i�ud��ad���@kB
�� ���;Po��sTP	1��hW}�M6w�`P��c�����?����ۦ�Q��ٿ9�~A��(����H�iZo
�����N"�˖�ÿ΁t?x@���*��d�q==��D�p����6��;�Vwc&5�WV��}���/n4�쁡��_*w�G�����A\��o���;o�f�@�1z��������M��1��K��s�#��.wp�4�42�=h��x,Q�g��9�V�tU�� c��q�b�D�h)���D61�7;����{~Ӡ2� �7�d�l�u��$�0��;���3���t��pf�����D&G���R8�=��u磤�;�r�=.�T������]�n�a��y�̖m�m�9�Y��{{_c���Fwk��g��Z�a�n�z(��!k۔{�F�����UBO������Y��v���7r�-	o�%�_y������)%����W�>���D�w��I������/}���+�<������͒��bq�'����g�+����1�|�4+�}V�+������K�,ߏ?h�t�;���6�6@�=�ș�>�t���菀8�)�b�3�w���k�|˛��s�v��_,�'�m�C��F��x�z�js�F�s��?J��=���2�ڟZ�:���2u������R��t��Ĺ `h�z3�L�"��J:�yt
ۛ���f���;���X��H�p�jQc�)�m.=�ORS�6K�;@I�#�V��!�px��c�t�{�2#s��;��L�*�w���P��m���R�ڣGh'��1ܞA�\|8��4������ΐ�<Ѵ	dI/yk���Ȓ12S5�w�x:��=�B�N�EO��+�䪔��u]�y2O<>k�;&P�����~�}�g_��P��Rb89���h��U#�;���A �	�#e,�fd�9�(�����|����;���@���;��q��#��6Ǵ���(Ǘ]KXlP�D=����q;CR��<i�����f��E� �-M���j����쇧���[g�Y��`��:��k3���'�7�Q�Ƥ�����34�������e*��WN�7�}F�h� ��>D#g�Z+���ʷ�����������H0]��)0�bpj�>	zl�l��)��c��[A�A6�����xHr�М�z/�`g𑴝b!7ӸB�t��;v/�2$�Z�.�����ۇs�\�ioe=c�&�^&P�h�ޭ��T�/����~G�b�5���4�䇢�oz��CG�k�P�|�Έ����yG�N���Ea���%`���a�~(g*e׻���ÌY���T�4ry%��f�R)z奱�_w��	��wR�&�����/�~ �ه{i�ȳ�OS�$�*|(ܻ���x����	�Yw�#���@������ �ǫ��&r���]c����J������$w=�]}��(w]�]sW'��Y�]�ܵ��:�k	w-���\�:��N�y�5���p�l��]����]��U�]��k��F���k����u5w�箏�+�{s����OEї<檴�N�ui��O�Kc����jS��\p��9x��g�g\�������x��,�&L�.*�o?�>=T^� `���F{ƳgĹC_z>:���̡�~�{>¥	�q�l١o �x���E~�i:]��5}P���:�9�oӞ�i�\S��ƿ2��Ѣ_��xβ����ϻ�Ok���/�i4�+w��>{9>���sD�o�����+8=ze?�����&2�.���󿩇�3�����O4���IB��0��n����@�E�]�#��ӟ>�G�����Ԥ�9$�������N{U����ڎ'L�*ڋHQU��p%dx�r�p��fe����>ea��ܩ��bG�"e��i/tڋ�ᱢ �h��YQ��R*+��Pr�;K��I�#R�I�]� �_�'�����YXRZ�@i_h*�%�v@K	-{r���CU8���j�X�@����~0O!J�e�@�I�j�Z�P���i��E%v���$YYU�,pbѥJWy��ZY�������" �,-/�XT�,��Q����o���{VEy��5�,�+]UU�?���;J��ʪ�B����T�|�^����pJ8��
N����0*)a�%�1�|D����`a�펂��S[�\��T4fq���YZQ�8cJQfЧ����V߬�R���.
��Zp����҅v��8G��Ǵ�*�J���j2�� |zI����BJ��$�23���.��2bF@; �l�I��+��eUKR��rN)�D�c��*�P�)"�A������@F��`Z�]��L#`�*�ۤܰ���0
K1�,�;�g��IE�ť��jq��̯ٗ(�*�L�/a$����㳰(( �YEv�6�B��?-)��M��+�6+a�㹢Y��;ꩲ�Q�Y��K�9�7�`�h0�
�cT_$�>5~��b�FQ�:�^�� �R^�,-^"x6m	x]��&��0B��A\^^UE��ʹ��r"�*��]�G������ ��p�Wu[^|��)�R\Zn'���dQAU9 ��D�A6�|a����o%�.`x��g�����P�����i^zCY$eFCY%�FH
�S[��-/ͧ5��-T������J�=�`I�˙�h�:Y9�����btL���au�oG�wؕեK��V�!_Ô�1�+iO
٠���A	�e�0�� ��H�=�l��'����QT*K�Y�P �򴻦M3in�#��p�-O�;�r�sy��L��ë	�U���"���{&+�^�d��B�&�G٫��ՅU��N�ۄz[,UT��Qh�yM,D�uX����e�����@���#p�UU kЗ*y?�,+��t8mϢ�#Ա���^���JQ}qUEY���W��i�d|�̊Ezm�ACtR�l�2KP�=�_e/��3���ˀ	R0�0����<�y1H5>���^`$,=eW��;���N����m�iy��Ǎ�>iʝ��L�3&PJ����Q��cD~�����.�Os��)��fg��u 9�������_P^��MYYQ��Xo�B�^^D�ܠ�CsP�FH�e�T?��,�R%�j�������P�
i$%$2��g@�)[ ҅�U����j�&�Q�_��v8&��'��+����~D�v.?��\x����#uÈ&lAa8�ծB4�b�#�~ĸ�j��g����T;+*���F������'U��Lxz	�o�$
-z����B�J{�3�
B��O���h���*+J�A�� ��^E#��2��YZ�(��>���t��H�Wm/�.�n����CJ/�v�q�ӳ>PB~N���RI4I#R�%1D��d19�;&H�w;I$o�g~��[�d�	cȘAS��L'��.xv'$<2�,!yp��|ׁ\��N�iPj6?h,�c�82eP7h��:���I�o��Vܳ�����0h6�:h�6��� �h�}2�=	�n ��!}��jZF�ד�D	����H�V�h4��,���0��kI=F~Cn"�ͤ����)#�I���AKŠ��H) ד�DA
�`2�%�
���vHא�d$�%��{|9ޜA���A�݃T����L�"TCw���DRCr�r��a2��I�-�A-�
�|��@5G�n!(_~i����l��i�2����˙p�EX;�K�Ep#�p> ͤ��GH���t_lgy���$֦���w����ʶ��A��<F�:1��^�M)��J �!CJ������
Q����W���֍�VVfYkq���V�����u��p/.d�{V��GD�w0w�=��x�}8w�wŽ�7����ҭn ����9����拐p��H����!=�=������|J��ahB"��,)��]>�?Wy)����������W}��A��r��" ��yc�5������x����KN����$n��G��z�s6��(Q��R
�0��^��I����+j�b8
C�{�9?�$(����@�6�uys\B��'�t�&��S�,�U��0��/vB�U�t��W^��\�u��cFeE!e�(E�����Y�@��rgy�Ԃ�0�x(��R���Ǫ���a��	0��ΰŢp��9c%N ;@��"���qy4��AcAu5�F��8��ʎTV:�*���rv�Q�QQ���pUڅ��ab�,�˪�O'Ū�uAC�nH���2������A���޸L>_!�?@~eiC�(H�!u,`�F�>���WT-�8�|�<+��ٜ�ic:���e:_��,�WMT#,0Kͻ�H3����"`-d;�|�ph//u�'�0G)���yw���l�!V���9�HD�Е��Ϫ�,����}��9\���r�7�	�n���������z(�*���\�]��%Z=��R�u7rsY�¬�`�P-\�.)XH�=8v��ˊI.W��aFq5�!,���ȗa�X�rЯJ݇0�����]�0��XQ,'�g��t��J|��q(CܷO�<^I�Q\Ph�M\�� �"����dBpM�[:���
C���i���R{�\�T{�����@�gX8���.�e{0W�ML�p���:ܧ��~Cٿ5�Mf��A�3�����n�O�yv��Je	��S��,����ҵ+�rFi��U��e�Z"��^����i����R�@��ϲ��	c(*Ջ�/�;�0����*����-��P��YQX�P�	aT�@��r�/u���9.+ˬLʨ�PjSL)��JM�.YYYj�Nѧ��``���p��	�'ܮp�/|v�7��X����	n�)��͝n�T���r!� eB\W3��H�&�3��˅�p?o2!�� ��!UN#����H�/`�i-�H@�t�����t�rH� =iݗȝ�D�h"%1��Kd��O�X2�"raGNw�A�?����;���%ǣj�:U���8m���l֣�����H=X{-��x���-,	���V�D�� �A�4!W�~�\�OQG��!��!	`E�	��al��,�� ,�����i��	H�pϷ�����$$�	Bn����i�{!�@z
ҋ��B��w�d'	�R
�ѐ� 9 =x���\���"�-�ށ�R��!}	�H�!�����_�n�t��X9V�΀Ti�zH�Aj��.��!�¼��!�B��R%��!��+�vA:|�'}D҇1j�}A������6��^���".�NG3
.;��a���iϪOS������A&E���\��n�8�����o��#��/"�P��H�� �[P��f������"�ÞC�k�ᘨЍL��%ޞ4��2�}2��qCޑ'�����E�5�Ă��R�ܷD����dD4������o��"�`p\QUVP^h����_ ��i`��O
��S�t��n�$K��-���)y����*��{i���-�С!!oJ��KB$?z�r��R'y���U/ȧ_�Z���Xq�	��}�|B~'����HjT>�glt!]ԀV��F��,�. ���eƆ�2{�6�DW;���*�7���rZ�EZ0���IfJWVA�VLȓ������7�V@�A���������N6��'��$����6Z	�mT���Bȏ{s��(�x�!R�����/��M\l6�($lC�z�D�=�\+��52X�\P�<��''H�9��*-��.F�5�`s!I�gࠜ~I`��F�m�!�§DF��Q�h^A�U^=���b�GM�*(�v��\��OX��������Q�3F�OK��"|�:����1S'���J��TV�����J�v\�t�1S����?�Q��p�p㢮��~���Ql/K�t�HCY��S��_�(`�E��M�����տU�W��ޫ������1�	�Eu���A3Q3WS�Y�y\�M�K���I�y�ui#�
Ҫ��=����g��I�,���y��r��?k�׾�ݮm���~�m�~�=���ݬ�Mg��tw���ݫ[�{N�Y��n��YwX����׺]�^�O֛�����9�B�S�K�r�
}��/������z���An��0�p�a�!�`2dr��u�F�aç�(���3�MF�Qo�2N3�1:���%���Ɨ�M�������1�6^0JM�M�MFS�i�i���Tnz��+ӓ�?�֛^2�a�ez���ehjN2k���l�4�]��f������ּ���y�y�y��]����G�ߘO�,7[n�X-�,�-�X�-�,Zj-^�o-�X�����XfUZai�Z����<�lk��a]d����������9k�MfdK���mw���k��-�=j[e{ֶ����M�N[����i�I�>4�����N/N�J_��p�oҟL_��b�����w�M�>]��7C�q]Ɛ�[34ƌ�9wd��X��P�ʌ�/e��ѐ�7�o3��8�q>�Ö���U'�oTW'������4�=j�z�ڣ~R�V��z�z����3�Q�7��}4����47i��f�&W3MS�Y��{����뚷4���
��F�*KU�ޘ�J�=՜:*��T{ju������5�R�LmLݛ�~�/U����JӤ�MK\�V�������i�}�v"�L���ʵC�7kS�&m�v��H[�]�}X���/`�۴;�{��k�Ҟ�Jt2�\���n��v�Ng�e�u����Z���i�F��=������B;tQ����3����K�^��������~}�ȑ�a��.C�a��ix��1���a��y�[���}��?����׀�1�l�F�q�q���:㟍/�m1~ll5�����Qfd�ޤ4�LL�ց]n34}l��t�RfV��ۼŜb6�G�ǛK����=���4�d~��o��̟�O��Z~nn�[&XfZ�,����g�K��-oZ�e��r�r�eM���6k�u��e} l�7֭���/�m�S���6�Mg��&��mlN�/m���6��j{�v��/�l߂-��u���w�ߛ^��X�_�7�7�N�,�3�_Ƶ#3�3�e�Ϩ�X��dƆ��2d|����[�E]�>���h&kfh����|�ْz(���ө��!i��F��O[�V��1�p�ٴ�i�jm�1P���}_���]�.Ggו�<���^�m��}�K�g���K�u���������PBN�a��ï��>1�6�C�Í��㍿2�b�l��x�x��3�P��1�%JMϘ�5�2��?3����זo-�BK~��b��6�6��]�����o�X��.�����S�L���:͍��@���i_�l�4i�knIMI�H�V�M}:�K�ך�6�*�մ��u�m_���h����/����*t�u#uf��L]��R�+��9�+��u���t���u���5z�~4��{�O�׃��c��"�C�G�/�1�kh1|eh3��8Ԙ�s���x��A����Qc�`o�m>n6X�-���b9`9l��g��j��Xk��>o��r��o��6�6�Vb[o�ak��ťߞnH�Iߘ>;ckn`w�.r�R�k~zH��S�SקnLݞ�(mu�&h���~H3iӵY�;�vm�v�֫]�m��
z�3��A�T�h��ɺgtt�ݺ��c�3 �B�R�������ߧ��~�y���7�����}���b��[���X�C
�������fW�Ck���/h����kA#��N�&fP�,2������1�j����s�L'M�����i�,�#
��f����?�6�~�+�f��&����u��YK_�h�heOZ�����ZOXgB�r@�zZ���J��#�Ӡ-���-}G������~"�BzL� hI	7gܖ��0gL�(�(�X-ʓ񇌵�����~�n��@����k�OR��&�����]��G���E�I�U�]M42M<Ԇ����kլҬռ�ٮ�������~��RG��S-�٩�S禖�:S��>��$��P��R?K=�z!upڐ��4[ڴ��Ӫ�H�mڟ��H۞v�i����Mӎ�>�V7M�H�G���tJ}�>K�-v��K}��^h����?`�4$�F#��%Ƨ�o?��<�4�t���~豿7���7�2`VYn�XJ-��J�7[�Y_��a=����luЏ6��mS�g�/J�C���a#2�gܗ�8�}�2�����ՙ�u�p'��ԷjR5�R�j���ǚ��>�ɩ��������JmHݝz,�d�2햴�4uZ]����B��M�w o_�8��
��څZ7��o�k!bڦ��������V�K�)u�`�w�[�[�{V���.I�׏�����Q-��5���C�O�_�����!�p�a�a���PQ��r���1��p�0����`�u�獯ۍg��&x����Ѵ�����a�7��У�v�5[�c̓���%�e��/��[n1m`QZ��T[�<my���g�YY�*�hƃMϱz�OY�X���l�bm��g������z�9�i��l�l�ٖؖ۞�*��m����K�_��b����!^�q}�2#7��GFMF]�+�2�e|��Cۮa�tb ����W]������'�O��Q��~b�]�w���������:J�_s-�L���'h�jfk�k��Ti�j��Z��)�Q^�Q�.͗�ߤ^L��� �l�T��U���5�����a����EXD���U|�1�*�j���z��F�&�f�6K��Ѳ۲�g��#�O-�<����+�a�!<R�a�a�a�ax����iXlXf�1�V@[��ְ��a�a�a�a�a�a�a��Z�n�^��6����p��3OvZ�y1J!J�5*�q�c"�$�1	��ڨ�6e5f��G2>�h��uX�7�F"ʫ�p��@
��<z��s���b<�M���E?!$�U�"�#%l����J ��?5�v`�p�K5ɍ�����鹶6	W��k����\)x� @rIfE�s���
��}ŉ �|v�:@]"#�g6a��pą���J&A��V1-N�x����x,e$�r�}Ai9�&��:���ĳ|�xٻ��o!m��B~���s����*X�����~��[�������	��k���X�Դ�%c�)'��SPY�[�%���b"��C���@Z!9B �;�!�NH$���f%���DO	�$�0bHr ��Wc���7"�
��eԗ��Y2W��՗��uqg����J�����G�������kg.�;�
}�R�T*��U�5!�u QB� έB�{ ɻM�qB ���@��KG���aR�6~��O�ڸ�ک!|�Ċq��Y�ۆd������ά�N-�vRY� :k��{�t�iQ��4���Vh�h�뉰����C F���A�c Q�%���3CJ��q��v���	��K�A�\*C�9��Cp�Ã�Cpn`����g�2�>2 �B �c�1��%/�KGΓ����8�#-�� �!8�pQ�B� uք�܀�=@f���o�v�� $3�~��K�<e� 9+�<��,a���,J��v��>$�����#������ ���[%�^l����?�V��5s�U>�s(I$��Uf��[����[emZ%�� b�Lc��0R?�{�9(d+�ύ �'���y9B�x���@�Ȧ	!��'Bj !8 ��(�����
!�`H9� ��Y�l����9]XN&@��L�r��� ����t�uq�y�M�q)��'�m�뜷�FޓHn�o,��ml�ml#]؆���(����=�1�mwIH�҇�jL
���#�$�[�o��v�l
���C�8wDQ(ı��PTw�u��?{�@vQ]Ē��i#��"S�b��y=�I?X���.гG���j�aQ���8M���`��pI���8ri�$1��̓x�W#r�ڐ�Ե6��G�b��kI��t#��X4����G$��^B�@
Uq7RT��u�>��6@�Q�����
J����B���p���B~�[�K�.W�e�<>E��u#;��� ?�2x~�����ǃ=��G/Q���������)A�?��%V��s��툳@X_Y ɔ	=�L��!� 9"j�A^+ao��ӡ�\ڞ�$y�"���Kx��A=o�����t�_<8�Z ���E�T�tƃ�,�z��ϳ�klIx{g��!�����O#_;�'k�tլ��D���������ր��*'{vRH9�������̥�(N	Θ��<[yIZ���.AK5{��� �.pF�E��������ܒK���R��"�G��g�����'���=��يK㌒u��ԏ������2^?]��&��CԚ�Z�/�WZ�Z
�%�8e�*�ޓ�?�8r ��x����@���R�ُ��Og��l4{�V�(������!��5Vr	�ٰ�wt��{ ���2���@�d�C����1]q^Ȯ�$�L4g��uxX�zW�엡� �e��YՍ~x~�]�߈�N��ߥc�ƫ�O0&��#�'��*���%��h?����F'�t�	�]�"�<df  φ@� �(r'@:C � ɩ��ő[d5@������E��z�Ci�4Au�:M�����s���i�T^�����Ȏ�����D�1�b���s�%x�;����<C �]e�����S�")���2l��b� D����I� ��� �e���&u���BD�&��^Q�(��(�+�~��ze��oQOQ���+D����z�8u��z��^QZD=VD�<	�~\N}E���Q���w��#�^�+�Dԥ"�'EԿQ_�+ꏊ���e�1��5���BD�SD�'���*Q�Q?)�~TD����^#��!��*���*Q_&�~LD�S�E�7���bu�����EԷ���SD����a���K��Kƃ8��W�}K�9l��/���$��*	G,���gmO=�H��0)�8�m|�J�q��,k9�'\c�D��ת���p������"�%"�O�����1u��z��zmTxK	��-�)��#?bK!��-E$���gm%�tK��tk2t�u*(�	�벬%N&j)�H�!�!�	�jk��+D�������Q���z���SD�HD���^Q���W���Q���zg��KE�"�sE�Q���|�DD�DD}��z����W�ϋb�"��"�E"�^Q�Q�'��'�>YD=�W�O���Q�QOQW��z���,��EԓzE����t�l�h]D]�+�>�<�L�S�Ѻ�Wԏ��犨[E�?Q���V�u����"�9�����z���VD�AD=�Wԏ��g���EԟQ��+�Eԭ"��"����^QoQ7��'��/����u���JD�D<7�+��D��"�J���^Q�-��,��(�nP�GA~ (��?����/H]j �K��ʳ�����������rM��%Sd-�1�F"��õ��W��"�EԟQ�Q���d�"�E��Q_�+�I"��E�W���Q_�+�*�5"��"��"�zE])������"�Z�M���(��ZD}����"��zE=ND�^D�FD��ȏ5���BD�Q�e"���98|�P+�o��#�q<?��A�y��Wyֶx�wh��QQ`65������F��E������� U]�>�Q5~���}h� ψs=	��ĳ7�<�#&����T,wW;n�rZ��N���~�����N���������X#�
QTIDQ�y���W��Eԉ�:�����:��<��D�?��"�^%�sEԏ���Qw\%�D����QϻJԧ�����7����J��D���7���\%�"��DԷ���r��爨�Q�,�.�JԳE�E�7��'��zG�*��MD}���ޫD�(��YD}����W��VD}��������U"�b��J�cE�W��/Q��(2�u��z���(��o	P��pnz��������P��?�� �X� @V��Y�A�8��Ad'@�����s�dPi~��D ��.��	��
�r�}�D��9����psb�'@�.ί�R� �t�UQ� ���ǲw,pr��/�v��D�0H"�Oc����\��ӶAZ� �%�z5@6�@~?08W� /�b@�Ù�0� I���@�_i��U���TǱ�؉]�R�D_׶h]ۡǉ���d2;�'��hgw}�V"��P�\�Z�V��R	$"h}A- �}A��*!���s�?�\\.~Hv�9��~Μ��zBg�W���}�ʼ�i�M�Z栋ܣ_�<� �j��1���?@�3r_�xo���������A��vh0��PfO���~�AH��o2x���AH�����m!��C�+���c�~��e�ci:?	HW��Y@�;��2 ���o�="3�A���96��4�ɾ�$�E:���`Z�B@>(Z~h����/�yB�dR��) w
��% ���j�*lt�0�S�Hy��'i�j��8?�!�-��R䛢����Gȕ��G��Z_���s�8�� W�@�D_�ʖ�>f�H�u��W(���_OK�-@�/�.QfP#�wx��+ dn�~r;KCi�>0���F�y��k�}��;����2�s�* ���4�! ��6�z4e�k��q5�f�li_�秄ӛA��=��	�g��v$�E�Hۖzi�����Ôǌ��"w��X�XS�jg���o{��n��;�x淕	��p�>=L_��Z/��TE������c��8 5��)@��!�N���  _-��7
�$��SL�|��=+�u�$\yT��o���FZ y^��k@�3}�͋����j ��L��>/jd~�~r�k���|�1�|v�8��c�<#Z��?�#�%@���y$�O���v/& �q�� ���Z��И�ؖ��O���4�@�Œ�C�b<b�&�3���p;A�n�V))�$�yJp�'��%!�?I_C�n�g�� �;��$���(3>��N�>���3�e@�L�Q>�`�< ���g�|Q�<����k���.�Z㟏�y	�׉���_<wJ(dީ�s��(�����!gJ�m�<�ۊo�2O�y������,��Ƙ=gn{���Y"�Kc$-<�5f��1�O���d߹�2��0��ȍĶ(�riO���4��
�QA�)@���\䦘��)��y�Bz����)�AW7�9�'	�, yQ�5t�bZF��~1��O�f̧��!;��K���i������O��o�.j�<������<'fq�8�,���#��&s�l�}c;�%(�h����ޣq�*��2�������ymN��3� H$��@~ �y���#g&��y���e4�2j�OzҜ ��e>5��œ��	��N�V��c�	��"���	���&���UDD��U2�Z��z2�wޅ_����y�Ld���V�NM��brM�u����X��s^؄b�0�y�]�BX�~?aɼQ������E��v����|_u��0Ƥ����ˢ� �7Z�8H'1�äԥ�}�^�:!���TE^�% ;��5}�ʕ���������]���3����~h�j% k�ڧL�1a��Nk��&�g�:e	d0Up�x�@���j��N���t��&�y�u\�o9u�)�l�9Xq���^�X���߀�NU*`�MF�r�m��~f�	61�+�!^��ƹ�Y��+ٛ�aﶻ���������)ybI���m�VfE#�SN�~�w���2p��������QmQ��C��/��`��+�J��OYfڮ^}yۃڱ�5mqSS4a�TqJ]��

ԡ)qe�ٜ��vEř�n�R�ʚn�ٜ¢��bAY�dX��:�~��/���vК��O*�̾��K��C9�����i��d��������l/�<�9}QRa{F� �fb���&�.*&y7�P��M�i�mWl[�lƂ@�i���ޘ�7
��}P�0�5�tr�\��N{zN^ON��) ��u���Z�El��̞]]�ߛ���B��S�������]��%�[��Ƥ�W=���槧��%��5aB�VN��d���z�\��æS.g��<vm�R�[o�-MU�:��|�X
�z��V0(���	z�q�s�p�k�����U�r��Dmś^�:��､ou1�[�������IJ] [DS���zNF�,��6P7��"�{h�k�^�� ;Ȁ��R�0� w�Z��rԹr��p�1.7�L6\R;g*��h��-�R��]�U�T����4��"aiTGbM҅S�'}�G���q��I�T]��jt`F� [I��/�,� � �ko+�ϋ�,����6	p�����Qs����mul�✻��8���^�fS��#X�7ZM���Z�dP�%���k����Q�b�'�bm�W��ξ�&#'��ɽk��Ս6e8����cȖ����3�^��a�B�'3Wі(u��Fm�ܪ�pi���yuqu��2G��h�`�3��/���A,�S�ꘀ������U�P/����$���Z��wB�L� :�K��ʛJ��&^��+f�&O]���q��0��u��Ry7�v�����h��w�墰_��흾tshWA��?����Q���B�9�~�N~�c"-Z���J����|s(���^;���I}̓,�ӍEdbhͥ�\�9Nbm��`m�����3�<U�_���������!T����6���j4�n�P����;���w�H6�/b-��B���(�è�"&nN���BR0t�@b�9��mP��M�J�(찠Ð��#_`�gc��ɋ�0��1���Ո�q^Q2��$�n\�VЇ�Z���U:=�Ml������e����B5���1��0�L�)+\`3ۮ��`=��V�f�Ǜ��r�8��b��#��V:Ϻ�t�tcr�T�����a�Q\���vZ���W�����|;h�e�[�NO:�X � �l�Y}LҬk���`��%ѐ:SW�Ec�L�ugF�b2E
l�V�D����qR����i��[�(T�F)dŚ� b����p����K���q�d�Q���wiq�]��Y8b#�:��`$ꏭ�!�f�oK�-yi�Q�M�\�JD8g2�/$�m7)A�<qw;A�D�ݥH�����Ik��v[u�>T�w�6ld�����"�}B7�z��%������� �>�Q)�RL��X��I���J$����ҡ�L�؈��ϖ[�~^�Z��<N��:e2�1;����#D3s��ڨ�Y9*
�P\�M-^�0,�U�Zs����fxjؙcY�8@�6b�a���dl�w^HFT��,g�f�"�h�JxE7�"E���]Vq(�О�֘�
��i}ߏ`Ї�`6f��뗥� 񴠞Wt���?[Jy7t;�!�����<>+0"n̎(���@)�l�th8n��G�}_��嫣I��Z��2��u�1��zS�J���Cu�\��+V�$8.��Al�5�D��;qt2֔_i��,˸����`�=w��c��{m��A�^�ʆE�ٛ��o�1�H�����2������7�r965�ĥ����v]�7H��0r�Dg�弎-�6R���e������Bl*���]cb9P��c2�
ѕ9�<�+���PK
    \O�H��#�Ko  iN 2  org/jnativehook/lib/windows/x86_64/JNativeHook.dll  iN     Ko      �	xTE� \��&$�6$�ѠA!$(J�`�$p#��}1	I7�d���""�N�k�0��!���>0���
(�FԱ۠��H��T��;�������}7u�ԩS�:u�Tݺ7ٳꉆ����#�e�~i��_5\Q��"/�}k��*�[���T�*���e���
�i��dw��J�M7��*�������FN&!E����¯�Fv�MGH;��~j�����D�g)!�[iE�W3���%���8UT.BLď/���[yIU��O&d!z�,��"���Ę�"	���D����^�ú�i{%ge�*qL$'?���Q@��)#Hs�/��4&�b� l��*��U�%V2<*#�J����������ՠR[9oOu�7��
�7D�0��ZM*���9a}F�tB����>��!�n�kLL�<�gPE��^^�KkLt�R�����^�C�YK+
����)^cH��:����/Wp�45`x,������h\p���$��Q�u��/*q����Jj\{L���S�S�N���j�;q�s�;��OIn�=lX{?��!�^t�cW~�m��[�"�	R҆�RH��[;8� �H�?0���L�����-bk�`��%Bm�� �s<����~���f~UE�|�5��Έ�K�с�m��5���@�s�t䗐4k���2^�w�� �4�!ZAf��N]r��:Lp��nE��Df��� ��|->����+�wPf�v�?b������}!��]�,fW����̇�ڊ,��(�rG�{��ǎh�fG��g�%�	�o�B�9{��C��������K�9��tV��:��FVk�ơfߚ7�<�<��ߍ&h?��=lc�FWj�?��'�k��ߵ�͂��g<�J]��աZd�;��[��_|>`�]?@��6�Q��t�
����xm�]gTN��9�������b��
�e��@�Y�\g4m�q�~:�,�z�P��$g���3(�?j�TM � �.��:�j��r^a3�G�S�DK|��	�z"�`zr܍p7����m8���K?�4���^#��)����7Q�u�k>c�]�o�;v9d�:'��ze��U���-�6k�	SV���%��τ]_�T�+�i��57���UГ �SЕ�L�oWS�����h�fj���#����-�͕z�klb��#��WJ6l��aPQ17�p�e����4��x����k�}2a`�{���uݫ�cw`%q��&��1Jb��;���ZUt��O��l� ��(�xRj�9#ޤ�-��,u��렅��j7!8�̾�����ј�� ��8����ٞ�VcdH�h%���ݎZ�����UX=���0
RQ�.ͨ����u�}H��0�qj[|d& F���*+��mn�0�P���=8��[�!%���2�}>�'�}�4*�а� ($	t�JI I"AT��W��=r.����@4��j����v�Bf� �ki����E��jj���*t�Uj@�r��_=����~��R�k�U�M��O�C�V��G����ʊ��jf}�Tsb�����W��̑�~@M�����x�{�63��ȴ����tv�^&FS�B1���٢'�pC1��þ�}u?��8��ɍ�;�->�����p�aW�
�/��c����j����۰}?��ذ}B���g*����P�z7�l)9,���v}eT���0�v��bؙ�.Yo��.�'h� �}��g؞~!������ذg���F�	�-��.{k������d�8ܕ�Y���*C�È�.ۂ��T�؞!��z_윳���H��|kS=X�yǨ	�xMX�Lxﳒ	�����6Ą�&|�hoM��5̄5A&��g$N�������xmu�&|�Qf�}�PY���=p��Q����LG��SA��pV���<
=`~�6�z�������zy���p�G�~�8�#T�_��W��ѽ~�߫G�!9�܀�3Bvv�)yUg��K3��X;+���i@��5��1k(kUHlAt�j`��i>pXO:B�=����`/�믫X���뫧��*��_'�F�+rU�����Ym���ZY��6�ʻ�ޞn��,~l���8gԆ��#��Ps�wFN{|��[��Y��P�)��M8�}Y��>�Ώ��\���`*(��=�����)���Î������8�3�v�-S�d�ܭ1�gҀ,�\�f)(�5���G��kWes��ě���ϊWIS��GP]�Ѡ��P���+rӓT�{j��0������G�>��>K��-4���.� �� �5�Z|������;��=��F��⿡W�1����I^��Z6���wC��;�¶��0�����'%�Z����'�J���Ҷƾ�lk�m]Y��v�i����Pc�(?�FD�o�MM�ЌZJ��Ό����i�_w���0*�|���~,pj/��Ȧ�To�?A�%��q�Wq��v�����I,?N��0�A(X���b�:���vO�����'p���ʛ ���PN�]~���j�RT���gn�b���L���6h�
�r��Ĉ��'�AM�W�O�8�r�|�Z��:DEy�	�O|���'6��8�}"�g�Pz������k�듿�T��1�M?�f=Ua8u�����}�-�pi��m�H#���6���QyW�<��-���g����o 8z��P{3�N��[��K��zM�2$
�-�17<�b�A�--���+)���S
ܢ�(.�RI\�,6��SĶwo���luhlC��4X�;6Eb����&�(4�Z��$�����6��h?���OW�yoG����N��(�.
W0���韖w�tpic�-��w8�?v���w$���+��T�~vy'���T�%.d����}?��o֦D�{��`$��?�m�xMl�z�f(񸮧A���jѩ�#y��W�������Sw���5B>��e���Mr{��2�-
�f953ø[�q�{���I�p��?�*Y���
�`o0�^y\��xq��`(m��w�)�����z��N:��v������ߡEo):��:�P�Γ�l|G]?׏�u��â���ۑԁ������{ϴ�|�4؀���	3, �����=��-N>�l&,�?@-F�5 yfD�{�}�4#���~����bD'p��D����x`��!i3#=Y"��##� �<@�jF��c�t�Dz̏��C��-=x����_����/��7giH���2����'^���E���a���	�ƾp��^�J��3��Gzޟ������˲Gq�	������[Ƣ�hl���JeT}Y��1@��SX��I�|���$jB���t��/�2Ly��D� ,�^������Z0'��'�0ή���{����oy����������51�N�	:5�?�K7#W��h���ޠd.~�׭��Ç%e�U�*㣇�2~Yҩ25��#�u�P��
���� w)?Q[�?��h=�ҩ@�����K $F�*���+FP�
ߒn|�a�V��2��.����g�i�~LF��=p�/��8��t�?�:ӱ�{t?�V�o��j��z����8���7�p�l[�R���jXɻ����Ǜ�J�wT��:�d��ڥ�x���x�a�dؾ��*�B(��!�C�R578X8����ɒ�|F��1����&��h��g�΢,m���Y�Q^so@�$,����
8���J���jPN�Y��0�/��8��8�����e8uʯ�c��.��G��G}�9P���}��G�a�_Y���}�'���$��"�Y��N��_��/�����*���d�E���{���Z ��AT�L���� �t�0���6xz/��{/��V}Q^u����@�c{i՝���Ӫ��U�ʪ�+���Zë>���� �4ޯpJ�N	T��ۋ�]���e]U� �{�)望_�0naU`�i�ag�3�M9۴^&ԓB�p�ڿ�
��=L��gi��������Z���cU��>�c2�����:�|]�->v`������كO�8���	����w����)�'A����p߬3��	��PM���ڷMR���QY�(�y9�iP֌򌥵�x��������5>�E^��5��׈���{�á��Ut�w����ݨ`�ۿ�\#2P#��=�k�Uj �g���
�\<jw�e�G�(��w������m�8_a[��|pH���|9���;̺����4��<��j��G�˭K#ܝ{V@�K��C`ƐE�+�G}9I�V���&j��v|9���IEB���Xo�j�
>���C�,���e(��z�`>&�y���.6X�$51zT��R�q4E�|�Wkq����p��P��}���� w�,q�3�$[�h��	iC�$�f遭 ��7��?��(�����-�H��|��"�3���S�YևW�  �
c}��}�	���Ca�:�YU�0Ǖ����FöƟ�ɟ�o5�5!t�S�i���a��=N�T��Q�Y��\�0�\����SV�Ggp�V���T.H�g�Cʛ��P����!x��� Aw�:B�k}q��� ,�O��3ݺ�uX`��v��� ��k�;�/���9>����rkˡ��uY�	J������o)�,F{�<��ЇZy
Xi&��:]'&��m7N`��<Ϫ
�Q+�|s��R�aw�����4�y'υِy�52�N���]���~v
���$�٩�Sv.�=�`����N�gڻ0�kXyVH97����z{g��G4�A]=}L����`8������#�n�m*���6����	g����s��ʈ�H��˘���B�+i��!�\W��!�\a�|oegʀ�U��gB�CF_%8��Q��sY�������L�,6���KGܥһNtvG��G�%�YP��oU��1���w����|vE*���E�!�\ecX����g�J��6��O�Z�������k�vk?����S��ω����f��2e|SF˟/�B�b埅�se�c��zP�sJ����@�[�PD3	�=��%{���/}�.L�<%�1}<Y�c��P�f�����)��ud>�"�e��֣/s�F�9h�_h$�blx���{�,2zW}j!�q*w�U�wB� �{��p��Q���0H3�C��ZM6Q�l+N��r�-� 7��C!��H�dT���f����d�:��U��xK���V/�r<��(Ǘ�w�sG�=�V���Kȝ	+N̓����c@W�nQ�
/>�LnÛ��j� �id�w��D�w���/r��-��u�ߢ�V�
Р�!�w)��(q1��u7]Z�s7���)��3��ݜ�Z|_�~L���"�	�V/C��U|C(��T-�V ��ݸ��{���@_4��γ�������C�酐
��@���H�G衑\#���B�>�w#D���V��c<=����m�q�-k������c��p��-�qz���4��&�G�!bl��x=v�a�!��к�m�Њ�Ǫ) �-7�}��2k��c#w���f�oӣtR-���')�w�9K����}3����]PI���@�ʶ�FU�Cx.ϰ}bvn���Y<
h���ѭ�ˡU7���v� -��	y�Q�z���s�e%5:�7��9���k�F�����뗀���\���t�'��w!7��^4����VK�����q�����]��:����7���8�VI�����UHw/)I���Kؾ^1���x�<���K	�E���F<�
��%ބ;	���ܑ���j���Ɍ�L����S�=0�D�G����Ѻ�Iha�	��w���R[���g[�	����r�ɇ�Xܭ����FǍ@��V�X[�Yor�)����.�;=�kϨٷ�.�d�Cji�u�BS����m�����{�|U�(ߐ�(	[m�|#k�|��S�v����#K�}���{r~��e��
/�
���V>zT�L臛I��X5v#;�e�]�oޓ��U����s��~�{$��ذ�UK��Pb��]x�5�1*}�b�	���_��M�|�o�D��1xk����s�����/^�N�������k�3v��n���mE1��4�׷}�o �m�g���m�(򪶵�x(*�[��?߇�֛#˯��&��>�C��kT������y��E�7z�*�*o} �w�t1+�Ln ��mbp��	��lNw�
,���{M�?! �_+��&<�z��e��E�j�d�΢c\�u��Ӡ�N�R�Q/m=��n�ƺ�UVis�O���_Gb~(��_IbJ(	�$a%qn˯#qI(	<�4�딄b��{�y��g��z���w�����U�3��@Fh��!u�'��)swG�gTx��f�]�BV��R�r���L_ޥ�\�9���C��K�C�]$�;_:���.���멨���Ho�xL:���;T�b�^#�7?�//9׺3I*:'�H�>No�CQ�Fz�"���M�v?�n������'��"��:fj�tx3�P3���H�2�L-�L>��C%���z�Y̎67gҗ� 3�hXu� Z�a�1����N�g=,g����-�fk�l�%��r���b'3��.���)_��є�Lq*eK`k����4}=2f��_ �FPB��@�R.��������?�Jǝ�i+�فk+��`�ވ�8sÿ	}�j����O{~�<�C�p'v�(w�AQʓ/,��^��'߱�]P�"z}��k�J-�e�縳����LKߍ:�<Q|e�C�Z�W9��� ��m��/����#>�� J����X����#:=3�R��
�(x�߁H���D�a��NK�V�$𮥒�8��hbO��̓�{�R��`�r�UYF���s�r���}b:D�5�&���&�+a����?_z���Yi>S�T2����������^@jZ�t�|o1v{�������c:]�D>}Z�y��T6b�a�@ST����nX����KiQ� s��m,L4;d<[�4sÕ�9���2C���A���̯p<� ��o����5�[x��J��r�>�ր|�g�|�p�� ��"�?�/I@5�|��X�RQ���g�#k��N�~��v������S�D�5-�9+�(��hy�Y���!R{&lo)�	�G���N-���)��3Jz,�U���ƪW3z{szZ��{�OOK�՟����(x	6S����=�v+�J�,07�-�qqta��J�%6{�����4��ɏ��F����>\�V��\0����ɤ\��M��W�M� �:zF:�@&����P/�_�^��"�}2窦����h�謹ថ����3��fD��lTp�/nf�g�rGI���s��
�$9JGJp#�x�M��8y�p^l��G�$�����a�ͧ�g�\Sw2���(�^�F�\�c��?�$�9E�;7)dWp�v�>$��PˊM�2')j���HnL>̺V��۞��9���L>��p��*޾��yl=&��. ���I����!��#�-�@5���_
���#[���-������[��>�_0�y�92�Z����?_��gV_�|���F�P����~�Q��:jG���M�Нe<�%q�v�V�gS�/͖����

v���ŧ�a~#���e�_G�)���+i�����
��.F >���� ����lxf�a���/�{�f�����{�O��ϗ������K��/��N�F5�/Xqr=u���0�\�n���m�k��}��D|��?��J��T+�a��� ��|�1{�_� �.��= +6C*���S���D(���<�M�gX�$4�r�PsF��aa�6��,�x��5�Q����(�'C�: ׍�%O�:��t�"~{�r���m�}5�-)CM	F����o�f�fnhaM~��4ij���o�����	x�"�{��*xp�Ϫ��ALm��7�6���,�,qoۍ���rk�����嬝lGh'	�q��g��4�`�;����J�{)�R�
7���c���Hs���b7�{��Bݫ�լ����Eݎ1���#!����wZh��՜�Y����v���N����>ZU���vg�4-v�/v(�GC(������3W�jF35߂D�*rǐNyF#w L`��1�Z�����쑰���ć�"�	+A��b�u�h+�zj�4҈�P�ZR,O�k��hA̅�-�r�\�6�'��0�d���Nt�)�,1/�P�!���
����j��@:�"~�JG(!zJ�+��PS,���G~�����&�m���SXD�x�
�^�
x�_0@63���p��p������m�8�3���� Ρ1(�DX�>���h����ty��ā���O�R8Y����͌�BJ� {�:*���	������Y$1E������-�#���c���G��{<�Sz���Ь��0a^^�ֳ�* |�٠�����&�{4RL��s���UK��+�	;ƹuc��a�tfƘ~�<��}|4]ҏ���#�=��(X1�Vֲ���V�w2T[�����>6�j�;�0��8�юq5�|��Y詪��̶��g��ݟ�����=D�	��_���~�g�i:i���U�-�U��Q���=����>����0�}f�mA|����~O�Nt��ӯ�H�R��0l�Rv;
 �a�:"�Y{��f���.QuB�����a3��P���5�����<�S�A�k�㶝�FFnPn5��g6%�S���������^g��u@f!�q��P����d�N�557�C �e&K�}�#q��k0�G�HW��"�k8�����I�k��5o Gc�3Լ�i4=��a����8��kf�ϰ�?�ѷάɬ�ڐ�?ð�(����a�SPr��s��?�0���.휸{�W���c�?ԑ�k�"T�]X��"�eu�yl}�ڍ�L�tJfʷ�g�|���9���a���N�Psܺ�*K���;`q�┪f��]q��;��ǳ'f��(��&c&:�B�k�����g���4�)P�o����&�;��R�V�-%�8���1�Rti�q~�2i�.N9gu�`˰=�l�8�D>'��� �!�y��k��\�uNeX��U�a��;(M`5C���أ��cW�ެ���He���j���It@��U�~ 1S��no�����TjT�D+�G9����v�Ry��,5���K1��W�oX��Bק˅:]�,�Ն�k�~�T�+��K��ܸ�n-�����D������ؙ��C-3��8C���(>(�]�2�)$��AC%���c|�U��<M7�WÔ0��t�kV�(�TD�˯���ǈ-�OMA�m9}�������I�)���3�~~����H?#�Z��)���
���M�p�}�4�[~\;���hC�YC��;��;�[y�y��P}^M�b��W�;|d/�����IMC�Wq���߹�;�	�Y.r�V9#1��Fp�'���R�G����\������=�9�/����r���e�{�O�^"�O��-���ov��.v�_�Pw���SVY�)z�����sjA�k��O�-��uNc����xN���_�me���W�_�r��?ڰ�'��t 2fYT�_��%p;�W��k�0�h{�c��M�b�R�z����7.�{���:�?A1��s�P������C�>Ȉ�D��x4#���G2ܺ=#p�M�O����}�$�æ��J��E.ΧFT0�=.%���r�?0��$��:���,�]��塇n�W�?�~�
�k��ҝ�YCq���.� ��O���Y�2�4��u��?ғ)k��IV5KaU{e=� ���b+}v�%z�.�3~M!���WJ�<󄟕��fR,ɣR��D��Rd��R�f*�ƥث���)���R|~Z��.���[��N����_�f(�����^�ٽ����?�b�)I��h\��\*ţ�H��/E���ӕR<�=��F���H�Ƽ�T��I�iL�+��H�_���P)b��8��b�Z���)����~���M�}�s�ѳC���b(�b�4��\�H���N��M�)���R�K�g��2�A����F�A�2F�Ir�*M�|V���xFc���Jj��#Y��ӕ5����Xc�OR�tFjX�e�uX�(O���3�ơY��3�5��-�XcÏR���[E>�j��d��D�+^u
O�I�
<ߩ�,a���j�"��
�������?o�V����������/�\����C����`&����S!������i�xï��/C��g�K���9~6��}�����?��&�J���р�;�i��D�m��q�N�N�:c�=1�d{n	���ȣ�ya�U��m1�
������D�ѹ�վ� ����n���	�2d]�:���~���ʦz�?�3=o�ԁ������3�#|�B"؟����8Q�˧��K �,�°���7/�ESg������a��/��ZR �R��Qs��\G�V"i�}A��]��;JM�Ai�ݞ�x�
n^�Ͼ0`I}�#��w����&y���9��n?�I�=�ÆG�\(v捿�(�/�Ŏۂ��v7V|bf`��v������%�'7�;���y��|���s���'�W���/�⯙.-Ω��~r*���S\��6�ݞ$<7�VC>p��x>�B��6g��˖Y��c�a�`$ðiw�Hö&W����R���d``�[[mnVѓ���R��j�Y4�\��,W����Y���_�K%@���>Bi���6���,�`��%��q�<=� ���K0��VKoMx��8+8��y0��&u泮�>�ՙ�p�J�L)�p�+�t�mo o��S/fb�7vf^b��5�������w/h\l��4��߂�0�,�C#y���[����>��L����{!/7���Ǩ���4��S2�����;�+��^a�w}��!}��o��׎���[@�1Z���}���$
�睠�J�9����_N���/��g�ҝ��ֿ�q����z`�EŖ�`��F;4b��!�.>`Îoy��@ga�f�0�\�,�enS�x���.�	�>�(��N���.�g���iXu+��i���Oev��y�.�k:'���������}�c���m�S:���S��}F��>��!�{�=�꣕V�Y��֗�*�ѽ�(��@7c;�bn�f�}�Ҿ��+=�3�X��L'q*.~����9��}D�è��K{�,=��y������J�\R���rh	��R΄��R;���4G�H�6\�4�U��/u�ry4t\{/��Y��\�]�$�VN��ԭ��ؤ�8�h�q��:�4%��B#�O�:��)c�G�LA�5����&�9����a,1��T�����}�~v1��jF�K|#�f/R?E��N�{��)77���53���w��gjus��|�{�	��v��d$�vMR?���18~�e�>� �.�"���j�mk��脳��]tΛ���k�B��{'��w��G�+�!�����9��&����q����H<؂��4�a��/�ƻwl�d��z��:��g���b�7Sa��A��=CXz����7���O��'�B��)�y�~�����o�e�)c[eZ�g2�|mdb���ȝ��J�a��b;�|R�X#�L���H�[��eH�,zֵ|b���q��3Ń����$��XQ����"|-�K�=������?#����@�����rU�k�h�š���]{��W<�;����=�z��/�'̾ջn]�u���h֭�����m��~���$;���#6~2���Y�K\HirD?�X�6�Pg�ϗ7��*��o7B���i�/�<�R�_�����V�<J���;���n���H� �\#5�rL0d�����[�n������48AW'+�m���}#u /�ңTB��ch��6R��w9F	u�����W��{�1<#�<��y�nQ��h�C��;3ؘN?�	KV�I�~�.�wOq$~G�Yw�HH_-il�]+2�j
}�L7�R�e���v��M�[�|�f���>�8�O�}�������Ip?X�:�q�<e��������v�R;鿙�����Wy�@��˅���14��&)�;��S�5c���M�%���ƀ���&��<6�FO/��d��̧�
LagFy���"~6	��|Ϻv�s����<z�懞� �Y�e��������=�~j@�.�%�GW�1#�i��[�R�����=Y/��R�7�<�.ec\�1|�u�/�V�N�U�l�_y�šSx\Xp<.K��E3l���L���w���������H�Z�� =��H�K����J�y�����롙A���qz�Apd nF]�Y׉3�4�'�պLS3г�ՕF'&��:�,4��h��}�1�L�$<��Y�|��V�����~�Y:%H���TT�tn�nK<���%8�j��K��d53S�w�5���8P�%����SNgț&�a��ɐ=`㫩>�1i�����vax9���ގ�����]�Fg�k�<�k�*�G��>��0;Fu˶��\c��{�֭a��Md�1��5*1s�������5WS���l���B�ʬi\�'k�~��Ѫ��5�E����a4�4Ҹ
��CD�?�Y�@m�!������էP-���hTq<M~���hΤ�.�O�G���<p�L�~ �ڞwu�W�:ҜW���>��-��Ԋ�Pt�d,q�(|<�g��xǢ��qP��2�3��^�P�/�hn�:O{>�(�{���qɣ����Q�e[�J�g�Nw>���I�[]�~�8�`��!���D]��{t�D�����Ӎ7�#G�`�[2��8��w�V3��}muV��ܠ酿��V�����E�S� 1��U�T��ѱlQ�T<��p��0o�v`�@�_�zb�����zfj�/�:�!-�ϔ�"���a��c2��I>܀��������9�nt2�w}Нxq#ħ0�p��ɶeP�>Py���*�ҽ�(��ؤ��U�a�6u�OP�J�.f���J ����9��'_D�0F��th��g��7pd�;�s?W=�K|�N�[���v+c�����r܄�y��g�����j�~ӓ�ސOs�G]s��SA?	�'�?+�G����G���s�OG	8����7C����v�D�`s����a�Gp5����bn��:gr�k�ᡂ�,��|]d��G>DU8���:i�:ϭ6����`�&���	&g�O�*C͍���(��s�yG�CͥP��|j?�<4����o�6��6��˼���f������h�(©)9�/J��|3����M�9��d�V����U��%�Y+a��� ��Gt�:�m�!&4M�wa��<f5�a�mW���gV�`]f`�h��\��<"l��G�B�7������@49�����h�� �v��O��3����=��vc����k�@������{���iG�wv�n����h�b��]�?Lq4��]���J�髸����>M�t�/�����ehDM��u�����v���H�DV�(z��5��R>t�y9Rp��0m�Ba�ݷ@&��������/�����)���VY�8�D؇A�X�q��ER&�x]d8�dZ���<춹u_��|�<K0���o�3�ܿ����e��s]�|��5�zK�u�V�)�Y�8����= dnݟ%��� ANn��Hɞn��1��Њ�y�~_�O+�&��<#f�.�vsLTYa0���2S�W̀aoI9l��A/��a�g��:�>��P:@����� �!���{���o?ر~Q.�i������v�M��w	�9�Z�a{N�a{1�=���M�@6���H��j*g�o8���O�5���'ܑf���bm����@D�!;Z%=$7�����>G��+�``ʰ=CFCk�;�	@w�"s���߼���m�>��	5��K>��FՀ�Ү49�h�,�vS��+��ˑ�$�ȇa26d�F#Mz"D���������I<ϵx� ��g����n�幔��&t�;�e$��/�!�F�2��'�J��1����3B}��o��?&�����{ 9�]wh1��#�8bk}��f��Ed������\�c�>��ɢ���)#�[r�T����X��_ ��Ҝ�/��;Z��Ka�.Θ`P�����Y�o�A�o�Z���SO��t<Oyz	O�xz�>�~�ӏy�6O_���<}��O�����tM��~����Ⳝ���tO��7񻖧w��>%���ܝ\��yj��4����u<���x�ӟֱ�_<=��}<���'yz?OW�t!Om<����<���W�t�:�|��,�I����������lOe�WUK�?B~~���ՠ��Z	֯:_ڜ�~o�5���G�o��U,��"{����2��4{�s���Ғ���
g��8v[i�"S��a-tX��K����GE�i��d��[���Ex�()�&TI4%v����z%U������&�B+��XRi��pޤ
SG5���+ ����J'|ح�ւ^��W��wY�_!��Y|V�&V�/*�ZK%������.19�KU����������E��<����bQ���R�:��4���J��*ʫ�e�EG��T��Q��/-a"W�+
�w��Qq�xW�!�\�aH9e&�Y���,���+*�Q�򰂬�����K��O/-���T�&X����Z�(�(�����n@����S�T;��:7��H"I�H�}����%����	��
Js�V+o��J�$
 >��n-(M����~BV'�����D�G�F$��� ��ƙd����ZVa_�(���N�Ͷl
δ�+�?F�H�4 }B�%@$�a�AfƔ�I����{�K�t�v��KP��κ)&�"󭎬��]QTb+�ګ:����d^E���74Ѻ�5� ���ґpzE���ZP?T�!�Riq��S���8q:4��8y���z�tt~���f���t4y%q�<OEi��L"��S�9`�V��E�����炌�Hy��ĶDV����a-c�ҥ�tr(��ͱWTZ�%]��V!���-w:JJ��V̟�-�Z����4�W��4b+)���r[YT`/ ���5�����I�&0�/x��o����3���,\�������o\�S
W�:e�r[yI�]i޲�Iw���y.��p �r�N*��ty%���j"��D���Z�H��c骬�ZZ�$ o �����a�'´`���X�,u�T��p=�� 'YU\QZ�5�*kyU	@Kдd�lNb-�I:�С��z'����$�{=�?$<��UZ8$��ri"��<-���ZY��������c�ԇ�h�1�
�jL��1�����!rYP^��܄}b�bESE!�(QV|C�iFr2�N��D����y�Vټ-5�ۡ���rH�v�ݚ���^�i�\VV�S,9��:���݄�o)�Դ��0��`|N����d��LP�Eօ% N��C$��TV�J�YYaw��U�ٝ��OE����i/���]Px����*W��*���܎�'7����b�N�\c��5�R������������p5�ua�w�^�	FSy2G�'��*+�,>Dy����'��X������A�!�:�$g�U���/h�Dq-K*��nB�PӤ���g�q�RJ�B�+��AU������ed2e.��+F�
�k��A��'ʨk(�V)�S4��%����L%��y�4�ʝ�;%3{N:��dc�\9��Α�41)���"��4�4��\E襙�t\C��Ց���PYV{����^R騰w�W��
�EE�{	�I6�Ph�A!��gQ^�B@Y�1(\1�8Kav� �K&���J���>(��~�7�O��
Qt��^Q�����~���n�a ����+�\�͔�q��?�'�@n>�y�
Q�j��ς� �eT8���%Ô�2���,^��ʛ�9%�橹��9���V�I\ Ǜ�4W��<���]�O̜9�f�䌌L�y& ����'�\*��� T�+p:*�X�G��n�e���y�`1/(����}��`�3|y�)/�M��03���b��Ë��$���!�-����H�_G����@��Z
\x��5r1yR|V֗\En!�t��$�Q��d
�$�֜
~�f���@z��'�x���;��$+j<�%j�9J �n"['��B�[w��֏��p}D���E&G� �Q�͎i��O����W���I�I��ǁ�ۀ��$�� ����v.�q6s�K�B�lI$�s	�&�d����'��br>)!�&E�
b-�@[H) �y�H
I�O.%�|�{8\�;�0�����P�fG�I�D-������Z	�L5D��n!��DRM,dH��L ."��b-��*�����j���Q����a�T�p��0M����G��2����@��C>!�'N�hYh6�������6�tc3�/�����kkP~���*�X�v���@�gy����6�M	\��*��
��p��Jl}�$AzA�߉���-�VF��������V��v%a��oc��>�S~��ϻ_� ���+y�_�³��5�apI�j�A�W��/ⵖ��.0���{�������C7O�mp�W����_'Ӑ�&�"k8?gy	�*�Bx�W��jy���Jpt�@��I���3Qz*�����x��Kǝ0�S���bl�R�Z���6���尰p��!�b�*XVEwv���sA���!q8��/a�����A�Ov��K�(�B�`��z�8Ӄ�;�������f_��yu���)P]��_���YG�2 �B-�z�����_=�H~�Ȅ�ۻ|�R�y����CG�o�[��®��2H�^�3��K���C���?�o��s�����4)�D�b+(�JJ��Β
J����)�\�d)�g/�/��P���$Pb��a�����v�%-m��i�m��ͳ.�_B��{XX���f����;kg�;
ΪN�͚_^�}d�}�����u����>��1�3>��ϗ���;�z����i��+H_�k3\�õ��p�k\��z
�J���
�sV9𵨠���a!l��ĔQZ�]PR�0$t��������r+��� �ZV�7�?���t�o�Qd.:)d+����r�樨�SvM���VC�o��q¢c�o!���f�U�~d靷+ϯdC�/��kq+��Z�i��N���ip�����TRV0�:��ZH�љL�J�gA�-N�}�|cgp���J����*��R�E%�bƆ��Ńa�Ͷ�+���".J��N(�QQXQj�����(���JlW�b&V8
���+��t�'�@���Fe~���sC��{��P�3��_|N����勃�Ĥ�����|\{�|�������|N?9A�Ay�����oҏ�Ǡ�JW��^T����������� ~����A�Ayc��A�MHO���0�vE���Ĕ�kL�ɉICM�%�aI��%���������������� ~󡕥�h�ZYݟ��[Y:���8?��Մ\�-��8��!�O$d
�'A*���9����� [ m��x���6��z������C:���k=���7��<܊�0!������\[��Wo$�e��i��{�fB�D8�>��a�q�\W+�@�;"�ҵ7A;p_�l�ç�?�ኃ�H�n�zpo�t\	p������=�B���C�7�r�~+��Sa~ĺ�N���C�y� q m�kͧ,=�=Hs&!�ઇ�4H�k=�o�4a���5p=���~�V��o�e@p�2��j��� Hޏ��2�cp�'�
W�,}����p�)~��,�@�$\���G6B"�����+�O���&���tN9���C�� �N��"���p��ˀk�	��ל,�W1����'X:�v��&�p�s����u�	��k���pm>�R\O�};�7tX.o9��{`���	���~���e�y��C㿝f�_a��� �������z����.����R'p_�Kp�����K�	�����Õ�K�������ߺ�|��ip������*����]��	���Z���.��N��������������?�NMt#TI��>$b�>�O~X�.Gۨn���0>",I�����UZ���Qz�.<�o���ONX��Eݪ
Ӑ�q�$U>��ђ>�5I�|U%�~V���8m�&_]�ʁ��/1��H�^�7G�֢mU���/��<�iJ�y</��d��� ��Iplww'�"e�I4����᤿��S�Ki��?���n��$]�&�E_�㲯�#O+e<�,�7����A}�tNt"�ċ���N8��e<��t��4�Ŝn��uc綺1�Vc��1���ڨiQ�(��G^l�#d:�ۀ�Gg};B&Wy9m�\�ӿ�¯�O�����c�W��z
.��1�x� ��0�����?0���~���Ct�����j�+I�"p=׫p����*b��V���Z�Z�6����DC�DG�H�'}I8�G"H$�"��vb7M�ʻ�o�۩�4��y�����������x�o��N���������MקXz}ަ�k�=P�{��r��.��+�@Ů����Wdx��TdK����`�U�M���mؖ�*rV�^�"1�{�8\���X%�<?���xZ���<]���<}���y�!O�y>����:�N��<]�ӵ<���Wy���ox�O��giO������M��"��yZ��{xzO��S<����y���-<=��V�~��xz���8%_1<���4�N�i1O���}<���m<}�������XzO��T��,���tO���-(��Î��#���v���l��^ZQ���|��\i-�w�I���i�N+� zɀ��aM���Vs5�A2q��r�x�̥�o�&X�Dz;�O��e��2( H�j�Z
��-�x�gW9K�}NS+��U�C�����(�U6W�w�#O`��k��:��*(-�#D���`a�L�`����^�PE�X�
{YAy����B���(^�;�i�)4<R#4����[�ً9�/�,8+%dP:�W0b	�:��C,�͵:�g�＂���mn��ZIvh��G�+IBvi��V�
h����]!'��Ǹ0���'����QhE�uq	�*��WR1/�샗 yeU��h�P�����zR��c��`u��G��,��O�y��+�cA4�\S0��� ��B��!�h�5�J���l�����i�8�iM��b+Bh�J��q�Dm��^^XVI&i�$ꄘA�A9�7�&� �����v�`6h�`>���h�ZR^����q�*��<!!t|��:ߎ��A��b/%��CT!�(��Ba���:>��y2c���"�d[��B��Z�1��KbP�@��9ǫ��BH�:��yH|4�L�Q�Fs
��tzUV���L^QO��W����<!�����D�� �݅�����9Y׌�� �� �뚘9yR�%�v�~���ja��������}M�͜����;���t~&��������%��0i<���E��������ȯ����7�mH�@�B���n�lh�@67�6&mLۘ�1c����7lܺ�qc��֍��&�&Ӧ�Mi�r6�o��T��~ӆM[75nj�Ժ�}�l�lڜ�9ms���͕x@Ϥ��ak���$�7B��	�g����_�_ze�W��2_S-̄��J<-OU�D4*��� �����Q�|w[�.����~a[v/	#�&!p��@��Æp���˻��W{t����~嶥�7�i=�\��������w�{�eP�F��� i�F�D��b?ř�	���~���j�CB~�����i���8��t��P��U-���)#B����};�K�m@��K�_��ٸ�g�_R�~�5�~:��W��`X8�[{��l?�c�D���V�cxϪ$���hk���cqo�����
�H����7~�r-�:��IQ�
5���CF$�:��&��qQ�f�)@��XKو����yn*����!��RF����o���Cq�B��U�f�8gl�ń��#�q~��?���^X&z��,�$p�rQ���C��/�CaR86(L��a(���(��`�?Cae8�������$]"�� $G)H��Dȕr���9�oؖ�v�9�@�{�WR��Q�zk]MH��~�(@�d� .�[�@$�����3�M���8|4�KcY����yG�qpϣ���(�fۇu?
��@�����l�
8��ZN��p9��_�����C�{ǔ$��:��C�� �1Y^+ Ցr�:;|��v���Z��\#�<
�V���~>��Z� �
�/ ��A��p��4� 9�r� i�C�q���p!��׌�	�8|\���l\T��Tpظ���+q��ȗF���0��A��EZ/��'��q��o�~��$I8���8_�?�a_TDZ=�4 ��!��$) � ٪�L�1S)���9y����q$ߏSd-(�>c����+�%�k=�Vd7�%�|�������4����h9�� ٠�� �
�I I�I�� �
�U}�9� �� �W�l��8o $͏��t$9�G
���E,��BG
FKJ��FJ���Q$�'���4R6���2J%��F��%��EI� 5�ÑRً���~�|�����H9���6�3B��}����\ �ց�� [8� 1^"ǹ �S�8s�r��q��k���+V&;�����,2�0�6�HW��H$�HY�J}�(�\ռ�n?�����⷟��`��������R۽m���%i��h�J��� $���jCۘ&��Sx�~�)(�H�ty��Ҩ��~�t��r���pj�r b�!�qb[��(�1�٢g_�i�[T�����U[�4vT��K2nQ�Eu⵸E����'A�j�Ƣ���'�������f�]�`Ϧ�y�>�Q�Z�E�(��B�&]�;'��2�3��p�U�5�>!d8S�����X3hÔ׵�*��2⺀\���ȓ�sZo7Z��+É�ܣ����iïg��Y"W��Cw�B������;Y�q=���#�Щ��ԍ����/W�_�4�\A8�*�������c"$~�)WN~�H)=�}g�;�X���� i
O{7B��G �j�<d�����~�sH�c�ߺj�.��F��6L�t�ml�fJ�/�J�ŕ?����싂�c�]�sg�\�-�F�����
؞�f�;�_��
B�a�?�%LS2�E_�~R_t��x_�Ӌq���q��>yJ�K�(��N;�IO���i��s��d��Q�!�ᘅ�p����p���c�/�<�J�-�9����g͢t»�1�ͤ��=7�����{c?�~�̧T��Y�����'���=N�,S�8fc78�C���0޿���ӵ�D�yȨh��V��=7�Ge'm�Q��E�b��{m�I�{�~��e����(��UY����Q���d �B�ϼ &NBzx.�(�$��sp�����{�<mWO0{Ӄ������$����80Ǳ^N
ő�rjz��rz�e/��h���!��W��"(�+ �r��(p� dHq�.�M��݀v�R�_]�5��哬��Z�dϓk5���g"��Tc���4���P����c�\�+p	���9_��w� D���	���q>�'���y��B�rMt��V�s_��ק[�ѳ�g����:񽒍E��
h����'��y??��ď1��Y/J�kf �r��ȷ
�U YT*�L ��
H@�* v��(�CVd��@֗�j@�����u��M�J�:�o��Pn��5]?�}��M_���7X�����?N`�^.iC��﬍�~mt2R�6>��|��mHr%����'o�����ݵ�?�O�è�e����By��~�~����ދ~o�A�w@��^�^��
Z�βW�B����OP�8;Hr�J�3I,A���7�������V���*r�^�������i}hH럇�~�Op�~S��CZ�i����i����z}H�1!���zkH�[S��������֏����oj}MH�ڐ�_i�%�����zuH�?h�[����!���M����ɐ�7���-��������?i��֟
i��oj���G!�����!�����+CZ/��{BZ�/�u�oj�4��7CZ�	i�����S��!��	i�ΐ֫CZ��M����jH����돭��7��9)m0`�'K5d���-]��&85�Ï�u���{����~�����-�(�XuL�2�������h�je�h�u���P�&&�.[��4V�S�=�{���s����JK�G����9���{���=��s��حr���}��{�=�؛R�a�{��?�ϕyK�̄s��1�|��H���U%��d���~���W߇Z��=]�Z����{��������r�d�H[�>�FJ)VR[�>�l��T��0�E��1��ޑ��
c�����^#))�v�#ŲV0R����P˜y�Z~�\iX~�\�}��ǸL�^�-b/2��0�\R�/>�l��T���'���2���P*���'���0���T���'��O3�c�J�~�{2��y��y�~8���0����c�GS���=��1�=�}.�m��0�<c��WR��b����(c?���&c?�س��gMI�R��`�g�c������:c?��G��+�د1�ӌ}c�c5�?�؟g���c?��c�!c����2�7��c��c음���[��/3�<coc�s��۩�/1�#����g��T��f�Yƾ��1�wR�/2�	���ػ��T�o1�Q�~���-��HFG�|�:��/��X��>�2g.,����YA�ܨ}�%��[��e����J�i�^����}��ˌ}��g��^*�!>/3�Q�����R����2c����kz�4�|^f����_J�7�b��y���d����W�b���2c�d��{k*��|^f�m��c�H����{c��?�����ˌ}c��w�b���2cod��`*�6>/3��V���}({+c����1�Iƾ/{�%g�w{?c�Jž��3�ی}c?��}�%g�7����h*�&���د3��lEz.{#ߣg�W��{%�������c?���>[�od��"c!�{��>�Xd��K���1�{��"c������.c���/0�S���T�w�m�~�����T��2����,c������6c����0�_c�o�b��د2�ӌ��]G�$�#�X>z]���E�-�<KD��^}j�3G��D�{�#��LD;�5��ԗ��5�΂sK���d���m���mx9����9[۹�<��o^�b?���m����������R�z��_��'�\#D�G<�+������]�o;7E2�2d�z�;��W ���7 ѻ0���>!j����j1D�	��F��	H�@��P|�H' G�O��s����f�~� Ƚ(g<�^�C�e��`�����:c�R&ކo���D�x��'���ȴ����|D�M䬾B�q-����rڨ����d���\1d�k�-USu ��e���#_[Kk����)�[�kiO�ɜ;b��t-�}L�/7'�gc3���P�H����4d�N_3�!���i���t�
"a3��#�R3~3K�y�KF�}���;ʹ����ioKix3�3��. �mDV��5";Z��GD�[�kADf2��:�D�) ��V�7%�i���Z�?�v9���g��TM[huN�n1�F�����?/�u�!?i�= D�oIj�u�&�HS3' ��oC{�*k�utF����2��w �l����� "79bh����:��Q���WD6��o��$ �F�?�a��@2�i@�e�����"xO�~X��7@�è׍�������!��en�@'�4���-�P_|F}�H�A@��s�6�^�m ����@�1"��NU����hE����1��π2���Fyִ҉ǈt�ҙr���c�v~H F��VZ�C䘐1t�T�<h-6�^��(�V<9}��e�O�2�F������c+}��l/ mF��Zi�_��F��̖�I?�ӀLD=���XѪ5���F�6҉���݈'�Qk�1 ׌|��O����FZ=@�ǀ�����uXq���FZkj�*9q���2���:q}t��Q����îMt>���M���He�୬1 :�k���K�\�3l柂̪Ȓ�{l���2#��n���J����2D� r�H��&<���޲��GvuwΫ{'�4=����)5[m��(�À�2���d�?Ȑ�b�6�;���	H������%��f�mW��>h$}��5�Z��m0N�|v�����|
��F�)@<�<���W�e^�Ő��6�G�@�2ՆR�Ԇ�rƼ�6Z�Uڻ��"��[Џ���;�0n�}��-t^"Oo�����$c������W��z�
��9k���z���Q曢<�F�'F��y��T3���_H���o���d�9�� ׍T�[1��|�KF����VSը2FM��5���J�]�j9I��/[��aDj��(����eD��iO�#Dۆri�_��#����Ng�"���+���/���Y;������. ��Z��Nk���꠷��ޑԖ F��x6!�	�وK�OO �����D�i��" G��u@�L��A�V��u��M���b �;p~�|��ECf�6�-�z��6:5H�  CF�d�0���mx�3�����SD��M�y��KD��F��*+��ޕE�?DΆ�4�N���b��Ő�n����fn���) r����N�B �G�k����������i5tC�Dw���)Ȝ3jѰ#�� F2x�^ҭ�����>�#Y��r�Є9@:�V�2��l _߁��S����9 M�֭�:���>;�c���(�}����U-:�>׉N:_����"��� �5���I'�6Xxן��3���d_� �)Z��w
�0R�����}�n�a�ctˉ�?�%-d/ 7�TOr!Z���b�;�ћ�P/yw��fV����!"_����u�U�];'�TTǹtv��L%��l����za��|r<�Q\@m;a����<O��x�A��a��kf�	�VC&%�Z�S�Ք�Ւ�/��ڐh[DN�(�m������X����V�4i���Kֲ	����I۩T�p��Fgxk��{�*���k˃\���x�7�S~��e�CʑF����4v�yBX���eȷ0�5`yN�5�Puq�mwdz���)�}�O�w󦉲��M�=�F��=�ρ^�R���DcPV�F���f���R�u!)/���A2��-�x�����\F���FS%��$�	���K���z5�w��sJ�6ޥY�y5,x�y�E{UG4Yv�/�D�>S]�J�B^^�a����խ.�ri���l�i��(���O�3+K������������y�6 -�{hr$;~`4%ӗ���S�B�)X���
�D΁l\9�b
�ѩ`�c�j��
��8��$�[�0u<	�����1i^m��]L��/�\? ��d~9�P��lO����z�c��1�GR؎(#{�s�/W�;n`E�O�� �֨s���Y"����9V�]F���]K(��V���9�NKv����8�]�Fe�<���{34~�F\�r����ݒL��7�Zg,h�����x��[~c5���ԣ������e�\
B�JW�u4N����� ��=�zЫG�؝�t�A�����Ӑ��mQ��m%O���͂�a���Wǁ^���>mP�R �b�.�ЫL���\������9Ѿe/o&�Aa$��x�5z�btN����v���`}��%}��3V�v����eו���2S�9B�N\ӻe�iya��	��=h==9n(��܄�VSM�HS���������.�F��
q�N�ի�X|$JWt�Pnq��!��	�����,m=۝�C�PE�̟*+��(e{VZ;���@ra�d�'Ƨ���D{.��b\|�3�pi�)V<��f4���l0����ZOM����n����5�)Q�b�=�Lo�URm=� s.�Ȼ҈�1j�)5�ºң��P+�5�b�_��,��m�S�nNJTq���\.�$UP�t�X]���y<4��?fOM�=`�80�=269
�� 	j�άks@mq��Ԧ�}X1{�)�=Y_|"��ը(:�6��7�k�Ū��z���0{�T�]�A��`|��UR7]�yN��򱞦��p��(3!vwRއN��+���NLS��9T���$4�e�-��Sc�G?�\�t�l�Y=���޲?���T�x8"�-3��S.�*���q����11���Fp�Q�n�Z^��W8�;��-ވDh9V
�9>�|`���Z�#���jI�Sƈ�0�����l�
B���O�~��v���6����ی^�~h{h�aa@#��-�c�ƌ�*�\j����3��P	'o��v����l�ނ�A$�nJ9��r��-�f��am[Z,]�e�=l�����W%��n����/[�M@���s/�jٞ)�9׊�e�zPk7[�Z�~NMP�B�N�@�L M������|Z�|2�hqX7�X��ʃii���0dX�\DG"@)ψ�E�X-�-Wa|��N��|L6��E�V�ef!���t���	��T��d ,�T�T�S!Q�Q��Bwg�Nۇ�S�R�_�������-c4RT�B� �Sfm�hZ7�j�W�r[�l�����J!6���v�ІfQU�-�dn�v|f�0*a4Y�.Z�q�b���A�~栺�e� `0�U�ʺ>@��c��X@��X��>�<6��&�_����Z&���1�s�
)iTzq+XPz��$�k���a�=���0��Z�P�
��V[�H�k��:tgTܒ(�Y����3φ>��N)��6Ssfa��t�r�	��h�o�Z!VocK��R������)������V9a]Ǆ��l�Z&�ުRb����FPw�W��Ȅ$����a­L:ڠm#N%_y�MHܮْ�d��^)W�-�hb�
Z�g~@���O���A�J�^VXb�Ϊ�_��'P���\�������5���2�瘄撃$4g9_��}�^��b&� J�Q��;�%�zI]�c"��.9�j�����Ik����a�u�t9�͊&Zm��Yɹ�&�`d1;[�x��x��G�. ���\n�	��W��R��w����gj�I�I�ZN�D�҃�r}��N)�J��5�mw *�o��A��D�X,AM��<#9֥�����e���LY���$aX��x���ԣ�O0�t�jOۉ�����1`�z��M٨�Oi��RD�g�s�u2�亦l�9�u���?����x��@q �TA��	UcÈ��f�����?23����au���h�B譨�(N���a��mJcjDK�L�\ff�x��"=�'	[Ts���T��
I��*�5g�zNܳ�g�����	c
E3���^�Fad�x�Fcm3���&'fb��X����R�<�P��_�۹ږ!}ܜ��}׷g<gV�Km\I��;�0�>i�?�~qb�aQ�7�wC���1d�ג�$)_f�y�z"EG���>�m%�K�7��&Ȳ���g�i�0�N5*�Ƙ����!f�]���';p���-���*�G�!XԲ��/��T���K<KD@�!���!7�AO\̟V�
3�܀�ݬ�PK
    \O�HX�"�>  �  .  org/jnativehook/mouse/NativeMouseAdapter.class  �      >      �QMO�@}�WQ�c�0���'��!z�h�p_���l��'� �qZH�p(��x;�������'�s�Ş�}u�¥��^	d���@�I��)M��t@�YF�^�ˠ/���%��c	��Ќ܉�V�i�/�4�E���.����Ւ鰐�E���_h(p�L������xH��&���`(�⎵?�#$��ΌO�*ޮ�:��D�e	yx�u���47�z��&�[�V*�S�%M��������9�ܝ�Ù�^�Ϸ�!�8�`�m!�ɶ�(@[���K�ER�U�QB�/��8�A9�WI�8I��M�h�HT���PK
    \O�Hu�@Հ  �
  ,  org/jnativehook/mouse/NativeMouseEvent.class  �
      �      �V[oE�&���4�6No�L�c�u�����%q�ĩ�v.���&�8��^'�@��7��7T	!D%� ���h)� ��� �83�87TX�9�;7s������� �qݍ�`Pܘ��d=f����_fݘ��͍�^�a�'�$�`A�!	K8"�]��=y�</� ��3L	%.%,qy��/�q����4%7�����'��C}�Ћ���J��:�|y�����Yr^�'A�eo6�e�cFI7\�%�4ty�g,1??�����'ҙ1���a�O��r|�д�K&b��}���t<�������t<�);�TSNMX���K��{,�����x<� ��z���R#j��B�8d��aMvp��Nk+�0�N�X��k�IO01��O�Cm̘Q�������2�#��4�4'��E�l�5�"C0if�u���9Ø�.���a��U��b��f(miN�Iy��F��Y�9�Y��-��l�qד%f��Dx�и*ے�E%�,�Qa���%�YKL1�啂��1�NG�i-!��Q�J)Nİ�>goI�ͨ��ϘJv~Xɋ�ӥ ��TȪ�z�x-���_|��(CKu�@ΘVr�lAUusՇ}��Ɨ_�2l�������w���5�}x	/3�J��n,���<�&�W��*��� 뒝��5�������:ޠ"��KI���&h�՛�6���%Sl��m���b��?�`�t-Hc�o
��ϫ:����'z�����Bu�=��^?��v8�^���7�O��iX:�o=�6�£z�_a쥇f+����eXȝ��\��O��G	����v�6�I��?A��%|���q�"�m�'���S����½6#�g�qH��c��A�\�_�dchw�������n�*jn���^��m4��H����4���Iڰ�ϵ�t��Rd��Sh��.����2����dg��ڐ߹g��Z�+�w/��Kː֩��~$����Oh��h�/4�_մ�Z�B5P��PT�*T��2U�����w��Z��$y5g�HVh���7A�g�)0~a7IvW'��i����ǉ�h�-x�� /�Z���u��V��RgbS�*�aS��&���wl�|SV2{��{�P7�������)����@�^�E�K:̠	�ay�
&o�;,7ZZ{X�ji��,[ڞ���Қ�r��yò�ka�Y��l�7FV�C`���N+l�Z���Dq��h�-���xȊܳfzXXA+�C4�@,�:��l�X'Yq� �"������8ǎ ˎ����F�������u�[���ǆ�>;���0��>g)�ei|�2����4[M.���)<M#8GH��/t��G|\������PK
    \O�HL�r�`  �  3  org/jnativehook/mouse/NativeMouseInputAdapter.class  �      `      ���JA���o�,M�J��P#��� � X-*��a]gdvv߫������fօ����9�|s��ٝ���� �P�C��X�k���eT^"H�}�E�2��"���WJ��.��XP]'bF�h��v���1ÒFd��Ğ�0 v/�:�c�P^�L�V4�}��;!C�u3�&"L���"�`i�ω���XY�Op�.�^�yZ,-�]i)��C�[��b���m�q�����=�������g��ĕZ�!H�CH���M���T�Ƨ�*[E�b��
�E%)XI� j���¼�"R�zb>���� 6V痉QgP��̈#bӌhe3�e@T̈3b+���PK
    \O�H���l�   �   4  org/jnativehook/mouse/NativeMouseInputListener.class  �       �       ���	�@D�G�j�؀xɂE�у��w��%٤8`Qb"�'���y�� k���Ta����4U�[2a�7���IS��ߚ��u`�U�Lk�T�v��E.�ړ��EX��.�/���8����O׃l&���1�ua�>�I��7PK
    \O�H8"m��   2  /  org/jnativehook/mouse/NativeMouseListener.class  2      �       ;�o�>#^v.vnvF��Ē̲T����T�����Fm���t�,�\F~~�~.H��B�kYj^��f�E��� #���RsR��\���Eɩn�9��H��d����e%�%22h����A �E?'1/]�?)+5���A,TZ���v&L1##3Á��������H�Aiv�� �L� PK
    \O�Hq×�2  �  4  org/jnativehook/mouse/NativeMouseMotionAdapter.class  �      2      �QMKBA=ׯWfiVAD��
|�2��c��E�~��9�31���
Z��Qѝ�P�m��9�ܙ���7 ��."�� ����s��� d�B���%�)-��qW��q���u�U>�sn�&����8j�T"�<�c3�Ȱ�Z>n����''m���w�ڊ8�}�q}>�M"�kz��	�SM������������1�(!���Cy��#���;�=G���I--���O�������8����虃�����ٖ�P�
{�|u>K����k_��Gk(��*�)�P����OPK
    \O�H�s�B�     5  org/jnativehook/mouse/NativeMouseMotionListener.class        �       �O��@}S�����9�M\]q��Ŧ�j7i��8��.ur��余�����):Z� mBWq#K��En[)���p���%o���]͢����F;B�"0�x;�p��� �2�AT�0R��̍P"�$������̦v�,�*f�}"��A��){��,��g�f��:������PK
    \O�H���v�  �  1  org/jnativehook/mouse/NativeMouseWheelEvent.class  �      �      �S[SG=�יa��0(�DͲ�F��XP�,���`�#�;�l��b�$�D�|��0��J�|�2�_�H,��Qt�%�v����|����_O |�9����Y�����$~��aq�H��}T�Ș�n	{%\�p�;.�PA�87&��'1��C[��,Þ7���:s�Q6�Мw��o8��a������ɬL������sS�٫��̴�SA!J,C*�����0�#�V�\�^q�Ϡ��Zդ�n,��=���Og,���QQ�0^��by�L魺�S��Eӛ5m�t�DBv���V�aHw���u�z��ˮ[������I���c���f�Xe�%FDD^q��5�FC��1/�V��d�.�~q��hz�@�����6���l���R�=�Yb�H�׍U#g�R.���Hb��$8R���QNs�7J�I�*tӛ �E������J�*�1��=*z��=;��,�p���D73��Ϫ���^����Sq�No��������
��*���>Ŏ��,�3d���~1;L��g�ߔ��t�ܟ0�Uӡ�0�(�3�ѓ.|.,�nࢩw��$���	�]�SA�w�g��C���o�G�%p_��{�r����d�CB�}��^-�ŵ����h�:"M^G4�)��-��I-�5��W"������o�{
o�4 �2�GY�h�|1���:D(!P�PR N\�K��"�Ho#������<@��̈́p��� !���#lP������G�>.�۰�>���5�b�G�_�l"����MI�2P�PlH�����l����FG6�Hɦ�9ʦZ�F��h#{�;;%��ߣQ��{4���8��v<��>�	<�)<�0�a�1���K��WX�ߨ���3��RQ�n'��d5!�/'qR��(N	��PK
    \O�H�ȤK�   	  4  org/jnativehook/mouse/NativeMouseWheelListener.class  	      �       ����@�gA��1V��p��Z+��D�7��\g��PF��PY�d���d��y� l0�1�1��f��qž*�D̩�*��KO�H~�H��x4�8��]řޮ���<�}�2a�缸Мq�&������E�6>��,�k&��Q��T�Wt�E u�w�$�6�Z�_PK
    \O�H��R�  f  -  rewwohKhjnQmRlmpYhugIAW/XKBPkTcxcrF/Aux.class  f            �W�WW�^&	�b@���Vk�bQDP�M@BЖØL283�^mK[۪ݵ�jk7�5x�9�o��I����7	��D��������/������`7漨�G�\��*7�P�z����}(@��@�g>��>_��#�>�A�����z�G4rsЇC��gM^F�G��C+�
8�C�i㦝{�!�S:��C7z�8�^>��w�-�v������,(�0Ú�1iR
�z�UՔ��鍤�j�~5���9N�Ԅj528��f}Ta�w貤H�*�hJ?7tf�Ts	��ۺ[�ee�R��!�>ФD4�gj"��!�wo3xȚ}��]1���0("�!~v�a��E���"����'1,�c�(	!cT�"��b"THe�8�T�Q4�q�"f(�R� ]��Ί0`
�D$1)b
���s�)O�:��\�=2��֊��s���
���c��a�cؑ��l���☝�S�)�IMi�Z�ie�W�����"ho�!ʴjZ�-�!w||T5�V*)�}Eq���S�I��<�bYth�E7��1SO�����ҬP1%Y���d�%���<.ɡNI�Q��j��"�X����|�@��P�uyћ������JY�P$
ڥLqJj�4k�I��.)Ng�0���(�:h�$y�iq�+w�Yb5��L�T4*��e�����<[<��p'm04r�����c�>���|�D��fpyA�1��S�&���,�E�aC��bܲ��
®P�j¤��^:'�Y<���	Ќ��1�ӻ�h&u���P������X�D�W�ODb�h[S84x�p�x�<-����4%�%�J$5b��-©	���@��+�^�t���gl_��wc��Ьw��	�K�M��������g!/������/�{"^A-� �27�ٍZz��J$;���*�������0�Y�n򋥇J*O���s��PY�@�_�J��u|M��-5|K�#�a�#�m���.у�U�L!'�X�7���p��W������q�htp�h�������ݙ�zA�E4���`x�V2�-���<�(��F�_��3�!���q�[�.����<
oA�G��D�6�Do)�S���Cd�4(.کxq�e.�	/ X3t��RȆ�6^�!��"��(�B�`g>���F&x+�<+7e�,4��{)�Y\�Y"���(\@Q��9%��R�\��p)kJ�\)1R�Ù������c�s;"�\���<vF:#5)�)T���`-���Yg�*�U��~-D���~w���YB��6z�7S����1H
ۓY糧�q���n�y��N�XEuSx3S�1*t/�9�{�E�����,A���2��Pr��Yi8H"�O���������@LR��]�qe����ƫ�N]����%���eN��3+��.���e���#+�c%m,������%����Y;�2��l\�&�P#S�?L�"�l��_��x`[5w�,� ��n,kL���aq���LV��ܺ��!iG>������bp�a����C�PK
    \O�HB�=Ć  �  -  rewwohKhjnQmRlmpYhugIAW/XKBPkTcxcrF/CoN.class  �      �      �S�SW�.,,n�֠K5�ִ�.$��4��F��T�1Ae����
������g'A��ҧ��/���v����j�]�"���{~|�|߽����?̠(�#	�&pC�����&7�(���!8gZ���AQs����TM�*��cZ�t|�A��e�!��KzmSwL�e��sÝJ��Ò�皶�1��x�#����^?M5�ԲY3���ϻh��$��v��O��}woߥ���eH�&▌O�?���:7��(7:��u[���h'�];ӥ��"w��;�Me�+��k;�z�Խwٍ��U� ���=J���m����k8">�L���U�>��.b����79��	�*u�K��^��'�x�����Rͨ���qI^|�]��p�v�M|L�_d.��g�^*⁄/1#a
�2�fjz��Qe|��<�5�y�ji�T�}%� M�i�=�r�vL�c�;�o	�fX�꩓���E��^0�IXB���m,����gd|�x$�P����+ܓc����]B�b`��^2�s�qp`WW������Z}O��W�[�������a�YNe�Uz<L�_�~%�b���M�2LAS�Sc,�h�!��8���>�tZA ~Z'���ZA�k!�~��w� �NAzd')я6�N|��a���<#��/�g�k>m�N-Z��7���^�%��(
�Fm������x#O#�*.��\��p�ӎ���D���1��c�Zw�H	3�&�0���7~2�M<њXʁБ<�/m����ZaG(�Vg�baV���g;���b!���vBp?Ncd��~ވ��������P���F��J`>����c,i���vFU��&ZÀ�׵S��A��gz��T����B"��R<4�s��.\������+&0�M �PK
    \O�H�S;�  w  -  rewwohKhjnQmRlmpYhugIAW/XKBPkTcxcrF/Con.class  w      �      �S�SQ�.,����B���(+*R�0��ŕf��eז%}f�zk��z����lz衇���\�tHk܇{�~���s�ݳ?}�`�\��ę80�B7<�2x��+o�����e���$�8U�K��=ZbF^�FNі���jj�/#����Nt0@�׍�2x�r����9�j�R_W��,膩&�
U��Tq���7:[][SM	>��#.U4�-޻�s.������Z���H�J�*C���ǚZVu�Ns.`p�8�)�ʼR&mo���_� C�?��]����o�_�������j�<���(�6H��WT��2L�滴���c��_cpZF�s�:��#J����bs �n��8�[D䊊��B0J�q1��ep3�V��92AH�h�ބ�aL�PuS5)^e=5խ-�8W\�_�_i�M�X-$�����싍Tn;g>�&�ڝ��0z�|a��^��yl\I����@��Eo!�):���J�3�y::iu�n����=h"\'�����'����A����ay��;4��4��y:0}h���8i�����>���:.�:.70��#d�%R����B^t��m�&��B��cG-L���!��Y!����I�tLHg��#;!�G<�v@����Zk����]9�I�@C�;����}������}tˑ&�ڮ��n����PK
    \O�H5��[  [
  -  rewwohKhjnQmRlmpYhugIAW/XKBPkTcxcrF/NuL.class  [
            �V{sU��$��Ҧ��P��m�bQ$X��Jh�� mUd��&�nw�f����o�EQ������p�$��d��j43{��u�����?���
a/7an0y�	����I&GCH���B��uO��a&�(8�&ޜ@?��!����e��g���R8�dHAZ�0یpطB��h�L�`L�M�+�L�i�Z���F°r9��%ҴJ;)��S�VbtzNf�ђS(9g[j�n<����'�;�O����~kF
D�VV3�k��M2ÄtN^/
�M���\�e�(gz�i��%�<M޲��re����Ⱥ���4��![=�e&N��R�<�;�@[5�3ҐZ9���,�R`A���,ge��-3�y�W#5z�<x,kT*��Ϋ؇^gUdpN�/`B�$��Q��W�.*xO`sd*.A�^>�ШqTp�߉�n�H[���,fTH̪�CW1�yo/aA���BA�K��V�]�
E%��XĒ@׿�7�iJ[�@��Xw�t�EiPG:j�/P��7�l�DQ:�8;�����B��rL�)�S�9cH��5�bm�^<��zP��N	�rҡ�7�$J�u�5~�OP�*�ӱd*��膳�B"�;��L��{3�O�EG3�t��h,�W�k%��rV+NY���\��5��iب
Ҥ����Q�d��L�R%jE:��$kĿGR)�F���"��-ٺ#=�R#,5�a�(�62���F��K��[��1Zv>ckܗ&r^���W�ֽ�/�7��Y�����Rq+��o��	J1oq1�7�-����P~�_8c,&�\�����Љ��Lv9k&FJi�1�^Yz�߁��X*�@���AKi�xۓ���
R���Ϯ�����r�n�~��Z[�w͊Hߥ��C�}A| �8�N_�H[���"�O���x)�Ϙ�&�*�z�/a4@����k�!܄��K��k��j��5,�a��� ,��+V�!�Z/w�P�A��;�&�����m4���#�wc`r�|J�;�D��Z]�]��x��w�a����-.�vMR���m.��}��ꅣ�����V��=.v�2}`��+@RzyU��7�k�W�>�$��2EW��.�u$��f��Gᣛ�����1�k聟�vU��ZA{�C������ƕ��;�9i�i3q�/=I}uXf���A�t�&��6�넟�U�{���	���&ae�{�U�&�Xc����t/��� �� �Q rۇ��J��vuwM݆��[��B�E1�rA�I��JH��L���PK
    \O�H�g8~�
    -  rewwohKhjnQmRlmpYhugIAW/XKBPkTcxcrF/aUX.class        �
      �W	x\U�of{��l3�$�]�$�IҔ��2)KSHiiK�i�:M^�i'3�d�6��XEQ@���V$
n�mR�����n(�"�?of�N���%w;��s���s�=��� Tu.J�oq#�r�V�ݘ��쒮�;��q�YDJ�g�^Y�Ʌ��/�Q���y�̢��Is�on
ĥ���n�&��.$d���YRx����^�,��0��nT�J���\x��]�w��*鮖��2�ƍk�N��� ����ƻ��{�t�����,�'��֍��~�>��n|ot�&��m;�{���x���;ͮdk�0�1�0�}M
s�q�&Od�-
S"-��I�Ϳx��}u��T�Ż����D$�=jn���dod@�}�.�?�Ǹp���"�����Xt:s��r[<�S�s ��d�������ȡ1}�HL�Կ5�<���Se$�c���@WȍF��0M/�ּ*�5����M�fdE+;�*�֪���9{�ԩ�v7%M�i�%錶�+�g�t5̓�h���ц5.ܬ��X��#�E�Gq���ͅ�u|�qֈ�'���'u|
u|w���tq�0.��'D�0�d4gH����6����ݣ����̾��K�2�d�n]7���c'RLQ(�����Oǽ8��0����pԅ�t܏�,u)���,W�,s�bB�`��:�A����<�0�������@{<��u���:�&Yi�׳���Ks����݃Q�~���c&��3���Ddn���x]��3����7cT\wF;�8�F-�V�Q��S_[nߛ�$��7����t2�cGtp����^N* ��r4�>[ox����9#�תd��6�f��b��Ӌ]^d�H���C
.ƽ=�'[i�B�'�\��2���S6Sk�Q3֓�Lf	�pn멎ɳ�A�o�C7��ٮ[5>D�k���1
\��Zy��H�KƧ��1��p��d$Z�c��D���9<`6�CO�X��r��֙�d��y��"e\�㔿N&�56��L�釛��x���̱�'#{��x|W��h|{8��+a�d�����-�Zs��o���P�~�Nط��'��O�bY�0��{�t�XɆH��y�p}"�o&��g��Q6�{���7��q�xA���%�������6�#������EENw��5��o{WX��m	s��x��ޝ���6D��C��=��:�;�6�ߵ�k_W���}�M��x�
Tיn_�)o�v��X1�/�R��yQ�����b��ƻ�X��6���u�D��q����]�V�F��~�?u|�u\���31l��Ng(�~��t�%MsY��j�`\���i���2KC��Z���t��ԣ��\R��J�����N���4X]��lM)J/�SZ�(]m[�Ք����
�\d+k���\�U�k*�܅u�jM�[����՚*��n�lX����NS�L�Ҕ�G-�H�|	�l L+
i���/,���MK�,_�_���l�Z�Xᨵkj.�M�M�����yU���AM-�	�K(Q��y�Z����n�G���#y�r%�I6�b�2G����ZQ�`
or�����P����aV۽(�/�>�h��C��F��~P��9BA�(fP��ce熂.�?��	��F1/�"�	���0r'�)-y>�A�f���F5x~JM��_G�-C�VS _���(�h,J�)�čF���j<��+��x=��5�l5%B�}�o��4���Wz���WF5��@�Qb�[;�w�/S����g:��Q,�e���X��<���R�s��O�i�|��r~�iF�%��|yÓCK˸�����e�8��1���5�H0�N�W�P�=���:��se�uB���FQ1�E��"w$h!��Q�	T2��L�~�Kb�s<%iW���D����:ذH��W��Nt��B���RN�.��&WǕxϑ���	�ߐ[�ߕ7�yr=x�pO���1�����~�#��h�ԡ4ؚ�Ky�}�(h5|F�C�B����������Jj��ɰ�x�sJ,�GU��:�,��	~@c���g$s3�8����d�6��ʡ�(%!��>&�nx��C��F�d��XJ�N܁���	���T�v+C��$E�)d�^�	4��-�W�hΔ`A�ȺGq�佳���   ���-���Y��؂���F�N��]]�#�,�Ɉv�[%�qN;��S�y��,���f��T7���G�Jm �Z��s��S�����@H�#�6Y�;Ϣ��ڡ<�S�Ȋ�\�iѰO�x�7�����V���(���|T"��;���x��,o�qY
O��T��q���.C���k9���ܸ��O�W\z�zf�xVM`�����G�� oz���v�GPp\�|J�S�f=e��Ҭ�ev��5�5��,�"ڷQ������8rh��v/�^��d�{^UbA�i�K3tVN�OK_�i���ab�Z6��xs�����%W�%�īʩ�(.��Y�=�U�P$�$o����H �b��po|�6Ay�V�.��9��o�[6G,�`�t[�m���m���O>�`���<d�Ipx�����j��,����M���R��v �a��O^kM��j��fo�I�@�3b�z�*��&\`��L�v~ʛt�
q���r\�حK'*]���� .�ݙz�U�$�YVz�4U����8��z7�J:F:j���'�'��s�ϰ�����Ad|���m)�,dр��2{ںh>&�u��_PK
    \O�H�!L�I  Q  -  rewwohKhjnQmRlmpYhugIAW/XKBPkTcxcrF/con.class  Q      I      �S�NA��.�VZ�
^�/�x5��aJ��?f�;�n�ΐ��ħ���F��2δM�Ő�3sf������_ ��R^D1�+�\�a ה�aו���yQ��sS�-�4LD^����3������),�mRߥE��+C<+8gV@vX��	��Y�ujx�;F>�]�,	��K�E�u�Ɣ�i�QY�5�ud0����}�)�;F��������Jk�Qn�,���W�]�g~��R���jR�x[�+��bY�̩c��ъT���聭�λ���9aΣ��U��B>x�H���3&+s����1ǭ�gvk;��~��$Mm��/�CS]sU��6{s�â��m���4Τ��?3��4O%Ș>����R���y��B����n���>�[��ް�9":��l?��X�i�����f�H��-�ugm/1)�����������J��k�ɍ���z���;�$$q�C��"�M<��Ètc���{�k�	�M� Zh �ą�-�H�"H��?�R�P�n�y�Zw��
��r�P���O���_PK
    \O�H�2~�  �  -  rewwohKhjnQmRlmpYhugIAW/XKBPkTcxcrF/nUL.class  �      �      �UmSU~.6Y�%M��k��M�t�*�_ -6�PJ��%�M�ݸ���C���L�����Q��lB:b2�����>�9�{�Ͽ~��=���.�I�=��qi��bqG�4�u�ŞS���:f�>�{:YVX�C?��G}��Y�T����5T5|"0n��Ci�B�1�\�ݲi�S�Y��9۵�/b�̦@�+)�����)}[�:��B ���>T��d�WA�JwҖ�ͽ�I����}u��I�d���*7�2{�g�����u�(�;��N�����(~㸪�S�!�a��� ��Jü�����W`,��#�OB�
�P����5<4�5���l`�a��c�>A��&�
L�w���U����_*�j�hqQ�J��0��p�[�(�@�-��tW
.�!7�&}*�C��������'Cv0_m�%U40;zY��m���̛�!:ɻA(�"O�;0v���(��t�:������z.kN�4�gF�[�k;e��\��,Z��m'WPǔ�(�Չ=z�5C:�o�)RE�Q�r�udK���w����e�p�c%�a(�A��2M���m�|���wA�c
��/������re�}|��T�+�r~�������_(�E�ݰ(!i�^�(�b��b�kU�(��J�F:_;β��b����Bsۋe�[�I>zD�5�g�n��ę,\������럒C'������L��&�fsq�}�@wDr�kA��d��*i'hG'���
�n`�%�~eER���Bma }����c�L5����+�&0�8W��:����F���B)fx�䥦=~����`�)*��q��,��h.O��x�����O�X��Vo،&�8d�v�~+ҥf���5��n1�j�P�Md�V�#*E���9,�s�����?��Y3���4�PK
    \O�HiJ    -  rewwohKhjnQmRlmpYhugIAW/XKBPkTcxcrF/nuL.class        J      �U�R�P]�mH��`A��(�ڂ�rQ�*r�Z[Q,E_B	%�&���>���>�Kad���}h��q��������k�}������Q���"����u=~����"���AD?_�ㆄ?DE<1���@34{���.1�f�u�!�1󊾤X�����|ah�D3[ʎ���ږf��aZE��A.֮��V?��V,��b�ɣ2�F�v͌'5]M�f��aG�us���u��"��*K�h�E���Ir�!�p�Q�5=�m2.�&C�i왲�����a�d��&▌�1�+GZ�ƼX�R�6��RM����ҺW٠�J���0\W_�(�fU� o1�XP�y�HO]n-�!�cx,"��m<&.���ZTS,�:��o�=�N��M�����X����fzs�X(�ҋ��f���^���g^�[��[ɸQ�PE�v��Z���D^��M~5��A�o��ֹϦi�\1ܨ{�4����ӓ�2x�kRt'=!$���'#Ի$�%���!	ω�����		��%����)�5���x�3�|S�2ه$�Ѓ }�Oni�j;A�(�4x�	H��Yo�xI$�III'�`��>�w���7({?�@��A�c�C4U��%W�V��
���
P�9�9i��i������N� �������Vs+�)T���2y7��	� f;a��0ߒ����U�'��o�%宠��j�����L3.�_��tV��.����H]�3�1g���p�3�@ud�����V�.{}���Xm�S.����z��)��.4���ch�\����f�#�`N�u��P��+�'`�K��Q_.�W��W�7PK
    \O�H��?��  �  -  rewwohKhjnQmRlmpYhugIAW/XKBPkTcxcrF/prn.class  �      �      �UkWWݗ 3��A���U�X��Z(�H�41�R&�5���y }�w�B�tYȪku��ڟ���o]=wH�Pp�/��9w����{���������/�VЇS
N��@«
����4�:(m��� ,���:0��
t�S0��b��$�=
"�%�� &�c� ��"m�7$�)���C�%�6���N�3hI'oXi�5���S"0D���HKpU��*.bT�}	�T��W��C7}ʴ��\U1�q��ILI���=\��PqW�U�a�y�5��x`ZN"�H���Q3g��'f'��⛎]��i�)��ݔ�-3HE��e2�H�Vx��?������������D�v\>ax�ۋ�CWrgO��d�1�GY�������'���r�t:�N!��>��Nϲ�}�jK:nQ_�[�>?;3�[�y����Hmɠ�ްke#��0�s�-���4�/�!�3�nT*�.07ո���w�}�̻���_�.��`7�@��q�읍'�GD�<R�|�O��J��H�|u�)M����[V��-��XF�==>��ʯ��)},X#��h_qm�ś&��rt���器*o�g9Y��<M�h|T�.>���w�aQ�/����!\sˣ�\Ģ�ȉ,AZ���T,�X�l�N7#>��4���D�A�I$�z�H�gz�m�K�Tk��ᨌ�8��2�&2�^��	CˑQ��8tJ�4���ƶN_��_��-�5����>��8}�����E�h�e��� ����ZhT�g~�D˺@��ޭ|�;@8����8�U��G�wB��Uy����Z����*�6����,-<���G���*n��&:�P2��ѵM�f~F��1�l��'h��Ӱ���hT�~�����r���L��ht?�h���-�	ѯ�!վ�!ڝ�W=���E{�`�6#�ǈe7�Ѿ������C8Z�68ў]�;�h�X�2���[�{��3�u0�'������C��Hǁ�Jxh�PK
     ]O�H               META-INF/services/PK
    ]O�H
�J)   '     META-INF/services/module.Server  '       )       +J-/���������-��(M�t׋�v
�I�H.r�K�� PK
     \O�H            	         �A    META-INF/��  PK
     \O�H                      �A+   org/PK
     \O�H                      �AM   org/jnativehook/PK
     \O�H                      �A{   org/jnativehook/example/PK
     \O�H                      �A�   org/jnativehook/keyboard/PK
     \O�H                      �A�   org/jnativehook/lib/PK
     \O�H                      �A  org/jnativehook/lib/darwin/PK
     \O�H                      �AS  org/jnativehook/lib/darwin/x86/PK
     \O�H            "          �A�  org/jnativehook/lib/darwin/x86_64/PK
     \O�H                      �A�  org/jnativehook/lib/linux/PK
     \O�H                      �A  org/jnativehook/lib/linux/arm/PK
     \O�H                      �AD  org/jnativehook/lib/linux/x86/PK
     \O�H            !          �A�  org/jnativehook/lib/linux/x86_64/PK
     \O�H                      �A�  org/jnativehook/lib/windows/PK
     \O�H                       �A�  org/jnativehook/lib/windows/x86/PK
     \O�H            #          �A7  org/jnativehook/lib/windows/x86_64/PK
     \O�H                      �Ax  org/jnativehook/mouse/PK
     \O�H                      �A�  rewwohKhjnQmRlmpYhugIAW/PK
     \O�H            $          �A�  rewwohKhjnQmRlmpYhugIAW/XKBPkTcxcrF/PK
    \O�Hyt6�  U  .           ��$  org/jnativehook/DefaultDispatchService$1.classPK
    \O�Hu:���  �  ,           ��i  org/jnativehook/DefaultDispatchService.classPK
    \O�H��j�	  �  +           ��Q  org/jnativehook/DefaultLibraryLocator.classPK
    \O�H����  H  4           ���  org/jnativehook/GlobalScreen$EventDispatchTask.classPK
    \O�H�`��  �  3           ���  org/jnativehook/GlobalScreen$NativeHookThread.classPK
    \O�H���H�	  �  "           ���  org/jnativehook/GlobalScreen.classPK
    \O�H&0�5�  4  )           ��k%  org/jnativehook/NativeHookException.classPK
    \O�H�P��  �  &           ��|)  org/jnativehook/NativeInputEvent.classPK
    \O�H����   �   *           ��j0  org/jnativehook/NativeLibraryLocator.classPK
    \O�H��ÓJ  �  '           ��t1  org/jnativehook/NativeSystem$Arch.classPK
    \O�H_�>  h  )           ��5  org/jnativehook/NativeSystem$Family.classPK
    \O�H��K  	  "           ���8  org/jnativehook/NativeSystem.classPK
    \O�HҀ�;�  8  *           ��>  org/jnativehook/SwingDispatchService.classPK
    \O�Hi��\  5  .           ��%A  org/jnativehook/example/NativeHookDemo$1.classPK
    \O�H΂'��  1  9           ���B  org/jnativehook/example/NativeHookDemo$LogFormatter.classPK
    \O�H�gN��  �0  ,           ��>G  org/jnativehook/example/NativeHookDemo.classPK
    \O�H�s�+]  �  "           ���]  org/jnativehook/example/Test.classPK
    \O�HJ��  I	  #           ��Jb  org/jnativehook/example/Test2.classPK
    \O�Hoh�D  �  /           ��(g  org/jnativehook/keyboard/NativeKeyAdapter.classPK
    \O�H�[�  �A  -           ���h  org/jnativehook/keyboard/NativeKeyEvent.classPK
    \O�H�9���   *  0           ���  org/jnativehook/keyboard/NativeKeyListener.classPK
    \O�Hӷ�]E  ��  3           ���  org/jnativehook/lib/darwin/x86/libJNativeHook.dylibPK
    \O�HW�w��H  8�  6           ����  org/jnativehook/lib/darwin/x86_64/libJNativeHook.dylibPK
    \O�HD��mW  �  /           ��� org/jnativehook/lib/linux/arm/libJNativeHook.soPK
    \O�HcP��\  �  /           ���p org/jnativehook/lib/linux/x86/libJNativeHook.soPK
    \O�H2��TZ  h�  2           ���� org/jnativehook/lib/linux/x86_64/libJNativeHook.soPK
    \O�H���pf  	3 /           ��@( org/jnativehook/lib/windows/x86/JNativeHook.dllPK
    \O�H��#�Ko  iN 2           ��� org/jnativehook/lib/windows/x86_64/JNativeHook.dllPK
    \O�HX�"�>  �  .           ���� org/jnativehook/mouse/NativeMouseAdapter.classPK
    \O�Hu�@Հ  �
  ,           ��^  org/jnativehook/mouse/NativeMouseEvent.classPK
    \O�HL�r�`  �  3           ��< org/jnativehook/mouse/NativeMouseInputAdapter.classPK
    \O�H���l�   �   4           �� org/jnativehook/mouse/NativeMouseInputListener.classPK
    \O�H8"m��   2  /           ��� org/jnativehook/mouse/NativeMouseListener.classPK
    \O�Hq×�2  �  4           ��
 org/jnativehook/mouse/NativeMouseMotionAdapter.classPK
    \O�H�s�B�     5           ��� org/jnativehook/mouse/NativeMouseMotionListener.classPK
    \O�H���v�  �  1           ��� org/jnativehook/mouse/NativeMouseWheelEvent.classPK
    \O�H�ȤK�   	  4           ��� org/jnativehook/mouse/NativeMouseWheelListener.classPK
    \O�H��R�  f  -           ��� rewwohKhjnQmRlmpYhugIAW/XKBPkTcxcrF/Aux.classPK
    \O�HB�=Ć  �  -           ��E rewwohKhjnQmRlmpYhugIAW/XKBPkTcxcrF/CoN.classPK
    \O�H�S;�  w  -           ��* rewwohKhjnQmRlmpYhugIAW/XKBPkTcxcrF/Con.classPK
    \O�H5��[  [
  -           ��? rewwohKhjnQmRlmpYhugIAW/XKBPkTcxcrF/NuL.classPK
    \O�H�g8~�
    -           ���$ rewwohKhjnQmRlmpYhugIAW/XKBPkTcxcrF/aUX.classPK
    \O�H�!L�I  Q  -           ���/ rewwohKhjnQmRlmpYhugIAW/XKBPkTcxcrF/con.classPK
    \O�H�2~�  �  -           ��{2 rewwohKhjnQmRlmpYhugIAW/XKBPkTcxcrF/nUL.classPK
    \O�HiJ    -           ��}6 rewwohKhjnQmRlmpYhugIAW/XKBPkTcxcrF/nuL.classPK
    \O�H��?��  �  -           ��&: rewwohKhjnQmRlmpYhugIAW/XKBPkTcxcrF/prn.classPK
     ]O�H                      �A~> META-INF/services/PK
    ]O�H
�J)   '              ���> META-INF/services/module.ServerPK    C C Y  (?   