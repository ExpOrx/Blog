PK
     �y�H            	  META-INF/��  PK
     �y�H               gjjkAkGlNmFoVoKv/PK
     �y�H            !   gjjkAkGlNmFoVoKv/OzIRjRnhwqtFRod/PK
    �y�HV�;�  �  *  gjjkAkGlNmFoVoKv/OzIRjRnhwqtFRod/Con.class  �      �      �U�[W�݄0�t�0l�h�j�a� ��"%6��C�%$c�0̄Ʉ�Z���s����>~���؇���)=w��>̽瞜�;��ܛ?���w �A��zp���m���v.��*�W�t�/]"JqM�ut��A/_n�)�uo���Ǘ[|����"⠷E���H�ָt�K�>0�PIǗ�A��̦���39k�2��B���Y/،䬃F����Z7��/{��(CI��T䈑�kѸ��g5e�/D��-�{!USz�����z*HH��"e���Z�]��XI(K5t����XX�Y�D$aX����x�A:���E�[9UK*��Q	c�0���I��x�$L����E	��c8}tذBFNO�b�(B��=�5i��b� �I���q�$4bV@BB�k�x !�9	*�1������'N,ɜ��sI1�YŲ(�,/�a��鬡�4�JVQDM���g�(�ԡ�c�YKY��I)��/1����mi<�Qt"�z,�Bo��m;*�JQ芜�j���+���Rix1�x�x������aQ������,��M��\�\v���EPX�mF{B3����KQ��_E5���'���Ce�%_{��$�kX���.����G"�X��zV1ɠ��?���a�?b��i��<oU�kt��H*���/���1�Y��G���E+4j$���Me	�f�ӧH���პᣟA��E��p�?�'����k���6�]�]�n<��]n|D�Iut��a�Re�u�97>�*y/��7\n|A�k�o���\��=ޫg�.��f��wt�K���A\�s�p����(Uk����M�j9�k�k������>C��2�g	�N)�������2�S\p�~�%0��{
�S87H�p��F��SX��:/r�li� �_�W��q��({�s�-���(�?|��<N�a�ۢȵ��j�<^��KNy�<�#��X���v���+Ⱦ����-ԭo�5�c�}�ַ�pF6l�5<Dy!��RD�'1�kD�����@}�P�$������#Z��4����%���Ó�z'	��ih��R���\�r�e��<*��pm�Z�����a8A�.�N�N��l3�	?�6@]�p��߃D�$u�����wK�K���!�m����C>�@,�'��.���e�jK�嵜�4����^���Ĝ�p���9C�ږ��ATs?G�PK
    �y�H~��  m  *  gjjkAkGlNmFoVoKv/OzIRjRnhwqtFRod/NUl.class  m            �SKS�P�.�Qb���"����ZEE奵V�8�4�E'���DC�Ǹ��\����0�ǅ�(���P�,Nn�9�w������� 0��
|h��	2�x8���<�eL��`�F�v�chԂ�B�ɘm�Nڰ7o���y|�=nW�b����v-8]0֌�e��Ȝ����0C�c��6Ӟ�&(*NᴊN��]P��̪eF�Lw�t�3o�\�UƼ�yQ �8O�i�ZrV�J[W]�L%_���9�]W<å=:�=X]Z2]gN����\�57FF��^��82h�3���&�z�`r�S�J�Y4moX�y�qp?�J��e��$����"�ɕC�24A\b�k�Gp��~YA7�T{bz9'S%��f����y{���Z� �}��4�up�tB<�ZSq��vc�x-��z��	�����-�d2��`���9Í���T���ܧ��%cU1x&�p� �ȶ�I����o�Ad��Ba9�<i%�΢3��y�-�ڹׯ��Y'I,X������|�6�(4��̤	���|�������1��7����Z�!��V���1@��` B�־�=�o�1�	abR=���?��]|��R��WL~�CH5��ڎ=����Mܸ��_�����F���^}�ʸ $� ��T�)�,�^ƨ��|%�T��7BI�k����]��)!�I��g�³�>:(���O���B(���k�S�X*}\�����~9�S��;]T����������[xXo�i����PK
     �y�H               META-INF/services/PK
    �y�HE�k0&   $     META-INF/services/module.Server  $       &       K���v�v���u���.����
��(/,q�O��� PK
     �y�H            	         �A    META-INF/��  PK
     �y�H                      �A+   gjjkAkGlNmFoVoKv/PK
     �y�H            !          �AZ   gjjkAkGlNmFoVoKv/OzIRjRnhwqtFRod/PK
    �y�HV�;�  �  *           ���   gjjkAkGlNmFoVoKv/OzIRjRnhwqtFRod/Con.classPK
    �y�H~��  m  *           ���  gjjkAkGlNmFoVoKv/OzIRjRnhwqtFRod/NUl.classPK
     �y�H                      �A	  META-INF/services/PK
    �y�HE�k0&   $              ��=	  META-INF/services/module.ServerPK        �	    