PK
     x�H               KOtupZesZNNfLlSPIX/PK
     x�H            +   KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/PK
     x�H            	  META-INF/��  PK
     x�H               _020_/PK
     x�H               _020_/resource/PK
    x�H3i6_  �  4  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/AUX.class  �      _      �R�J�@=Ӌ��j��Zŷ�`�<*��bl����۶n$6&��U?KP� ?J�D�AD���9sv�����`��0�#�!���P�0�!G��v<G�R{��$��~[�u8��ʓ0�E[9�W�����P4/DO�V�'=e�F��0�Z���4��0B�E(Wx�F�u!ۊP��h:]%=��p~��W>a�<,��+Kv�R�6�j�aX��^�s\�Ү^�vNm�H�����E�,��zԊ)�[k�	~�t���rl��w��4f��a5��x�	�Ai�_@��P���`����~�֑�d�A+/H>pA�p��j`�3D��<�����$#���\y=#���u�q�PK
    x�H�I,9a  �  4  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/AUx.class  �      a      ���N�@����ZD��xC�;��zYbLqa�@DP�`J
��R�D�q��P�)Ɛtsf��;gr�|��8Ė�6"c!�y�Kؔ�'���BE��	I�n1���5M~�B��\ö*��m��ۄ��eC�����!�\�0��z��n���&���BB���Lfu�r��[.a�_P5.��Cf�����ڄ}�����j|��J�jV+g7����z�Ν��jԻֵ>.*���'P�'V��=��2~�y_���5�}�ӗ�*֢Hb��篳?@, ;�BaÀ�	o�pV@H��N|D@��l#�zA�Q�����
��Ln)с�� 4�J�>�r����_\����PK
    x�HZ��t_  �  4  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/AuX.class  �      _      ���N�@����ڊ��h�!$��Rcb�c"��� SR�����L4>�e�V���nΜ��gfN��Ϸw �XQ����$&4�cIANAZA�0�g���'$J^���Ŝ:�m�t�Yi���V�oy�oV�F�������A(9���:!;L� ���IB&T9���f��!�/hط���'��A�D�a�8�����o�r�2�Z��R7�^�Կ��U���]X�	�/��sg�@͈�A�2�a'������)V"��g��S��4a#Z�h��?֤���~e&�;��b�?
���hh�8br�
��3��G�#�2�}W0�Y ��d����~Kj�Zx_�����*OR��/PK
    x�H��7 _  �  4  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/CON.class  �      _      ���N�@����ZD�xWиCH��%���
D�� S,�V��X&���2NѸ0����3s���o� v��"��E0�iq	�ľi��*8-NH�N�YU暬a�so�9qm�	1��c��k8n�����LcC����v8�yq~�JH�(HE� I��T��Z���MAH��f_p���`ƫj;�!l�'%qwS��z�h�V�||��j�n�̽5�Q���F����⅕'P�'V(=��2~�yG-���?n,G1�9��� yqlH�!��'���X�8��[���#��s$[�=�^x�+�*ǅ��e�Q�(+����w��S��'P���������9|PK
    x�H%�k�^  �  4  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/COn.class  �      ^      �R�J�@=�Vcc�7ﶊoՂ���R|c#�۷m�)�i�i��Y�����Q�$�"BXfvΙ�;����7 ,$����!��Ü�����ax�r,����mI��nK�g³DӖ'A �E˷\�Pz���d��X�/�@h����@:��Bv�|s��P������,!�l�t4�y)[>��'Q���t�G������뻄5}��o��ߨ�L�>>ܻ���A�{�]��<��v��Ɓ��j�S{��Q��	��Q�j8,F���}ޢY���0��r�V�M�F��`�4�(�4�X1���Q��j1>@r�T~A��B���W��!̦��A����WQ�J��zF�7_����s�PK
    x�HHY��_  �  4  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/CoN.class  �      _      �R[KA���67�K�Ң7Kh�� ��hSɲ�m\gkuۭu��YAQ���GE�=D���9߅��Ϸw �����(�TLbIAVABA�0�k9��#DJn�Һk0��<��l~�B��r�*�L׻�m�jN�>��@h����!~_\�2� 
2q(H�C�͜K���pC��u�'��=B8��G.]�������i�^�\6u�V=�К�~�{�ݚܬ]��f�ߗ��]$��r|?j4+�eiF�5�0���ƣ?9�,Ƒ�4a3�r0�|
�d����%S��LVHHń���6B� ��'P��G9b��}/0+;�yĥ����Q�F#�zA�/_�嫒?-w�PK
    x�HL+Љ]  �  4  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/Con.class  �      ]      �R�N�P=�b��,�{|CH��#�������nI��Z*�g�h4>�~�q��cH��Lf�3�����|{���"XVŔ�I,)XU�P�$�훶�"�)	i�i�R���[����hx�c��k8nW6	��-�BO�}i{��r����K��(���8��!�vK+�۲�V�%�fϓ�t	�??�r<����������ՊEC�*��k��P�w:g�!�Jwй2j��/�<a/���Q=�X��Y�?��F(���8�Gӄ�`���#�`E�v%S�&�*��Q1���\� ��e�@�W�� �8�}70���<�<��3?�]��(5[�=�^��W�*󧹇/PK
    x�H}���Z  �  4  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/NUL.class  �      Z      �R[KA��Z���i����
�.�F�C�id7�m���\wk�,VP=��Q�Y�"�e�pΜ�2����;�M,$���������yi���9j��(����5��p�D���+O�BH��r|�H���%a�`^��0Ľ2dGz���A�¾�|F��hȧ�a���\�]���l(���D�i+�ɀ/���+_��u��n,ٶ�e�t�G��խu����֖v�u�<��C�P2ʧn��U��	����d3�`t	�ȶ��8�i̤�E��M9*��h Pf,��\�8>:��v���� ɕ'��+�<�\'����n
)"���}�J_��>�^����:�s��PK
    x�H=`�^�  �@  4  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/NUl.class  �@      �      �Y	|�O�[�� �P�-d��4��8۱�a�yl�dt`rM�6$�\� i��j���Hb��i�#��n7�n���{�M���W�B��f$���N~~�|��������_��2[���2���3�/&���?�|�ɿ3�.�c�&����L�a�/L��䟙|��?1��t���5	����vq�����:���D@�����!�M�1�4�,x�ɷ%��l|W�ϭ���cŷ% ��4�% ��i�/1y������L�L^gr�� �ט���&�Ę�cr���L�0y����$�!|�����y?��ON؂/�Y?fs~"��p-s���%��Z�E	�m���	;���ڹ��vr�k'\������s�n�Nn��	]ܾ焽���	��}�	~n� �?sB/�������?u�An�~j��	!?σw��}�	��K ~�����o�w��{�����ȸ?I�gn������,�+��g��KL��mL�L�P�p�$���\&yy�ıN�q���<��'bw'R��8	'����զ:�,�pw�KH����3$��ĳO9����e�{���H}�7i��T����F��4F#FP�&�+��2b�ݕQ��S�l�������]vM��iR*I�H�TF#�` 9Z����~]g���j}���Dc������.��/RVRz���˸x9�lCpT;U�BOЫ��)!��ǯ�2!Yd�/��?t>
��u���[�\](��(d��0�T��
o���0f�� 4k(`S�f�DX�P@sv��_@�z�a�9�PjNTM�5�&h{��V�s8�R��*H�2��� ��K�`�V�7�p����%��X�/�q.F�[	�d\�Ke\����Mjh�L�zD�d^YE&e*�U�Bƕ�J��L��\�b���p��p���qV�+�V�X�5��X�W˔�kd܌	����m��Mx-�f	[dlŭ2n��2��6&�2v�N�{2 U���`�r#�ux�����w󈊌{p��^��S��]��n���'�>ܯ������߫�r�����2���v;��$�� �$����e��~	d���7�,7��Mx����x+��x���v�`��~���KMƏb�ЄT��a����G�/Qj(#Q���@@[��o\����N�A�gX3i0�v���J��s_�b�Hq�!�[�T��0��"���`�r�BK*�j8yɟYfsi��)���A
\�6�g����ٸyi�F#>YE(���c�1�\W�g�/�Y��h�q^�bL��P[2�P�j��S(�a��W)\����!��˾C�V�9KܚN_Dc��^U0@����c1��Ծ�`H��F�L.aB�_�^S���a��t�0���FL�ߝ�K�{��f	o���t��y���|�<�Z�c�\7�j�-J�b���̰7ͩ���=d9⩩��o�C����J�y]z�Ԍ�MJH��U��!x\�dĤ�Ʒm��@�i��Ӕ�2�1L�̷���2HF�N!�\K�R�
M��6�VZ}}�u�+�b��n#TC�D���M~ū�%�\�h��FX豮W���)�v����)¶ݕ��x�Ks�1�:s�ih�����?�pia^�q%%
dև��{�����;D�D���#�n���\Q��u���n=�\�X>o�j(��&=u�*�������M�|���.����å�Wt�	O4�GG>�,2��F��/Á���'�f���Zz���$�K6�>:�Arz\O�3�W�Z��Aޜs	�����	��������66��j¦]��N�7�R$�����C�P�)"M���KH� �d=���7р��^�	���?�-��w�j�i��!�s�bY�'�5j�{�@wd�V\UJH�4�>�B0�U��J��p/]!4�Ծ���!�����A�U?��֠�?r�]�Y*>_ LU���U�M��x7~�_ޟ���F���:������Hh�:^�m�	��D�+~��}��?����s���7,�?�����|US�
���R{�5G ��3R�x���^.@�w��+�p�|�������F�������������.����~GY�@�����C�Ԯ����ۻڷ��Ue[���b��,�vPRS�B�^���F�gm݂m��������0y��cLN0y��q&�2y��i&�1y��CL�2���1&0y��I&���ge|^��x�y�&��(��2�
���<|�q6#��Y#ΐ8����<^���Pq�#�.�y�8�g��<e���qv+N��E��}5
ov
U��)([����1K�ٚ����P�&�5i�'�<diRE�yd%e�lg��i%����&.�u�]qUٖFE�aU�Yf����Y>��:gz����gz�ߴ��W6.-��$o�mZT�.�[�nua.�OǮOU�{�r���.��_�\Y���4mǼ�M�����ݚ�EzL��U�����2g��\�@���9�:��x�x����`��l�NM�0Qh�1&"U嚈���i"��D��H7c��H�D�f�����h��f2="��d��SLLѢn�j���d���[�}�nZUu]��/�V9Lɺ��Z�f!�t^�\�,�Z��6o]qϸI���ݟ�	P��`^&@�n�+`�w&@�>�B*��߸�_Z]^�k[l"=�K� ����V�UfzzV҅wB]h^��q%Krm���"׶�� �t�:�/W���u���p���=~�c[yo��5�蚼cl�!�a��@uɬ�e��sm�(��f�s�<���Lͷ�=�ڧ��n1����h��"��u�i�=��'��1�}ToO��q����|��u�Cz���>�������ޯ���-]�D{D���-,���{�ӴG���b��F�w�y���'�+D'i\|�_�� I�s]����u�>\����/Cة��ݶs�Y(�q���}������3�ar�y�b/¿����'�1�]�p���X�M|��Rj�<@t�Y��Eo�K۷�D&��iܞt����Xw wd���@>i�=�J�0�k%��[ܸ.gT������>s�\+�{�z��F8iTw���"+�?�t����m����yY�~�2��ے�ߖ�^5���#�9Vt5�-�p]�/��u��Ǩa�BRH�+"U�YN�4�T��T�I�٭����n����r�m#�۸Q�_���?f�y�0��QV�ב:P0*W�G�;0~������he�:1]�0��jW���w;��ܥ���$���޶��<��`�9(9$����مW��ɩ������V���pf� o
CV�3�Z���������Y�0�,\1*etҺ�#t`�8pĺE#t�xTxں#=BKFŁ�; �Ё���q�8G���Qp �ɻ�f��٥1�t�M枆)�nw�l�	���<;t���xv�vw4�W��ܭGfȭ��l_��b�p����c�P>Zd�m����²+
�R޸I��N�kH|�N�qw2��`Ps��� /¬6-%s5{��������-)�#�!�/5��:R�Ei�7�B�:�'�f'R����\���ն����Ŏ�6^��9-��+R�ڠ9��nN���\ �������G��ʗMth] �U��C'��'��ʽ�X"�y�5��{�O^�����Q6n�H.=a��C����P��%�`� ,�:���U��
cg�����Ym�1v�;���:cg������h�l2v*��Jc��ة6vj��Zc�N,ӫ��5`_��W��L��泰��͌x�rȶ���CC�r��7�P{MBr-�c�r�Ù���H�ʸ��2����#�6�m�U)��tIv0�M�V�pK�q$ig\���I�
�q$�ɸ�nm
W��#����%p�)�=G�݌Sn]
'��H��q^�[���HǑ��q��mHᖧ�H�Ÿn�ۘ�%~�L�H��q>�۔oz:�$��_�*R���8���#p�)\N:�$��*�+NǑ��q�:�+JǑ$ĸ��դp+�q$�0.*p�)��8�d\��եp��q$�g� �����<��Ay���������wKn-�z|.��+�{��_l��6�.�eM�l`�L���3pG�$�&��2Uf֪άU�Y�.����Z���2k�ӊ�G�p\�YmE��Vf�Z�Ykuf�5���f�*Ϭ�.��z�p��.*+��1b�+�݉+ J�p\Zb�q�ЊL�o:)��m����<�� �L���!-�Q2����ڌ�*�"}�7_Jr��ri�Y��l�uf�r�9��j�L 6��^iƬ5cV��Qg�d! ��̘��d�̀�G��X�<��r�{G���=K��ś��z��j��v�[{w|�/I����E�5b{~��E�r��/��u�~���d���\wNQ�t��N����������߷��'.]j
�o�����H��6|,4>;�F�nO>8�Gݱ>�*<��'�?s)�ݭMpr�e'0���o![������lU��NڣЂ߳{h��!4{�@�!�t ��E�v�d�����)P��J�`���q���8+����_��Y��W����)��ЁU��+�Q��M���S���?j/��8f=ycG���QI�i��Z�ǧ��ue+���u�X�=f���P]��PK
    x�H�+��]  �  4  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/Nul.class  �      ]      ���N�@����ZD��x�;��zYbLqa�@��0%��j)��e�Ѹ�|(�Ɛts��9�w�d�|���ú��b�b.�Y�J�IHHH��p	���愴j��y��5M~�B��\öj��m��ۄ���e#������\�ȗ{yi느�$���CB���U&�:J���-���T���-��yo~�c�6aG=���[��JEW�z��F��^�ܹӹ^�{׺v���J��,��#�烮�j�V�PO��8��G��`�C��AQ���)o�0VH�G�N�6#$�X�Q|� �(nY��wX�,#&��c���w��SɅ'P�Ὸ��ˢ=|PK
    x�H��-�_  �  4  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/Prn.class  �      _      ���N�@����ZD��x�;��zYbLqa�@��0%��j)��e�Ѹ�|(�Ɛtsf��;gf�|���ú��b�b.�Y�J�IHHH��p	���愴j��y��5M~�B��\öj��m��ۄ���e#������\�ȗ{���!;I !��!�Lfu�j��[.!�/��[�!��^�H�vmzZu��h������ɍ�=4F�޹s�s����u�ߗ�ʥY"P3 Vs,c��|�q�U��i�����2V�Hc���s0@���AQ���)o�0VH�G�N�6#$�X�Q|� �(NY��wX�]Ft ��0���
���O��+�q��E&.j�PK
    x�H��3^  �  4  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/aUX.class  �      ^      ���N�@����ZD��x�;��zYbLqa�@D�`J
��RA�D�q��P�)Ɛtsf��;gf�|��8���6"c!�y�K�H�I�f��p�	���ᄤj��Yg��Z&��!�ڮa[��3��VV�S��U��[�r2��z��N���&���BB���Lfu�r���.!�/�C�[�!�^�P�vmz^v�n4>�J%]5�����=4G���s�s�:��u���R�,��c���1�a��8�C'�}��8�U�E��"a�_g�x=���n��La��p������,��X#�f����8dS�,a��R�	>��~_h<��{�_��˿�,2QQ�PK
    x�Hx�8�`  �  4  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/aUx.class  �      `      ���N�@����ZD��x�;��zYbLqa�@DP�`J
��R�D�q��P�)Ɛts��9�w�d�|��8���6"c!�y�K�H�I�f��p�	���愤j��Yg���&��!�Z�a[����m�VV�!S��U��[�r2��zya�NHOHHG!!A�OT&�:J���-���T���-��Yo~�c�6aO=/���h������ٍ�=4��ޥs�s����u킏�J�f������0�w��԰nX�$�}��?9�U�E��"a��d�� l�!�'���Ya 	+�:;�YqFr��3��Gq#�"��;X�20�Rb	>��~_h<��{�_��˿�,*Q��PK
    x�Hb���_  �  4  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/auX.class  �      _      ���N�@����ZD��x�;��zYbLqa�@D�0%��j)��e�Ѹ�|(�Ɛtsf��;gf�|��8���6"c!�y�K�H�I�f�tSw�	���ᄤj��Qc��Z�r!�ڎn�nk�=��VV�1S��Q����r�IN�}a�FHOHHG!!A�{*��]����C������&�	���?Ե�������m�������Y]i>4����}�q�:��o���/*�k�@��O���.��Y�㼫rs4 �}���8�U�E��"a�_g�x?����~��La��������lD@��\#�zA�Q�����
��x���@��`��W%�@�W���/.�LT��PK
    x�H�d��`  �  4  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/aux.class  �      `      ���N�@����ZD��x�;��zYbLqa�@DQ�`J
��R.>��F���S4.�!��̙s������|{p�M!lD�B�X����'���BE��	I�n2���5L~�B�5]ö*��m��[����aC�����!�\�d"9���N���&���BB���Lf��r�Û.!�/�}�[�!���P�vmz^vw�k������٭�=ԇ��s�s��uot킏�J��,��c���1�a��:���Y�P�MO��(V�E��]����-,�0(��v
g��$�����gA����Ϡō ����`	��$K�	$��~�}��Tr�	�E�/.�ⲨDE_PK
    x�H|Tx�Y  �  4  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/cON.class  �      Y      �R�N�@=��JE�yb|CH��#����Qޖ�%��j���e�����Q�-�!i6���3'�{>>�����!�uQ,Șǚ�����$a���M��8NH��άsMֶ��	�{�c׸k8�w�y��FLacO�#n{��r����!; a#	)Br����U�v��!�/Q5���K������9�]�T��nZ|تVժ�N���Cs��7�q��h����R��ʄ�|P��G�b�Vb�Z`��G�~�v�MF+`KX'
aP2�k
G��qd̉�YQ�!$+<���?��q���%�a�� .����z	�	J.4�Ϡ����_�,���PK
    x�H���^  �  4  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/cOn.class  �      ^      �R]KQ=���f���Mo�Ж=AHѦ�w�]�������4VP=��QѬE�ra��sΜ{����� ��8bX�1�qcXа�aBC�0�c���%Ċ^]ҦW΅�mQu�Y��l�=����mY'�f̦�Ct�!;�U�^����� ���4��>�n�(W�����M�NIW��h&�kx�#l��euS�w�R�2���+�һ�Z'��%��v�uiU��C�(�;�v&,'УjH�Z�e1��jO�ˡu�8�9�'��$a#��p�	��AC`����@��a�������ĳO��+��\�g����l	D쁩z�>J�^�A/����|�����PK
    x�H�*�_  �  4  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/coN.class  �      _      ���N�@�����Z��4��e�11ą�Ea7��J���>��F���S4.�!����9�w�����|{��u�)�bN�,V%d$�$�	S�mz��H�isBRwZ̪1�dM�_��c-�t�
w���6a#�wِil�i|�mO;K��}a�FHOHH��� ��*������G������6w	��?�q<��������4J%C����k��P�z����jԻ2g����.�����S�1F���_5l������*���"�y�v��� �|l
E!��'���W!a	K";=vY!�*�z��У8dS�,`�R�	^���+4�J�=�����_\U��PK
    x�H�1��  *  4  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/con.class  *      �      �U[WU��d�a�P��z)IhH��K-��)! ��$�tH&��d�	��OY�>�]��&.q����(q�	�PX���a��ٗo��gf����?��"��>\ǀ� }xEn4eoK�/��w��!b����]�yOD�!��Rw՘n�7����0w���]���$��k�ź}:��Mݾ�0��2�p�A�[�����V���ih��0��u�l(���G���e|�["�e��*����f)�h��V4��1���NoC��j�:x0*c}2b�s&c�fkjg�m��K�KU�|����2�l�X�6�M��c��g�����!Z���\0[��e͠uW[��Nu�[���L۩�;�k�n�\a'��j�v,fZ���B(�c����a�XԪ"><Q�D\k���H�]�3t�4"��W�j� �B��eNB��V�$e��c^�	�L�qC��R$�[��yQeL���SĴ����SK��<h�Z��UH9��!&yN���n�4.D4��`��\m)��,�8�^�j�d$8����%��ㄌ$�;�@Ģ�%�(=_V�36A"���Y�A�������u�[��.�v�sJ��(P��e��v-��X��Nr~Ѯ�d�Z&�*&����F,s��no/W�-jŕ���z1����cy�$x�I�z��ԚA��j�hy(2�ƛ2�A7���8\��:��]��{s^����y��ك���?�b7I�N��vt�9#�V�GW����Kz�>xi��c�!�*-�k�Sa,��g-����E��&�&�
oó�ix�}�����F��nA��	��Tj\̮��9ezܝ�����h@���#B]��$�h��|
Gb$x&B�O;��)pO��u�%%����ĕ�deZ�7Td�%�E����������o��v�C�i{^�(�!��݂/)�dX�!:���&�(��k��������h���n�QW?z��&���ցۑ�H�ƻ��/ ����e2��=v����s�T�u�PK
    x�HQ<�^  �  4  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/nUL.class  �      ^      �R�J�@=�VccԶ���V-��A�blŻ}۶��&�V?KP� ?J�D�AD���9sv��������4R��чaC��0�aDC�п�x��"��~Sr���Qw�q#���;����$,�K���)Sv�������S�� s4d	��
�eV뗲��-�FIO�d>��j��'�Y{Uu{U�7�JŶܣ��s�v�m��k[�G�^�̮�˻�Y9qK��|\N�G��bމ�b$��]��Uc���cS�6��(a5��x�	��A}`��2�P���`�����֑��WA�$� �9N|50��l"���7��d��W.
O�g$~�����Q��PK
    x�H1�2��    4  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/nUl.class        �      ���NA��Qv�E)��*Z�E/�M/����HK��f�Y����e�5�41մ�Їj��`L�dϞ9��ٙ�������&�xb`;I��X@J�g�<'�\��s�5�H^�A�$ZԫQߥM�}Q� *x��S�Âb� ��-��!�=�;v5�]��'�	���V`!��*^XX�K5M[��$��D{�1���!���Az��
��<�EU�֌���.�H���UF�P�1���c�:�P_�������}M@(����J08k�~�\vJ^��xb7���n����0������4ٯ�Ϳz�K5�z}fa��͇������]��lg��F$A��	��ѽ��H��B}�~���׈�@��J�	,��Yl ���|v��ϴ�x+�|�5=�s���)B�Xh�5!����� �PK
    x�H�J	�^  �  4  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/nuL.class  �      ^      �R[KA���67�[����ڲG#�!�T�,}uVV���]�~VP=��QѬE�2p8g�wa�����@���!#��X����'���B%��	I�j3��l��~�B��]�2���,{�;����c#�����7]�x9���N������BB���fv�J���.!�/Q����&��~�k�aO=����&w�岦����|h����N�Zm0�_k�s~_R�WF�p����������!�6��*���r�X�"�aן�?�x
�E������HV@HƜ���>� ��(���Q��X&�
�B�D�'(9��?�^�˗����_PK
    x�H��^  �  4  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/nul.class  �      ^      �R�JQ]�K���{Z�f
M٣��M*Y������35�Z�E}@����a8�ٗ��b����;�6#aCF2�.!#!&!N�9�M�9"�JV����fF��:k���k;�eV��Y��w[Y���LaG�cn:ʱ9q��N������BB��P3�J���m������C���&���P�r,zVqF�M>l�˚jԪ�7J�1��/�;�k����5��}I)_E�A�/�գ�O1s�#�5�bⰊo���*֢H"E����A��ma�0�a@�)��1'����G@< �{�_|!"��� K"��� *�0�������s��3���|��/~J��PK
    x�H���\_  �  4  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/prn.class  �      _      �R�J�P=Ӈ���Z��*�j��R��c[��fw���ؘh�~��(.� ?J�Tq!R�y�3����Ϸw XL �q��ż�����4ah�r,�+�-I��nSا³DÖ�A �Dӷ\�*=���d����/EOh���dO:��ۇ����)!;� ���qB������*�K��	������#=B4쏵]�%����ڐ]�\6u�V�?׌�z��9�nLi֮�:g�q(�KZ���"l��r=j���#A�w/\�����I�b.�&��6�#�)Xf�����MvV��b���\�#�H�@�WD� $8N0��������?�D�(�P/>�^��W�*�'x�/PK
    x�H��ؤG  B    _020_/resource/1.png  B      G      B���PNG

   IHDR           szz�   sBIT|d�   	pHYs  �  ��o�d   tEXtCreation Time 08/02/08���   tEXtSoftware Adobe FireworksO�N  �IDATX�ŗ{�^E�3����Wwi����k�-B� (���%����Qj��?$�$�!��`���"�(T�HP�啲�[��v��~���9�q�v�P|�IN�w�;�wΜsfF�ds�ϟڠN\r���]=�8��k���g^���+�����"�_ ��<�˵j��/�qa�7�z?�����]�EL��[&n���Ķ�؎Ƕ=���O�þ�_��T���?�������h�)t�րM��`#�0����'w15��������g= o�G �_V<b�g/��{��ÝR@9��d !�6H��k�	���6\}�_\��m��/�-�-9qņ��-���� � 8Ep��X<�N�;�g��-�~云[���+:Vy��[�CG�~:�S ��"���r�� ��u�����x��y���=������(UXy���V[] Q��T�en�լ/ ���oS�Q�<�@w��[��#��h������˷�����U˱��V�|�^�-���3�.I� ���}p�`]*��z�إw�#��V��V��J�K *}�Pnj�ʖ�� ��Y�e�Yl�6$� ��x�iH�i� T��k����ƃ~�	������lh�R��P� J�E:��H�f ��m설�C���Ю���*���C�mP���Za���׉�~� ա���`���%I�\��C}�E��q����[�uf�$��P�?���j����~�G�wN�W�CX� 7�ٷ}�$,��Wٵ�>�����:h��5�x�ѭ�=�ߧX-c������C:�� ����V�?\>	�X|��g��S�D�x`B\'O��uP�N��+O�aϳ�y�b��4�TB0���מc��g��@4q�i�5	&D�A�A+��y���+�5Z�����
Q�q=-�����
,^.��T�	@"�	8��6ԧ�4��K�Hlb�ƀX��y �Q���.��js@��IK�@ir�rjaV��r�f*6�[��F�I�dN���q4�	R8��*���4וs�(��mgd����q&I�Mblb�y A����Z�;��3�bY6H��
Ӂ���X4g�i�b����D�(�D�}L%oΫc�㿏ۍ:d�4���R�i/u��[�:H��F&u�6&�Sn�8�h5��y��{���sf^+�V�!�"���V�~	P:-L���lG$�Jb�%%%C|�Ąa�"y�e�é "bG~���΅]�_GO��˜M��+�a�Ji�R(�瞵�׫�r|�=~5N�w���6�բ�|��W*U "1.���;{��|�:�=BCeQ���LG�*��2X�_}� g s[�����vܩ?a�S56����+������M0�v��N����i�g7��w���V}~�ϾQJ1�@��*?q)��G�c�$hC�blW��Q7�3��@Ý��hō�ݚ?�С��$�(tV�����|��P�4b�;�kt�<�?n�0��8ɓ��HҬ�r��u 
��}�z@)� �k�W'\sɲ_w/�̉r��y�m��6�/�)VP&LS0KV��U�&(l���ԣ�I�5lc��^�ɗ��+��Y.��N�f � n9���y�>�={
�w��$A�}�"��WV ~'(%1N2C��2��f�d�hL��mw��^m�t�]r3ГU��ּ3�R������Xsن�[.]x�ӱr]���Ib�#QD{8$��#&���f���mm�}����E�\Ң�^�z(�<�	8���W_)~uh��j���[@zQ^	�\P:=A�6�=E2�����۱�����a��
� j"��{�JI\�~~����۸xq�i���A�����*.�����&jL�Z�{vL������ox��i-Gmy��z��S����TN]��Oˬю�#ƴ�@����.x�GB��������4p��q��P�j    IEND�B`�PK
    x�H[���w	  r	    _020_/resource/10.png  r	      w	      r	���PNG

   IHDR           szz�   sBIT|d�   	pHYs  �  ��o�d   tEXtCreation Time 08/02/08���   tEXtSoftware Adobe FireworksO�N  �IDATX�ŗy�U��?�.�ݷ��f��AP@E�B@+�[-*����(ZZ�1m3�j�6%iԸUMk���jI�J#jEpAa�q��a�af�����v���U�ƪ��I~���9�����9���	�_�0���b�sg,��M������qrv��c��m=/�mQJ��.���l��o}���铖D�N5�2����|���I/���=���m���'����� 	am\��U.8뻉��G�D�K�>H�[4�ː;�C�CO���?�P���`[Itƴ�~�rᗦbEA
:(d�w�˃$L�mmx�Owo�uʹ��>@����?��[��bS���6TTC(V��@8�xaތB�bU0i�e�U���>+q��s�|A����Ry|ZӍ�o��?;��Q�l��[߄���!Np��i�aA����l��`7�HbMkb⒦{��]��3n"2��˞-�5-���VU ��W����=P7��UR��#��#G���U���|�U�k'�^��0�	�V�� �]�����M�H c3s�
nx�N"*�ŗ3�A'T��pBѢ�D�x�<�]���q�#w�����0&��r��'<�/6z]�ܦ�x�p�cQ��yHr�o7Ѹ�2�{��aHT��3���W6Sr�\�zn3�y�lmE� �-��(m,���ɥK?�t,�w�ī�.�P^���6�+�r�ZbŅ�n�ȇO?���GWy�B8`k��d��\|�m�4�qz�aƇ�C�Q#}�|���ݯ��C�QBh���}]DC�jp��~8�������v�ZZZZ��ng�_�k�܅ҁ�A���U��︍]�v�l�2֬Y����/g�h����"��s��a��X`U%� %h������d3iZZZ�������˗s�%�P>n<#��tN��J�����w����y��ǹr�
*�T �O�|�"�Ku���GԝV�Ĉ�	<�O��Ī�9t��{�1�����j^��2
?g�R���J�H��c}�mmexh�h,ξ}��P����%%�V�y�(�HU�]W�n�PD��>���O����5�W����Mk��Axit͇�f���lcFc-��&��y^j�;��v3��/	�$�I�(5���'�8fy�}���<s�=l��V*�圳�\F�� J�s1a���x��뾹������z�y�Q����|�/A��( 鸃�s�-:�&�1��7���o`ɜi�K2�o�F,��e�QR�o����$*Pdv�L��m4?��%��x~����(�|_�����c��[��� {� �a�X�(���*(����.e�~���~D�sn%��"]��s�?���ڻyR*��P2VF�@)PZ(B�$� ]\��U AQ�}|���́́t@J�� ��q	\?��F�
ƅn�m�w��h}�,�,H<�?��常+(E ��g�pAf���������vՎCr���RA���ϕM.��E���tt��\ӏ��x�	��.�bh�!���*0,���H�&������+�_/��J�@x�Ń��z6�p�f�O��#��ɀ��w���i�&?�V�?~/�E�r玃;d�s��`q�B��%Ju�ͯ�7ZZ��"h�_�J3��2��+#ˀ�M�N����L���KM�m�]t\��N��nwߪ!�j

p !��'��/�?���w4�D�:�0�oX�K6@�`�Q����O����s��]��mB���ڇn�x�<�u��8���� ���fQ�PJ!�Ѐ��s�/o�S��2+@G[hV� L���z�w`W4�}%s�z~ጠ�,ұ�l�����=��}�A�����@�R�� @��R��˾2���)��rD8V Y(-��r��Q¥�y�T2(�t;���rY��>�]��;w�7��ϋεb�{�R�QU�B/~�Y�U��Y�4v�>��20-�B�� 4��@�� ��(�%p��0�������;�i�r�'��0(��O,ˋ�(�$T>�]7ez��D�8�3��,��	BG) �(�&H�w$w� ]mG�<�����V<�Y ��r>W_ 
$ ����X��6T\[9�L&K�XB�4��� ����`.w����c����~��#�է�_�s7�~�8�1��rfj�Q�2猨}=}l[������������^H�H�    IEND�B`�PK
    x�H#o���  �    _020_/resource/11.png  �      �      �X��PNG

   IHDR           szz�   sBIT|d�   	pHYs  �  ��o�d   tEXtCreation Time 08/02/08���   tEXtSoftware Adobe FireworksO�N  IDATX�ŗi�^U��n�>�0e��t�����C�B!D
�1� !FC$c�_PH�cL��AæY(��.1�ah�Li;���y�����N�#��%������=��=���y�0��q^�ɼ�ԥ����..vv�e;n���֪�&��_��@�1&<Y ��xdP,>�\�ֿ�BG�n��f;�#�����*�g�au�@������������� [�����K��Zַ*���|�h	:����`L���gf�ۏ�����>��y�?�㵥�/���5Ck�R;(�N0`T�
�$ ,�+���ߨ���sÆ;F9)�Wn^z��/^�L۪��ၕ��@�ޫ���g�)�p�4�#��ed�[��z��	����CW}O��O�^�Q� V,w��>�f:�.��F��D� <��w^�s���|�5�p���m���u�@	X^jx�3���l,�`sp�t�=V
뵃� ߽������t���C�q�wv�Z�78�.�[Ɍ�)�eʘT�H��.���R9��:�������m���5�n��%0"(ۃ\	�bv1U�.����IoD*����������������uh�m��>0�ۺ�rw�K�dm���D�wp[z)-?;�\�Y�S$Y��H&FiN�a�6��2�]9�Q
�����~3�Sk��wv�1x6��"Out��ZG+AT���E�~��5[ ��@6A���p�C/?F0y�|���Y8����@�c��7�=:i�<��ʭ�����/;��[*��
,�@ұb-��T�Z��OO2��)\WPZ��&��Dɀ�=���h	�>�L I��x��s���,3?C+��Xb�i��� ����˜�]AŠ,��P?��x%��[�F��o_�F3�&B�'9e��k7B؄f�:�9X��uFK�RX��b��R�-c��4�T������`�[yV��sY;/?a"����$x�\��|j�	�p�t�]��Z�h�Q�6} l[t�vA��l �V��V/��N�h�/lzK(e
�B�~���1(I�i��$���T��- PI<mTd0�H[�3��*VV�����yMH�\'�8IRoU��ҸPa
a"P%:I�R΍��`vv����v�`�o1�U���0�6�eN��q�P*�YJ�a���9S¨Ũ8F�12N��<� ~}�i���p>��f��TB�*/���I���5�f=�8��fU<o\'	2�	�dA�`m}L�V�o����>\�7�,�|�E��Q�uP�`f�:p��LE�0J�(F�q�]�j����/��3W�iyŬ���k�p�q@�M5�6[I(cp&����Y*-�(?@�!�����|Ə6�2pW�)m��1�x�O#u�u~�u��d�`h/�&�6iSs7㜺�B�2Z
E,K��!���=Oe�)*^�8�0D*�QD�����! 䀺":���{�iC�7�����bLL�a_EkK���9I-Ba��؏ʯ�V��o?"7�%d��@�st,|c�=�� f�� ��l���?�m�[��'-�1�� ^�z
���ѱ�+0cF��x'&�N)�G��Y���ۅ�bLѬE���������l��0� ���ҭ��t�˟h?�-���(�����N%�����J��H��	:��a�(�9�Wtc��^����;W<l���}G�1�\C���=���#O�^=92�(F��$d�C�2q���J\d�"��TJy(�LEUm�	{���`���?f�I�B���f�����g�Uvk/�m������4ccR�̖"BUT�]f��6w�Y���Gy83n�05g�}M���;����7�^�sM�%y�u	"�N)]
ac�&	��rf|?�}��/Dwo�a�4�YcL���"%q u�鬻���zw^Tj�Z�:Z�\��v��
5UҘ��걑���;�����E^�<͇���Ny��p�J.*��l�Sk�G�yc�(/}�	����φ����c��r�H."�i    IEND�B`�PK
    x�Hw�B	  =	    _020_/resource/12.png  =	      B	      =	���PNG

   IHDR           szz�   sBIT|d�   	pHYs  �  ��o�d   tEXtCreation Time 08/02/08���   tEXtSoftware Adobe FireworksO�N  �IDATX�ŗy�U��?�.ｙyo�a�aG�e�`�R��T��5V���RjJ��&M�?j;֚����J]���kmc�B�0VQ���0ì��{ﾻ��܇8���%���$'���9�����9��gٜ�Y�����&]<��ʆ�E��6jx�Hvo���//�m1��g �]�l�>���k'�seE}�L����v,G���!:�T��~v�H�ı��n��Ē��=�5�R!R=x��ƹ���;��J�Z���#�!��&��S>�L�o��y�������U��^���f�Uu�;��Qe� T	L�l�"��Ƚ�n����[��~� v�>�YW������U��XI��*�x����sv%8�.y��]t���?8r��x����7��i[X�N@eC,��DTP�A,���&���
l�z <���ɡ?w�2g��p�w����4�w�T�4�)�cx�È�J�g.&�8��8��" w`'��&C2	M�'P5~2d����]���v�/����e������鳧b��8�}Q���ťTf���~�o���3Jd&�o l�~�9��9����ڦ���Opx�K4�As[\2c�s�0�a`�?X /\c�k�1�6+U��]]�3���%Wӵ�-6=�num�Vs�����:���#U�h_�����S�ɕ"�-��a��B�>�`�i�Y�ug�5�`��V���\�Be��Sә6w!�6m���KGGsf��dO7-�L��$�ù��K�g׮����լ_��ٳf�u�V��9���^�R$*4M���c B��u�r�H����j�B���Ge͚5�\����~6n|���1�VbFN�dƒt-6lx��˗�v�Z�(bݺu$lp꧃���Td��r��2*�\�,IUg��
��q�$,0ưj�*�0`ʔ�[7�@Xl+N�T*EGGcǎ���%^�
4h�qK��������ƵO��I�T2��T�=��ܰ�����"�V��ߺ��`n�K���q��w���@gg'����g�ߏ@*x��Q
���T�;T*���e,t���i������2�*vwu��{Tg*�fGHȣ؎��al���/Q;�:��{7=�>`���(�;�u���� ��m3a�m�zA$PA =�T������R���N�����^�R����-u}�=NP����F���ۨ�oFJ��)1J�1�Q *
��
�(�\�SA�{
�A�)�-Hq�L��@]�&�7���V� �q�i��:��R��Q �\�K���v��ˆ�*{@��Q3ұ�6$!�ئ�c�.šBT��F�P��*��o�zAz�<�?s��"�"���G���"P��⵪��*;��Q�qEH?��E��
β��k��f߫l�^�Q`�vkG��`��:D%�B����²$ɤ­�����X� ����0 ,�f�~�k�G�1�����׶�-��^Y������4H_�U߂�T���*G��J:�p��h�����>:ȏ�o�~�C��H�1F; ��u?�0�a]�x�E��ul?��%����������I����83��B����~Gf�14җB�  ,��:=��$�B����֟O[0i�]Y��`YH��Ը�tF"�^�Ro| @���� ي��
�\�}�'?��#���q�������e�
������Ԇɻ'Lo�`,���"v�C�ԁS�b�a�1J�e���ho ҳ�:��� �8�덯����F��K�~c̈u�:!x����3���k�#,�0�r��ԣu-m��Q�FI'�(�FŸ́��D5&�E�]��޳��eqȸ�No4��o��|��M��%���BF)d ����d�"�H�@�J%P:5�h���uX������@cY/��1Ѩ+���yׅ��\>��[��5��ւ�B؉���i�)���q��R5|���c�]�F���Sl.�`<-��K������*״�5�Ȍ�rj�#R��T��/l���D>�4���;u��='���������"�3���] bP����.K]�:�Ც��6����NfllW��AQE�!���u���o߾���W�Q�1�o>��%��q����ҩ�pYU���4h���d��=�k_{�=c������Y|���d��c���    IEND�B`�PK
    x�H��Z�{	  v	    _020_/resource/13.png  v	      {	      v	���PNG

   IHDR           szz�   sBIT|d�   	pHYs  �  ��o�d   tEXtCreation Time 08/02/08���   tEXtSoftware Adobe FireworksO�N  �IDATX�ŗ{�T��?��;w����vaU��A�J��D+�"���ք��Ѥ�Xb��Rk���ML۔�F�T�MlĠ�B�H��*�V\D\���>ffg�޹�sN��E�&��G�%���qs���=��{c�������5]���tK�+kב����߆����'jی1��N�����oｵ���Kɖ�'�l�l�hat�]�c�Zq�xy���S��|������5��B$�=��ö+|�a�Ld J��@�����	 ��R�?���?�r����������]�rճ-��ͲR-� a�0`�8�ګ?	X "�;y�?��/w_v��'.`���Kgy���y	L�2��8@4}"�Εjc����O��N���ȥ�����xmu��?u�7_o�1�Aِh']�U;�F�r��5�=���p�MSK��+zz���^�_������G��M4|}��[�\=�@�w�G�E�yr'�s�V���k�}۟�m[LsϵH�f��!bb��N�:A��7xkǡşy���	p|�}��n�SĲ�l�r�ǎi���dC��w�Ӡ���p�cU!q���(d�a��7���N9B��I�v(������꛵���� `�m���3g�!��	<Μ,�u�.�>�\{+=�n$l�r�8�����C�&��ߵk}}}8�f͢�]D4: ����p�wj��?+ f^��;Sm9A�e��It-"�qX�~=K�,���c�Ux�_OD;�;�'�5��^��5k�0g�֭[�# ӵ ׋��X¡�3{�!����H4uNY&lЀ!�4m�ٵk7`���<���ٳ�l�d��B�!m����/P(ظq#===�]��|~���)kb�!��u��.{��R|�]��Lz:Z�P`�T��F.�c�֭lٲ����eՓ�(��:Ĳm�oߎ�������!1[����c��)��}�+��1�&˱��r�G���bT���l�L�z�)V�X��m۸����/�0(�H�)�;�-7�`�lڴ�r��c�=F���Zy���R@<aϝ���I^��@���tA��&����Υ�����^ 
�~��Dt�ӘF����K/����ihh���7�Z�u�:C�B8&BZ�c@`�-�*�Q���d�$�YR��1l�"cm�p�Fq���XD���䏽�����s��U}�sſ�6��Ji: �C:>���J�'��������E]�12Q�tԅ-b��{A����^�M�?��<a{��=�0(ޥ M�Vhbi5�خ[}#
���v �R�.Y��-��""�5��!L�����~Or���)ǆ�9L�.q�D�����QD"& ��_�u���N��*�,��5�S�*��D�6��8Q��[�	@���*�)ʱ"�Q>��`,�XD�¯E�&ԁg^�m�U�D��d�D
��}�SA9E*�9J��9����AT���@T��1��j�Pq
��ī�N���h��&�wO x�mSK���I�!9��B�'���2�/�Dz��8���0���(5����!����084{��)L9<u�f
!�b�"J��g�vM�J�%q�8�w@Y ��P@3
��Vw�qѦ�%"�����x�W�^��Rȩ��oFk�@#B૿��y��鮆�7,M��e�C�X�Da�s}(� ,�mK&7k3(&2�`|2�@zL�.
:�r8<��o�F���� ����rk|�Y6sV��1�"�ii��IR2�БS$u���#�$�zx�1d��`�V����SR�+�C��|��7�}'\J@Ӹ�����R/���ڴ���d���)I�R��O���1��hF`	t�H��e�
eܠ�W
!��r�O�䖧ͣ�ы���c��  9�<q�s}����Φx�N#�	l+�%R�d�:���1�B�(�L�0��|ta}f���Tq���R� o��L����!D_�U��N�y{���i
�iD�$R$@�����5Z�h�����GNS>}28�7���͆��*����T4a(u)���	�Mw��qinUCnj��NE$��é��''Fkkho��xw�=Νع�U�G?�+��
��1�����Ā�ۗs�W'n��h]�nj�K7g�D��t��
�:���^1r$?�{�[�����L�g>b���n^"_���T���e�i�<�3o���{����1#�����m�O��d*����e    IEND�B`�PK
    x�H��i6	  1	    _020_/resource/14.png  1	      6	      1	���PNG

   IHDR           szz�   sBIT|d�   	pHYs  �  ��o�d   tEXtCreation Time 08/02/08���   tEXtSoftware Adobe FireworksO�N  �IDATX�ŗ{�U���}ι����0/`�aFdD:�����5il#�&jQS5�B��Wm4�!���U�M�i�����E��Ed�afd�a^w��<���vjk�����s���Y�^k�[c�2�s>�_�A\�vե�V��-��X�����sG��q��h�1�?_ ��"�B�h��}��:�m�T]�űT�4۱�F���U�;Y�s��w�����տ����"�ԓ�?ܰh�����*+�hZ��@�`B0>�qǆ�8��r�o�<��WM����K�|��u�,��u� a�0`T  偉@X���ɓ�}���҇�^8/���Z�/���oL��3M��@[���0,;6��z�*�����3.�N��ｮ���g_`睙K�����5󗦰S�:����h�dk34/]�S=�|�� ���ȍ� ,�ghZ8�)��{9�{���<<��s"�жj\|�����y�=��ū�%���{�b����4@��c�1����Mߤ��J�|o7�ѝ�[Ҋz(?���~��[Ã�r���7~RQ��$G��x|1�+�:^���Dߌ9|���W�����'��@����� Q���n��P+����d��Z�/o{��?X ��d77.��J�!�83"i�l5�qc�����6�Ё;< �,2w�����e+�ͮ]����!iA[�b��N��0��Q�������)@�u_�=��Ci��q���������Ú5kظq#���s�NZ,��C��)��!��I��sϽ�[����6o�L҆��x�I�*Nc[�� !��Y�7�x�AF!�L6�e��-[�c�=F�XdÆ$��XNt��B�/�ŗ^&�n���ٳY�v-�b�L}3ƪ*��l���7������:W'���hBb	*  ��e��̙@mm- v<��B��X�Ŷm�Ð��A��8 �Z���q,�</�8נ���٫���E��B��"� T�~�z���صk,`ӦMx�Gܑ�IeL�>���7�h�"�{�9�(�'� �I�����h0Ja	H�b_��Tu�Ӷ��A�d�*1���3g6���E?---X���P/�N	M��
FO����ر���n���hkk��S�3��DI�V
�¶�=�l[�	"�
��%
�k�S;/H�2���"���X��]Y5r'ޥ@ggg�y �x���ZJ�����Ĕ�(7*0_�l��������י�[���2OF%)�A�sgA"��!��|o�W�a9X�qjF��V#(	:��R�}S ���n�Wى�]ޕB�K��G��)���B�r�2�| U �)C2؆<� q�~�.F[��C�!:�a������`�u�
���U�lQT�C��F�"Hdd��Y��-ǌ��!0�A��9�:��~��FS��u�K�?�;�v+ n���DVr.�@Ax��eUQ���
|��� ��0 �B���`�ѹ��W�[��s�O-ʃp�&�8��q�n��rQ���<��-��A@!��M�!�B�\+�pw�3��񨜆bee�՝�h(��p���qlw7:�(C�r���\��� t�|�>���@�	!>=��<:kӼ%m�U),'V�S1����OMҸ�Y�Ռ��@��&��}�(���H��e�x����
@L E@���9u���\d���K����1/Oz޵$��˭��
�i��}�dCE2�H����|�_��?�,�, V�"�:[�!���'��;�k�%,�� ��,�h퐬��r�%�Yd`�d�ʦU��H�|���?��}@�",%���@��������6�7� D�62����m��`��� �d"C�4J�Q�ڤ@7�����-ϛ_!p�M�dB��Wй���g�6]d�̂�4p�;F!2mX�Pc�Ac���V�^5���P����������cg�F�
! �v4�|���3n�NoI:5-�d��ee������G{cȉ>��������O��Jŗ�IcL����L� ���tܲ2��Y��+���c�;���c�h�J**��n�L���={��۰�����s�_�|.��Y!V̙��t�%���k���3�O���Wx�5&�?����ŗ<��]�v�o�     IEND�B`�PK
    x�H�5>/	  
	    _020_/resource/15.png  
	      	      
	���PNG

   IHDR           szz�   	pHYs   H   H F�k>   	vpAg         ����   bKGD � � �����  3IDATX��W{PT�>�.��_$1����g����ѤCb����?G�H�I}��hښ�I����:1�64���dQP@E@@P7�򆅕��XVޏ��;�^M���Qf������}���8g��?��is$O �%����(�GE���bm�j�Z�At(��@����t�X*"������{(7�����w
4��_�k@�#��Dw�0x�#P�OQ
r�	�@��o%����FU��z�w�Ռ���h'z	�! �i���O��9M(ݦJ!�^�(&�7��b��m�>�n=�ƕ�f n_�:��%�?	H�&^$^!��m���LM+��?�B�&2��l�{Z�jh�Y�g��J��u"�WD��XA,ez�ѭ�@W ��+�~��7��l��{�iy��К��<;HBL���SFO! �}��q-��ߣ�z�����	#Ux¸֣�9[/Ү�'�sw%=T�چp_h��9�B�}�)x�x�}�ŧL�)h-{�S��*,81PE�0��u<q�șC�J�w��N�<�Q �}O�VV�)?h������c.\?F��!H���b�/sþA0	�����ǉX"�H�U������+Oq}�w)tH��c����̱�	i�7��B���l�?
��Is�8�����|�귭@$ߓk�~*�cTO2P-{M�(�ͦ��C�1w��
�s�RF$7=a�J+��U��Y�̌J��̱��Q�u�|�G�(���v��|���Y���p	8�����PU����KD��g��A*l�i�#*�`T�F2lI�AU�$P�5XE�x5s\]�;�E�}�hYٺ�D�@�)!�C�M�u!�?����CC�1"��g�K'�p0��S�y�0l�g#�F���H8WYP���=�؞���=��^uD%]�������������6q����*�H|JZjQ�;JE�4��)��������z>Ѧ�Ņ>�h~�0�"�cN�#���i�������ޭ�f��'��=Uo#i}>__�����}��Ŝ�͏#�cZ�a
�b�Jgdѵ�"G-k��5��MO��{������yҽ����*
Ʃ�|FA�[����,h����զ�n�ġ`��A���(4�/1D��r\S��s��7L�d��\��� $���,�T��|IƱ[�0z�V`���>k��O�((��`�O���hI_cD,�]�P'�*4��c<M�V$��)u~�O��a"�8A��Y��A���N�E���H�3���pb�1H���QN�(�p����h�� �i7����y%�~$�ǈ����33�45[2�"&�-�*�g���$+7_��(T�����o��r�(���fy�1�'o9m�����/��,#�����X|6mWy�^�g����i*0�g���v��)vYw���s��jr�mE/G�ׁ�ժ��"���ž�Zl˭Dx�r ����D�b��L���E"��e��@�b:ͻ���8xLN�B�-\A�������a;<"����q�Eg/�;Ĩ�D"�H!RMA���{�uLm�l�~��q���؊?�8p���,r�7�EX��������aѫ����CęEz�H0Du2�ʝy�!��Ky���VҨw�����(��J�m8�h��g�x��U8�1��jhS��m��4��|�/ZO�˔�6$#��_��ߘ����$ٱ8%��q���(ڿ��ěG>A	۩��\��ul1�_�7B����b�D��0�m��k�e�tOw�)[���-�FQs;rݭHw� �7�`J��PO��W�;��|�#��Xx�^477�09\�z�|ϗхI�:W{�ݨ�v�R�u���E�U�������O'��ݕ"�v��t:a;���p1=��@��+��*�(%���ٍ��^T�v��؊?_�@$�!�]kBЩ�벒��YT1yN��ݰ߄�]S�
7��%��g�j!��[`��G�)�ͨ"y1Ӑ]�Żl�]�j]�g�u��Y\|��h���*^�&��`~�&�}��y���D;I\��c�U�XӮ�����ִL����>r(6�w�%��\;����$ٿsE�*U   %tEXtdate:create 2010-02-10T02:38:05-06:00���   %tEXtdate:modify 2004-08-29T12:30:22-05:00��*|    IEND�B`�PK
    x�HD3��  �    _020_/resource/16.png  �      �      �#��PNG

   IHDR           szz�   	pHYs   H   H F�k>   	vpAg         ����   bKGD � � �����  IDATX��W{l[��}��3~$��vk�PF6B�� Z��0m���4�v��!h�V:F�[��	��!MEc�@����@�2#yl��	�BI��q�8�����vε�����?�IG����w~��9���XG���4͓����"U�s�E����������5���7���/�r��T*����b����T鞢מ I^ I� '�r��7���  �L&TU���,����F�111��1��H��� ��]!��d�d���ݺu�566^YWW���*TVV����n��l.��2�l6���>n+:�7����2���W���t����x-\��kkku��|(++��b�B7N�G&����f��vm�-]�`c���~:�S���� �H���a�ʕ��x;e �}g �
^�
�0��#�뭓p߱K�Q��1\���I�W���K!��9�D<]�������$�DI���4Iyt۰�?�tg��{�v��ID�	�~. ʂ�,��{l�&��(z��{~������xw�z��<h�P�	�sOr߱���:�����N��(9f:�,�9��~�S�x��O�lYE��䎉���Ԓ@<�I)��������v�pl�X�z��0(�'''A��,�>:�X�Y�_��$�@4��G?�й"��ܲ!�s�!���z��6�zοA���á8������S
�:*k���z��W��։�l��4j�K�C�`8�nf<{lD��R{>��aE�,C|�s0�*p������M�w���Mg ��B,����=dcl<�N�^2  �u�`��uM�2���gض/��v/Y��3��nl�<����J �\�[�g�ሦG����r��l%P��,RJ�;2W8]��P(�+�E���9�!�i��/J�_rô����F����O������Z��3�s��g��z�E��:ṱ�N�D�>��HB�%�����}X�G��K�n�����JC����4�蓋@08*,F�0� ���a�js�ywM�ٴ��� $:#�h|��==f^4���$��a���c���Q���Eyy9***�!e���j�*����;I9�!���n;E���As@9��1�عEb�%�� ��4�K X ������44�p���(r�4`sZ�x%
���Qc��L饚�8!��H�X/�̘$�B�/�V]�;�p����Z8�GA��D6{�������e��P�"���(p��wq�h�ڍI������Ι��k���hx7��K�Ih�
޹�=ak�?�͌k��c�)�n!+��2E�DA%�ͤ1)&y�YU�P�YC 6,�(5�cCf����p�B���mVP�Z/��&�ǭ����Bc�Y�5�xsT�E����0�~�=M�O�C|s��p`c.'��L���7�}] )�~� ��+�~	a)�36n: C���d�#k�������R�|��c�g�a�V���Nb�Gj�4k�UH���x����lQ��%�~zx��~�-MCvll�2|�F����a' *�в\�^婲w��W3{ļ�ƾ�ۅyׁ����!D�<�o��hD��]��#�u]�,����H�X(2
A5{����U�F�Q)%\a9M�R�$a�C����c�pS%��7Q
����t�f�݉᧷)2<r\R���DBƚ�e��G�"]�Ydl���O�R@��|�^���a�7"�J-���
)x��{q�5_�B��v�8��6H��ƞ|�K��<���$��VбpFd^���O�t����=}��A�M7�_,���m�n�ȥf��Eh�
�~�8�)|��e��/��Xn*����7q��i�]�E� 9���&�n|�q ��A�-+r��]h�����p�g��ţ�&�pU�a�=��8�?��]��}�8(�0E�f(T�V*3���vgq�s9Jhf&4��<�T�@V-�g7�"�FJ��J ؒ�#5��+��ͿAۉ��G����}m'U�-������v��h7~�ء�0�׿\C�܋�   %tEXtdate:create 2010-02-10T02:38:05-06:00���   %tEXtdate:modify 2004-08-29T12:30:24-05:00�LF    IEND�B`�PK
    x�H�d���  �    _020_/resource/17.png  �      �      �O��PNG

   IHDR           szz�   	pHYs   H   H F�k>   	vpAg         ����   bKGD � � �����  �IDATX��W{PT�>w��@)���X'�h��i#I��I@#i�Q�0ik�Љm��v�Z��:Q���FCQ	ъ�#�OQy���%��,y�v�]�~��h&m��d�;��������{|�\!����}<��_]��Ns����'�U���O��������}g}|�X|$X$�o��]m���}��sz.
�J0����q9x�X{?�}��W�5�'���R�R���`�8h�:�KV���o���.F���א6���Eb�Wb^�#�Wy>���ۋ��P ))	��z��
t>Hr��M�eh%nެ�ƍ���L4߬�.�������[�����H�������Z�:�5�b��b�v�\ܺu�7o���;8f̘���>�U�C�sv���,�Ṣ�!7f�����`u�ӧO����@��F5���3����m�6������W����Ʉ��Wp��C�������\�wv��Qz���HKKæM�0}�t������uuu05v
���������������7.\���a�����a5hP!���/��P �7��J�S�w���6����زe�����ݍ��t�.nS fR�[�0�ł��h���A��chh��լ�P
uGo��%�\�ϑSٚ�p��(���%(--Fkk�ށ�ttt���%E�1n�2�R����"U�$�B�d
�]�������ت�l��	(}C�uD�<I
��i
�2V#?/�BJ�����8��ms���w�'�ֶy���PW-�_�������5U� K�����yw�ox� �U`�4����P�Ϊg0fr���7"k�<B�a������;��������0̹���jAFL
��ۆ�Nr�dN�J�!����h ��b�т2��/�4�^��
��x�XJ�,�#Tt�`�+�_n�D��8�(q����$��D�'��	M�a܇$��'��*��u.�z�]�����25���*���O q�H'.9D)�#	�I�+N/�"h͘G,$�n^�¤�Hݾ��8�#�Q,\=-�^�s�M���8v�piJ�	�Ft;Sau�Ø]S�.�� ��7��(W���Ǽ��}p�Mݗ��L
�"�򑂫!�(���-���n/:�PM"��T)�*Ҡ�e� ;|&�"_���?�G4��$��`0�]���6�(�������ޘ;�lvE^R�U��8��{��7�����E��\�ي�)�h��	��t�����I��������z\9u�W�G��f-��d2�N���=w��04�]�49��nW!�~*�=��j�����%�t���R��|�?��ާ=0���U��YU�(��&����H��C�@����]���QW3!D�H;W+���tJ�{�s��=9�A8���˧!��i�������Ky��P@v��Mh6��܉B�K���o#�@�SP�}
���f�XtƼO��H@���{������Ӑ䊌u�8��)��8����
�?������_�ˊ��{enr���;�@�RO��{��80�W���-Z���*�7�x4[!��c�:_%5�Z��un�%}D�>����&�#������j��Й���t!�")`��8�C7T,Rо����g�*�ޕ���i�@�L��@�"P����2E�}d�?	j��<�=�E�_h3�=�Q����y k��(P�� ��;��!<�p�o	Ը	u�n��1\�H7��.�<�Qx<�m�O��2M;�8���8E�Z�>�A����NUk��Z�Hڲ�ci�#�l�U��22��C���_�X�Ś��ۦ���U;N!�'�*h����GA��b������[-
	����Bo�gV�n�����QH��>��^��N��;��Q)�(Wɚ�� #��"ӿ3�~�ŭ�������/�����ᤅ��G:�=&�(�(C�S����5�]��8���}��O�1\��   %tEXtdate:create 2010-02-10T02:38:05-06:00���   %tEXtdate:modify 2004-08-29T12:30:04-05:00�i;    IEND�B`�PK
    x�HO�0      _020_/resource/18.png              ���PNG

   IHDR           szz�   	pHYs   H   H F�k>   	vpAg         ����   bKGD � � �����  >IDATX��ylU���b "TDFY"��H�R [HM\�C(*�)Z@�He+-e)eo��Rh��k_��-��ǣ}��ݙ[/E)�	��2��f�|�;瞹O������jm�z���2�t��A^#�ɧ$�_}�Ӣ�����*c���[��UY<��㮨�b���d>3�|��1�v|D���	��(��U@�Y�B�I�@�e�~],M�K4!�y�w[��$�Ǿ#��y_`�\�y����W���6z���Th@����AA~@DD$�i���| ���N->q�BK��!SG dz B�CN�t�Χ8s#8��{Bڑ�r?J�D�6Ά�ܑ}ē-	>��+����m��L�^��+��'���n@_3���g�(2��$���]a������.�܊���bg8sE��=s�Bμ$��? u��#�,2��IƓg(�#J�	鄕!��� ��`�R�$��~I�/u�z���5g[�<A�Lr��R���z���"s�<��2�	��y?	pm�i��F��V.���U
`������Xj�`]�Vr	�ȦS�E�1n��=�'F����A���dy�.�Sd>�?߬ Zt�� �,h� �vY� ��u�L���אkD�ט�������Z��K�+S8>GՃ) n��hcen���gp��H��8L���_ᘕ�PX���R���� ��L�g�yl �GpL��1�
�F���l�E���7X��XQ�T߬�f�ycY,�'g4x�\1;(Pu�i!�D�k�� C�2����xd|eaJ:Sds��W��T2m�'��|�?��� k@ւCb<9̇Okpn3��>�T\�Mp������f���%�q���t:X��G�5�i�9�.�co �}�S@�r�}sͥ�>t��$� )����b^�1a���9�t��M�̻�d� �`�J��Ԍ�]o���+ �kMU�i]LS!K�f��$���ِrRC<�A3s��6�mo�썌����o�ΥcGe������y�;I,�orW��(t�芲-���Vg)��"\���;yR<'g(��_�T���D+����d��DH'��ĥ�Pgym'E�<K�pn7�b�X���ip���ʅ=$�W���Dȗ�(7���u.T�����(W�Z�.8SV���f\���R!���\ �I�������Ը�=�$q����*����6LC�se3.lQ���W��N�"�TJRUm���iJ\�z��;��ΰ?Mn�������� �+��7��	J�L�y9KU�IJ�t�7��ߓڝF�����~�X���𬿉��.���T]V�T�&Q�����p��b�~i�~ٿm	ZQD����5׋M�5�C��Ҳ_��Rĥ��ͬr�)����-�ثCi�բe�n\�+�HG��!Zv�&�l��۫?sZ�/��צ`�4�/(7��|�l5�:;�U�ɭ\�#���o�{�O��.td.��	|�[j6�y����r����C�񇷵��ò/"���Σao�2�ׁ������ql���.T�=�8�   %tEXtdate:create 2010-02-10T02:38:05-06:00���   %tEXtdate:modify 2004-08-29T12:30:00-05:00I&<(    IEND�B`�PK
    x�H�%��  �    _020_/resource/19.png  �      �      ���PNG

   IHDR           szz�   	pHYs   H   H F�k>   	vpAg         ����   bKGD � � �����  "IDATX��kl[���9�kǎ�$��4�
iR��Jɪ�U\�R`cA��ا����� PW�7`�R.�V�
�P.miQ@"	b�HY�5�����8N��9/|��:�&n�{�G����������/�5�woY�vMs��|4���T"ͱ��?ʾ���7��X6�����k�����p��������\R��b��|��'_�bϷ"��b�r6�.��Z�����$�x�s���%����EW j���'�S:}�{��׎��Z{��߷�ލ�_,���s�yB~|�Z�v��rXȇ�"��;Rj��F���JJ9GjI�|�&�n ����=�m����_�����C�~�<�y�qFG� $�(�y+�T 	dL�l�6O㰳�1�l�����X�?C�����V���:C�˘p6��
C���,�<���HPs^�xJ�go9[�H6mZ@E�P�,矟FQ��§9���v�~�.��@S���?r���ʪZ�iC�ꠢ�>ph�!�����,�^�����|2�����ĉ�/I�ț��&�j%��쨩�@-`�1�PGJ�i��m<<;��L`?PTfy`�!Ia�%��*�����X��� ����Ϋ`Y�o�E�� =z�h�2a~)0����܀(��}`�b��S�n9+�Nh��7�v32�̩�*>���":��G�}�Pu���)����Z�N.��J��<WRcp�s=��z�@��}1��E�0bǁT�k2��`���=�]�e�ZύNg���#1xj��l��,�mO+Nr��^�Ћ@r͟�dqG�� `h��!�̃�>V�+ �,q�,�Qʫ:��U��pQ����~��u�g	�A i�c��z�3@d|R:��@���� �����4+,�m)���7��g@�%�AR�F}::V�2#�6�:8��&�<qp� 8�9�<Kk�Y��i&�p��i�$���E`ls@���
-�v�����}���i�q'uA�����yr�B��T]��D�>"�F�4�EA�|[���" ����B��$J��󙷼@@Ni׋HdJ�H󹕘(A@��b&
@�}��/���5�)K��8���2��± �����0�p�wM�q�����h����H����1� K�0��Cr^���aK�l���a���R4(����WL#�-x@"�0�)����/Ǯ�5��}\�+����05�h��j�(����ad�䟶*��YǱ�y�7�7q������HH���R��d%dAf!z�d��o�����Կ���J?���.��NY}6)�z���W]
�k[.O0;���g䁝���a�Y����cIF���-�U=��)TU�*QT��czn��r=\=v�Ou�M�!�%���N���m�x�8��3�A}��u�d�KE�v2?Ǚ��ۺa�Kvt5p��G�HAKDb���\w�7�����x,I���w�X�giS��]Q�ȀX"������>���˞�3�|�[�r`�7���x�WWT����#�   %tEXtdate:create 2010-02-10T02:38:05-06:00���   %tEXtdate:modify 2004-08-29T12:30:24-05:00�LF    IEND�B`�PK
    x�HSZX	  S	    _020_/resource/2.png  S	      X	      S	���PNG

   IHDR           szz�   sBIT|d�   	pHYs  �  ��o�d   tEXtCreation Time 08/02/08���   tEXtSoftware Adobe FireworksO�N  �IDATX�ŗk�U��{�s�=�9/f�����@��(�Z[�Gc��@�R1�R#�Z��Ri5�!�P��h�Q�Q[���"�8��T��'̝��s�y���^ԩ�Jq''��d����k��_[c�*�}6�_�R\<�ɗ'j�/��� zn�?�������k��Ƙ����O6�!__2g~�s��W׎����-m�F���U�ۗ/f{�Ny���]O��}��0[瑇�,4��;��OH'�
t: �����4��Nz~�L���s�����[��']���qS&X�*P�U��Qe TL B� �]��c_���o����ɳ�y�������1MILDd��2@XZ�*�rK߬ة�
�����ڮ���}��/�����Snj~��qj�DM�96D����r��s�i��&�h �\�({���~���:�~!�]B���Ӣ�j/�x42�C���ɞt1�!�JP?~���P�-m}���!�����}�]���L���F"��=���=Ͻ�4k���s��'�5c&���h����u36c6�t��#xϫ�W =r�ݐ����Kz���P�4!%�c�yc+����&H�Uɱ��(0�_$��s�!��&�.�$��ZZ��-����Ҳ�6<�;]K�K8~��0�N%��V����sb���K&��b���l�^���Sx�G@J*�+���S1�3&^q�ͩ��J��]�1�7i*6<ƯV�`ŊL�8���m4L���' bӾ��g����8�W�f��;���f�������_	*O4�vD՝�BȊ�C��(�.N�(|��?�ҥKY�h��ݬ]�5u�H��PNCF�f۶mlڴ�x�3f�f�V�^M]uS;], OG���z1j ��y�,'�n<s��A��c��ͬ\��Q�J�F���Î����o�I�P��m,�`ǎ���s0��ضC�K� 0�i�U�c�Q>��t��w�|�cժUTTT�.�����G7�=م��@��ٳعs'���cӦM ̙3�����R��|m@�3�&K��AD@;��i:?�3#'^�[--�r.�t�l��hx�v��L*��p+S�L��g���d2/^���H�w`�D��²6 ��D� (���N��������M��q�D�"�����5��^�3]���a��P�X���:���6��1a� ���Q���*�D�q*#�����K��!k��}���r�c�G"�E��N��E���*�\t�� �� �B__���K�X�*9/�t�(��|R�tI�t (*��1�������A�a���}��}�����$<�n狡��a��� �`r@�dM��}��@��v2�=ئD�@���о�¢O��
�O�'��H�L�(��bO���%1F��V|���
�	&@�DJ���<��P���=��ov���S>	`�ч~;����U�dT�%�G����i1�؏�!�G֒!$R
��)�e+�@�(}[� �{�[(���<r���%/��!�7�h`�_����Y^1TF�B2���o!���Hu
tY�Ϥ�Ǧ�~FҍA���6��WQX�bɹ�/���`� 1 '��>������)#�Z�8�q(�t����}�n�����cB0���Z�	�܌��2a%,����Q�w����e �N� B��}O���6�~X���+3T�@�sH5-@���>��1 c(A�{�ޭ��CX�a<�|���ޭV*-$)�"F�W"���qѝ��z����1�"�pȝ*ғ��h�+�F(��xg� l����E�m�S/��$���Ow��r��U��ƍ�w��r ��	cLp �࡫���.oXW�P'V��P~��7��f�a" -�	��^��~R����݄�@��|���p������s	x@�1�0�%BX@=�;��_S��~x�+3�*l�F�veDI�m�X�G��B�{���#�����]�����4��ٔ�w���a�3�'�66�ߜ���C�ZD$�6�1�4&(�'	{�p;r�h��5�x�?�.�@
�}��K�D���mc�x�e�u���\���IVWX���F+��W��S���j���޾}o��{����Z4_p�gs9}�Rq��s�,�b������̾�v���/��d��w����|��R[MX�+e9    IEND�B`�PK
    x�H:��  �    _020_/resource/20.png  �      �      �W��PNG

   IHDR           szz�   	pHYs   H   H F�k>   	vpAg         ����   bKGD � � �����  �IDATX��W{l�U�S1bf��`D#��H�K�c"BL�Bѐ@$�!� 8�5��F�e/�`���ֵ{t�֎��nm�����"���&'��w��9���{�W!����ψ�o^j���f������ߙ��������xĿAj��E1���u��\%P�(P�$�9,��'P���m� ǽ	�D�������ı��ĵ��^r#��(�^ ^��h���v+��8����=a��w�s���8���:r� 蘋�o��InZ�.��&�#F ��ڽ*#b�_%�:G��mx��477+���pW�A��>�{h�������e�ޫhhh��\�|�є�"����{%BrKźh�;�hkkî]�����@ ���F8����QL�y8<������V$''#77W	q:W��r��E��Sv�o��ޮ�o�b���_c������AGG�_��ΆG���C�,F�EOOf̘��'&&�b������{me�A�����n3Ys�wT$������jA�����eee�8c��Iջ�nE� "::Z͍��B||<3��ñ��"�M��k9����#9X��@G屢/$���	��鈉���I�PZZ��
�|�0BU�ھ$$$ 22�'O&�6�v�"
��.�I��^w��i���oB�5�f�j�*B�߯ kl�ۑ}�:܆�R�hn��+K��ݭ��Ly<U6��]cw�M��������[0���~�`B��Z����H�VUU����YY���������#z��{PRR�˥�e�yyy���4�U0��B�2��}�<B'R�w���&ӆ���	r3v��T\�X���/��sn�-��Gڪ�"?e�23�����,����x���j����x�U^��'������\���T�$�ahMpS����u|�#�LF��i�e<�G��z���n
1Έ>��F��U���Sx�l�]Տ\b�	�8�h�O�3L_1��9VMxL�A��{
���t�G�c,Z.�F��A�45D��	�@Ц��θz�_3@�>�0�+q��@eD���B#ѢEH�� #��pb����&�b�ZrT�'��
Hvп'��D.QL���"���Z��d����,�M.EW��j�Z��������H"�Gu����(�C/�ў��3Ҫ��W����1�=�}%��k�9��X����YH!���o��~"�5:ni�&uk��3v�9J@�τ�>4��pǏw(C��B��#`!~'.��+Q��85Y��vj�
�ib�z�ɺ� ���;a�����j�)�+:e:�rMX�ŕj���y<kxؘm�;��"����%���-w!Kq��iʳD&qQ)�b�5��gY�<�5��!P�QB�I9��@^����DD���)�L�Y����Y��`������b��n��iѹ��"B�=���7��I�ߛ��\�kg�0�Ӌ�|>Ms��K4��Ko���[e_�]�gp�5�Y`A��͕EH��=$-����˰ncd�0p�5g�\�N���y���Bٜ��@�M�[�gC��%(˿�+حp1~���E]��+G��.fʽAu���ئ����8�)�L�����N���GW���W���r8-G�ΕH[���ͫV�t��˙Bs����4�3���I�[l*�Xmj`݃�;�¶�ΒmO�d/��%?0ճ�p���G����} xPMV�   %tEXtdate:create 2010-02-10T02:38:04-06:00d�   %tEXtdate:modify 2004-08-29T12:31:16-05:00	�b�    IEND�B`�PK
    x�H�m.	  )	    _020_/resource/3.png  )	      .	      )	���PNG

   IHDR           szz�   sBIT|d�   	pHYs  �  ��o�d   tEXtCreation Time 08/02/08���   tEXtSoftware Adobe FireworksO�N  �IDATX�ŗ{�\U�?�>fgvv:������.}�m��Z��"�!HDK�Ɗ6�S��Ǣ6J�&��b�Ð�RR)B�J
t-��ۥ�����̝�:��ǝ>V��p�_���9��9�����9Bk�'٬����/�K�_�pEe]��e׫�sܱ�����]�7;��������mb��^uc��s�N�6̱�զeX%��Q�#'Wt�#�����:�{�o��*|�X.D����Z_���o���U�*@���BP(����ΉA2�=������zF�� ^�5�p���n���x���)@� �,x K�`��;D��;���:o_����x��i�Ͻ���W�jK�c b`T�aF �f/]�N�ͬ�*��G!��A=��k���o�X /�V5�����%	T*�"�XKA���K�E�e�
��`$���/@���q{;y�O���_?��#�"q���v����Ĩ3���dN8h'QUI���O7I�J <r�2�7J�STT@Ì�$�̀�Ap�&�K��}_۲M�����x��߭�5o&�BɀC�_%h����-�25���w9���1�Dj�\pF����3*�a�E�P��Dn��������_hlm��Mjb�q�g�?
,�G ��k�����aē`�|�Յ9�&�/����o��כ�'4кr-�{�H�0��+�%/�m�Z�ϓOl#W
X��62v��`H@�nL/�'}��[�����)��!��,�]���[�������������C��ϑD&�z���ݻ�;���|�ys�s�Nf^����o -%���k��' !���4y���@�_r�׷�+زe�֭c͚5�i�#��&�]��J5Qal��V�^����	����	V�,ps�'�T��;�-�b`�uֲ��T+J��l�<1�ִ����> --�X;CL#
�x<NGGMMM 477G�lB�%�e���V]�ڠ��mS���f
�C�a�&`{��?߸�t:M�X�����~�f�'�H�>�6	�%��q���SWWGgg'�-��6�x��a��DK�! ���S 1���4���Aؠ�4LTz��y����E>�0!UI6;F,<�i9�Kꚪ8�<������{�&O���#�R�Xh顤-1M��0MQ+ҋ B+����a��ӔRs0cU��P� 1ÅP�
0+,�k�Ƚ�^���)��̾LM~'�a�
Ct���+������hW �rbV�j{���4@X�ӵ@��ď�sCe$��@���NIT�� �'��8�R.�%}�R�"aF��Y�1P
���HE�dAR�S���J�����}������K��o>:�<�=���"�E�ϰ�3����+�Q���
)]�ڹ
Bק���
��'�Kn6�.�)8��@>��'���c��EyEd�Ez��Q��_���n�w��Ze�F�QN��*,�	P�~��(ȕ8�N*QVA9@��0B6_M�zH�Ez.��ȏ���}���q!�qj+>�r����h-CCe��M�/${��?
:��B��%��:��!s|����0�ѥ,ҍ��E����@�l!��r��1�'�.��άL`�6�!��2\�{tf�[d���!@+��4�AU_J���$�v?D�[���C�����?R+� >�
Bk������3�M��8U�mcP��Ìo�-x��X��D�o�0���PQ��r��ܣ/ AX*�=�☫6�(W}�e��T�bk��N@��,��֖�5��q%L�X����|D�RHυ�0��XVB��M��
�оh�IX̡
�x�<�V߹a�~�/��i��S
  ?]e.�nE����5;���È�q0hL�
�A	�{(�Q�By�-��C�F������/n�����֥qG2!�	4�Ӷf�ğ5Nk�e�'�]VaƢ�Z�4�4Z��0J5U�"3G��+�=0v�W�`[ٹƀZ��C�e%��ꟺ�r]kk�-��S�Vz
"^V2�_�h(�\T�a�g�0�{�w�r����[t�#����Ǻ������1�+�_�4���du}���M�)�ZI�W�Aa�q�C=�ûw�w���E^-���q�gs9}�
q��s�2Y�bôꔒ�W����җ��u�~7�7�O��Be�ES��a    IEND�B`�PK
    x�Hl�4��  �    _020_/resource/4.png  �      �      �3��PNG

   IHDR           szz�   sBIT|d�   	pHYs  �  ��o�d   tEXtCreation Time 08/02/08���   tEXtSoftware Adobe FireworksO�N  (IDATX�ŗy�]U�?�n�yo潙�t��v�B[JgԖ�"(
B�D������1��Z�c!Ť)�RJ���vZ�v��������9�q�L;�A�n�˽y�������������Ӽ����߮/\����M��ݬB���o��������Z�g ��O������ʛsۮN5��k��r�eX%��QAU�B�͏)��yt�k��o�7�k�N!������.�R?kA��� ��
@��}�.� 헩�1���t�yσ��G�#�]��W�w�O6-�Xa�A
f�-c dt � L0p�)��W��w��Տ�=uV �n]����BnI{�p�H�aFF��.�j��YV&���!�v���}�ݿ��#?�D /ݞY��d�^�B9џ�)0�`ا �F_Y�^63`7�V�*��Gp����}�#C��`L>�/Djզ��m[�"'J<92��l|�D`f*R�J@��'�N#�&�-�Xؾ豗osVl���%?��d�b�hg:����AK�&�R��x�|� R'H76�;g)�u`&A���l4�}a��gT��M�ܖ�+�5�i��TA	�ՁY)`�㚰�Iҿ�U��\�X|=���݇?|�E��&ۚ��~0�� +7��%��b��B�퀓�$�`F�}"��[�����Ѱ`%�`���4��J�c��a�%��8u-�����Ι{�p@Ea�����.��{�Ǝ�倊�N���0�EX~�Mط��_���_�
���$�l�m��@�E�!U�|~Ǎb�� ��ζ/~�n;�M�	V��g�P7Ց~j#�}{�����ӱA�xcGpi�q�2�l��w�A[[۶m#����6P�N�TH�Cy�P��f�?�rJkn�����Y��#�CǱ�ձ��΀�)|�:����}��X	CG5���OWW�|� �J;�� DK��C@2e�����L�ih���aXe(+0�`$�.^A�e6a�V�'���D��Ç���#C֬Y÷���r���m�e����4�?�4E� H/p�6C�s'#�-�0-���<��\��ïp�ƍ�=Ή�h�	�m�Q��
T��-%h�� \KO�]%6N�\y�aGk�<*HfS��2z�Dnօ���O�Ћ9���*��� ��wo@�P�~u��H�S-�d��Nd@�#��)A�����n�V4�D8s(�G�>��	����OkÓ�=VK%�{��e�
�e�%'�x�s9��JbQ�V#�Ff&=��M%WA@��Ԫ������O�e7�?��8�2��8IX:sL��r� I/Z!���*Ț��<��|����z��i Zk��}NUKS
��Ba4@��8QP�8=&��SU�BX%_���u����<JE��{^�C!DRaLY���}]��� ��2�����b�r�c}�R/�F�㨂�E~/*�'��>&NN|#9]�#�(�_q�8��@����=����g:�g֥0L�պ�	�����,�yl3�4��A+��4�iD�֓Zt9����<F�[��n��A������|`(�5B.��}���׆�a�T`�:8���"�R��؏r'@��H5a7�#�IcU��S��]�@��hϣRt��������Z��uq� ��e��[=�8;�T��pR�@�u��#��Bv$Z"oP>ԆQ����B8�F4߁$�P��R��=����ԏ�q/�@��:�R h��F��+fw5�nJ�hD�i��DF���3��D��о�R*�WE�Te���I�߯��k��?���j�k���Bh��~�53պ`�3;�XI���vmD�F+��!:�ZM��ȉ��U�,>�y2N��"0��θ)���f4?so�}K���R?s^���C$��JOY�ր���E��'��}���;~��{�w�+����':�����X�����s�θ,�k^j���f��Ĵ�V�UdP�V��}#�#{����塗x51��?��%��p��Kť�۸,���0�JɪW����M��bU����l���>���nD`�A�    IEND�B`�PK
    x�H��]3�  �    _020_/resource/5.png  �      �      ���PNG

   IHDR           szz�   sBIT|d�   	pHYs  �  ��o�d   tEXtCreation Time 08/02/08���   tEXtSoftware Adobe FireworksO�N  OIDATX�ŗy�U���.��7o�3Î��e�j�5�4�[���RjJ��&M�?j�MIjZL�R�h�Zc�-b�Zi��VFQ������ü7ｻ�s��}��V�ē|977���w��mGh��$�u&��%q���^Z�P�iٍ*\,�o����Wm�vj��3������O����ڙs/��7-�3U��eX%�
Q�+#�P����{�=t���W�*~��X%�����ml\r��sSfTN5 @IP1�T:탎�a	wd��#������ۮxZ�� ^�!�t�57<R?�B3[R�0 4hY@z�#`��?Hί�ݯv޴tc��g��-3.Zx���מE�@��H�aF Nv/}�n�ά�:�O@܋�~ݯ�u����� ^��z����uִ�ȠRPՐ(ǂT�dP9� Q.�`��΂�ӂ�������?w޸x��֏�U��m��[M�:F5���3:⢅C�����j��hbz�(�`���ΑNCӬ�d�͂�Apߢx�K������[�}�2�{�~�0o�����w�B�t!�/\EUn�݇8�ڟ�5�#7k!��`B�OqB�e�y�S�4��P/G�=G��_ink��Mnr�q�gg>�� ���Ufk��E7N,����0���+��k����6�IM��^��~��(d�z�/�eϡ}�z�~��=B��X��FF�vJ��������fy�m5W}(��՟�����FJd~ߙ�YKV�c�~z��lڴ�ŋ���M��/R��c��v�5tt�����{�a���ڵ�9�]J!���-%��M3�n�' !�Q3�u�H�@@�8��	l߾�6�v�Z���غ�j&�]���M!ml�r/k֬a�ƍDQ�w�A��~��D��L.���׈�|`���JgR�%A�X��r��Zk֭[G� ̞�|k;)�Q�4v�M�61e� ZZZ�u� �A��
�2D�Y�'���>�r�1s�� ;7	;�T��-���P.�Y�n���u�G��!�6ۧ0Z��;嵐����N�-[��6o��	�a��DK�!����&X 3���4��
Aؠ�&+?��EW����b�eR��|~�T|�r!�4L����s�.�����Kϱ�i�6	�G��.x��2@I	Zb�L� `��^	d� �.�����f��x���j
�G�����C�@E�i���A
�<DP����F�Ç1�/SW�t���h)A�� �'�4�H������pbL��8Ut�aA�s]�;jTb�Q���)��#T��x|& x�B���t�L�W
�RR��Ӌ�J
�xAR�S�������A�CT�q�L��o<��"�?��e�2�%�����iϥD���rR'd�BJ�R������hB�`�~\����Pn����4% N9>�N}+]P>2�~��A�
B/�{Ȏ	 Zk��~Z��X`b�#d�t+���Cz��	|TP_[�,�!!�q2��{[q�D�C)��GE��DaT�x�bYN֫2(�H�#���*�>�m�T�"����x-Q~z�' �;B����+[�)�2�-�mb/�З�/��=��^�����k��w@3P�H�
��w=�%}��y��c�°m�e��S��t�����d��)�@II��De�"[��0%�_@z!�碃��X��P?LB�+��6�}��{~�;�݃��]�R���=E:S�乳��:�t��1�o,F�*rͭ�Ϙ���"%SH�FG����qH�讗��*��ɎH���+�UW_ڲ���>C�agVa9`9Va&��V
���GF>*�P���˨� ��q��?��v�h��> ���ބ�LaV�'���]3��3Z�5S���A��$]�$cj��J�e���PS^9z�B߱r���ۿ��T�k`�ZGڔV,Q������U�ښ��M��X5�N#XY0�%ё��F�G�q�p��o�}��|��/�u��"!� y��,��%�W��6\��ml���5f:gb�B+�
�2*�p��`�P������'o�W*;��G\�ę\N�X\<g.�d�Yn�V�R�<�v/}�)�u�������a�	� S�/ƽ�Q    IEND�B`�PK
    x�H�4��)	  $	    _020_/resource/6.png  $	      )	      $	���PNG

   IHDR           szz�   sBIT|d�   	pHYs  �  ��o�d   tEXtCreation Time 08/02/08���   tEXtSoftware Adobe FireworksO�N  �IDATX�ŗy�U�����޼���73�TQ@�
Q�B��-T,�M��bmp!Z�6�&�5��mmS-��VԢ۸�Eh�Ұ��03o��̛�/����D���x�/��������|�RJ>Ϧ��䷮3�.�rE���BU�ԅ�c���={�����{[Ji�)��OX5U��Ⓓ��M�W�5�&F�xZ�M
���xf����G�ڼ��Y�����f��ss��M�����1q%���>��.H��C��}]��{}�6������51e��WjΞv����@�PK H�A����P �n
�w�>��-S���:#�-w���y���?5�����R�(e �d}`C`���8h������v�>�����9��S���JL���%o'&M��Ad��	���=��	PS�)z=&i擻l�OZֵ�=�&��뿳�n�4vϾ��R[7�q�Ɠ9��SpJ�&�%o�IH������`��N4?Ä�4x����:������~����g���M=�B�4 t?n4�nX���//� �Œ$��`��ng�?�0�l�õ�\ڒ�����7�z��S^&F>���C�q_��j����(]]]8��a�;z���n.�:<p?x9p�%�Ϫ������$*�QS]Ex���mۘ���#}L�n�����/x�\��3�л7�G�Ff(�RJL�$��`�&A���y��'��8�/��y�L��x��[8w�lۤ��l�"�uY�;$��w��(��z��(׾7�Ce�%��@�uR��b��G����qg�g�l�m��0��9x���|�r\ǣ���u�̵,˲pl��[�7[E�'�C'<P����-�.�oa��i�aP(p�u	� ���>����c$�I񀎎cd2�����5aZ��>'vp@�ī��M���Aj۶�}���ys/bxc�<�ۍ�*,�"�ˑ��9��Z��hi��2謙�a�sW���h�B*�"K�vj�붅R�]R�[��ȕ?��dLOJ]�?q�#ߨ�����������f�e�ĒE�p]�TTDy���,r	���Nho㛭�ycŭT%����^�M�s��*��n����m_I/H��5]y�$Q���{_�gpB��:Z���_����̈́l/x&�vI
L<o8��M�*���[�;{"+W&4ϭc����C���U;��F��7>5a֌;�U�*�5�}!;��7%��k��2�H}-�Xn9��4��lP\��P�s`'m�}h8LhPi����"=�
OO|�Z:x�wv��yF�5�J���#M0}F#Dc(%k{�r���J	Iz �ςl�3�c���`X��"=���;.������n웟�(^W9@ �۲N�"����r:�R"O��C��@�8J?��8.���Z�ܺ7�6�d )ex��/�M����DP��Q2�<�.&��Q!�`�*
B((�@�((�^�P�6�I����86��P�w����/"�R�Pس�me���U�R"8>��i�{6P��HM�r\��Nt���q/%BS�z��r!@%�K�]�fۿ��@� �Bg0�}l�O�MkZ��:J,���M���B�����R"�z�(*���6�D,��ŷ-�M:3����(�@� �L��_}����F��������wt�?���n��r	J�� v>L<�ߏ�[E��`�;�k��{��\�DʙX��%
���b.����5Ս�*�x�b֦7~=�e!��BN�����(���m+Id�#|��p��X䃽��7�"���iRJ�8 �0��^�ξ��ƕՍ5:�h�$�k�wF0P5��ld�
!}T/G��C�+Q���Ahtc����#�k_�����2RJkHE$�P������|M���4�W+G@�M�</��+)Q|4i�J�@��Gh�	r�(t1�����Wy��\�@���;eU\�DPk�����K[ZnJՏ�iU��0D$�)a"=����ϵav��h�ۿ^�<��N�I� 
RJ�S�D�D�[&p�sb�G����H׵D5UjEJE���xY��w��dz6o�a�q��������8���K����63'�d��j�a��%wg:ٸp�R���o�Ϻ)|��ߒ��6���    IEND�B`�PK
    x�H�5��g	  b	    _020_/resource/7.png  b	      g	      b	���PNG

   IHDR           szz�   sBIT|d�   	pHYs  �  ��o�d   tEXtCreation Time 08/02/08���   tEXtSoftware Adobe FireworksO�N  �IDATX�ŗy�T��?�z�]��Z`��GD�C���I�(BY	�bE�DŤ*�)C��R5��#�J(Q0�d���..�����o�ٝ?f��e��(���z��~��v���-��|�%p2�_��8gش�sbU���@�Zy�i�S;���n���}]km�,��w
<;Y��Ƌ�*6�h�S��X��Z9(��]�/g��?�n�p`�{��������!D���]=���%�ƌH�|P(��m�v�N������_hyq�헾��G o.�O��`�3�c����
�Y @��� 6�y�.�`�`u�wpw����&����Il�u�yc�_�����qtD�0�(x����fᛌA Q�sz�;L����}�1�>��+l\�?���7�5�EA�AF���<p|�&��Bg��`)hUP����C��{�y���;�|)�mBDo����L<g�U�(��"�M�@��\�� ��J��D߄�V������/o�<}���_n�%�g���q��ֿ�6�B� �`���y>�M����}\P��_?ɞ��%��@k�V�f6r��	Jj+����p����.��ƌ��H���Jq�҇�e��8�Q��e�1�ʚa���;ؽ{/�ky{s�~�4��.`�i�|	�O���Sf�7��>�k�@�j˦��^v�*0y��J��	K|7��1��yǏ��gݺuttt�h�"ƍǦM�0MH��f�1�\�X~��}��ի�D",Y�������XE�ᣫn^��sP��ܹ�nm�@]�y�����w=��lٲ���׳c�R��e'�0�ݺ����rYV�ZŐ!CX�r%���<��C���ƭ�)|3����2�0.zV������vӝ�����с
�[�n����H$B{{;�\�H$̪�>BiY)=�ݜq�t<ϣ�����:b�۷o'
��:,����P%Ċ��� G�%�_<���˦A��c�2\v�zC�x�b,X�m�,]����z�㩇��3g���kY��.***�?>+V� r��"aV�x��S��Ҹ}i�v��o
���h��́b[&�=)̼ży�hkk'��0j�H �{�Xf
��2�$S} �u�]\u�5�B!����.��Y�%��Xy���C�H)*����1�XBy���3���AJ�4$��N�I�v0�i d��2i8��$�f�$	
��Z�{�:Qc+�%�(�C�h��N��m���$�ly~	�ړ�J�rZG�$ �]�VJ럗s��T���sh�!dT�8d0*o�9.��P���<�@����w�i2�`�2�`t� ��
F#x.�f��L���;�DZ�c��,��y�8(��s\<�;������F��YJ���5h�.*f@D��ŢUѐ܂��?)�/��x��_�\�rțn���q���-+�ڋ2��&xY��
���e����=�'��&(e����m��ʱq�~�����Z�w����q�����E� �@nx���L0W��rx�nR����o[(�&�v>���	!"B���Զ6���-�*I�l Grg�jo���,��l����@Dt?�F�#MW��H:�·
������k��� �B�v�zϠU���EƢ2�C�^I��X7 3�E����������)<_�P�*�F��B��O�>���,,�#G�ݓ~�� 	d��!g@�s�6��v�6� 9��
�oƑؙ>��a���"d#ZI�t0�D���X��w^>��mriK���_��M� %��Z�?0����9�օ�+��#JH�P��`�b��l(��ݡ�w�zw�~�k[a�]/ׇ���d�k�����G�����k���
  ~s���9uk+�*��+�8"AF��E#��C�y�c��Fy
e�(+��u���e���y��}��`G���~G2!�jo�T&/�[�@�кFY6��� >ˊ� m��h�Ѿ��
[M�S���iϽ�'����x�\i�Gk�~ᡴ�D9 +����b�45�^WR38(��TC ^LN��]���K�av��Б��`��ć�W|��Z�_�^ 
$��a4㮜���������`��L�K$2(��Qv�w�����j;v����;�?,�Ȗ�,�%�/q2�ӧg�Y#F2;�`�!UJ���׻��+��u�~7������A���l�    IEND�B`�PK
    x�H�?	  �    _020_/resource/8.png  �      	      � ��PNG

   IHDR           szz�   sBIT|d�   	pHYs  �  ��o�d   tEXtCreation Time 08/02/08���   tEXtSoftware Adobe FireworksO�N  [IDATX�ŗyl\�����ݷk���U�8��8qlR�)��"�"P[H�*"D�U+�O[�VH��TMqHhچr5\�R�6@1�#"���}���]3�?vMbJ)�!F�4�O����������ֱ���W���\p^�*u�iE�U�9nzb��޽�.�<��v�@�;ܿP4|�����u�TMK$��0-�(���
8�9wb��L߇�ھ��������aw�s���'�rs�3�]
PT* ��A�����d�����~�E��C���J�t媭�y��%� � �-� �<� ��`�1��;���7,����cx�֙gͿ��'+�,,AGAD���aF ,�^� ��3+V�`�>�]t��yۼ�߿�3�p]iۢk�;˛�QQHT�cA4	A�+��+(Wy���Q2�a�@Ąt7�q{;9�������� �	����z��g��(�f�wu��&^����T��3�/��az_{��lb)L�'U��n~�>��2����v/\����/����|�GUsZg�-�ؿ����4.]N"Y�P�>�{�9���'y�|pGQ�þ�A5]L��5 �p`�_ɿ�����AGI�VsO��	X�q ���̆�y�7v	X&�]]��N۲K���&[~��HY�������8$*����ܫ���<���Y��Gy�y��@�\����My]���;�/�D���\[ZSAJ���=�OZ̖-[��]w�n�:�Z[���~�9d���M������L~�!�ݴ���~.��
~�~=M�'�����$��R3���B�3V�h�y��	_�}���ڵkY�z5���l��AyU-D����*`���Y�t)�^z) �tt �hy#���&�d����M���SWX��d3J��"r�h�ioo��} ��
�F�(�r1E @KK��r�T
�%K�7� 4(PRaY�h8��,�e4,l�в�$҇�#�,#����y�r�z�����r����o^�����Ii<`�������\���R)V�Zź�~F:�p_a��DK�!��GN�f�xY�B���eSS���M�����Lơ,�`b"M4<�i9��TΨd��Y���lذU<TiG!>� ���()AKL��i �)R�@ �@�`�I�n҇!�l���29p�DB*@hEm�Gn��O�E�*�8v�eb��*�a����M��?���Ѯ@��=V��� ���` ,őZ�}P!%v��9p��B���� �0���i ���.�;g���YP^,8�b��R��.F�P��
�rϦ��5(-}� }���~@�=����[�O�N&�.�+H��0a�(I�;[��we�����Ѭ|�{(�G��w�i��q��Ewbb�)8Ņ�R2�(�Ss�ȷ��G���a�-Z����z�^�k��ZM�<����,0����<�
����$��I}��<�L��Ƨ9 ����G��ݿwo��7d������(�����'34����&A>��<��ˮ��̀�!D���}�냉4���BP4�.*Q�b&�N0,�>�Oϛ�T��h�%̻h/�Ș���Gx�@�B\��S��\��qN]chX��4q�<0�$��v�Кi�e���`lp���nʞ4��Fv���C����إ�S- R�E��ZS�G��KXr몦m���&f4��q��xaXX��a"��ϻ8#Ā �R/ua�I������=c/�U߻j��P]�e��ZS  5 ?��\~�y��+�Sqb��H	f�M7���<B?@k��1�@�|���~:�����A�Z���ǻ�c?Y���E��Z����La�~��,\���u3���3 R��a�V�H1�+4!����wZT�5ot�ɏ���8tۚ��77��40��>�)-Z�0SP��M����u�&k�����v5X%`D@�hMក��@b���C8�����m�y����&���g������z�
��U+J*��#%�r3�41#B+��r2Ȏ9^f��@���?�<���k@��ӟr��r9������'����E�iU)%/����ům�iW������=>���I��p"�    IEND�B`�PK
    x�Hbȩ$O	  J	    _020_/resource/9.png  J	      O	      J	���PNG

   IHDR           szz�   sBIT|d�   	pHYs  �  ��o�d   tEXtCreation Time 08/02/08���   tEXtSoftware Adobe FireworksO�N  �IDATX�ŗ{���?g��}��ݽ��.�P`��"�M%�b[����RK�ck#�&XH��%�T��T����ƚJ�����.� E`aa���޽�;�sN��W�U�ƓLf&3���9������l�{y��O��&_>wq���"Ӷ�T�W�b~��C����~�/Z��{�I�G?&&]x�����4��:ˎ�R�eZ)�
PAE�B�͍���N>{�o�×�[��_� D��,]��{ѪdǤ��4�H	:��A��]�e*�aƎ�������ʇ��������^s�o[fΟaƛA��A�:��Z�`���p�uw`Ǯ�zo?��=켽�ʙ˾�����(�#�U����U�������c��e����ӿwxͻx�	Ͻ�k�ϛg�"O�a6D 띆�\�U�e��`'@���!,Cq �c���9���f�>�����!�oY�z���wa&A،:H!碍�x���/%��ձ��U0<���f	E�����4L��a��|l�zm��?+>�/�p�O���ezo�(�ʛ/�����I���D���o���g��[�a�l���?����J�%����I!3̱}Oіy�Ιݠlm)���z�z!fm��?� x�xO��+E���Ğ}D�~��˗�s�N��zNsӗ��T� aq�͜ym;��|�]��J ��#�'S(3w�

�P�?��hlk�z��o�S`������R�!�d/�f�a���ٸq#�ׯg���=}����(��t�f=f\q-�v�d�w��]w�E���ٶ�1z.^H>l�� (Iĉ��n�Y!�|F�XS�ī�m�!�mS�x��[��իY�b�����H�N�H�?��h'j�l�tK�,aݺu(�X��,"�Yh7W+�q��y/�h]2n����h2>�0 |,�@y%������\��r����S�"Qa��f�g��86l������ l��<h�QRa����"��m=������/1�F�t����p�uY�j˗�\f��!b����r�h�Z:;;���cΜ9�}��T���@i���! �X�S q.6*���B`���5��3�_;��)��4&c��
8�Ӫ�'Iw6p��S�z�@ߎ����,(}�T��Kt�
�"�0�8�R4�b�U(iy��L`�T[�`�q�	��.�����L��?��y-mT�c�m'urb��%��� b>B��8 �]���L�]Px��)�T��j�iX�s���0��@���B�C�Fa�'J�Sy ��F��� �����n%�C*A�EY[�#8864�+V�mF��~g)@bR߇l �0P@�*����2	�pp\���S��
	 a@����f ��|�<��w��!��s����`��>]A倲$�p�`�8��mv�ya���l@��cy�研7�aa<�,���:H�P(��U��2���ė>o�S�˹\�	!m@�-ز�A� ~��y���܏S�A�HK��´ lPH'�T����}BGa�5���~���tkC{R�L�G�� ����Z����D��\�A{�|��PQ�j��A�H¸��.O[��W���;k�o������_7+�֧aA�!p|�t
3��%#�j�	�',�)g�XA�Yt��
��	Le��fܓ6�+Fj^9�d!��D�l\]:qrk{�BD}�d�0�L�)�XQ;�0T(	�*A�
Jo�!b� D&4��B�j��{�m#>E U�VPF]S�A�=z����PEj䁩	� O��3�Tg��-��T�B	ڻi�<�H�XH%��V�U��G�<ɓ�t.���Z�5u�l�������:ZliF�q�C�"laX��V
�H�E.ګ"�
�-�ʣx�S8R޴x�^��R+>0��.��dB��]�%_�j¦�I�S�Ɖ`7�� �H-#
��5Z)�ѡ��=��G��)���QX��A ]W�d�9�h\(�+�������9o�Wڻ#VS7�I���UM��EU��c�TF�2tr�-ϻ?��n^���2��Z��j_PO- o����,p���L/J�Zg�ɖF3�41"B+����/e��������K�p�x��l���x{�����\���X8m��I曦�VJV��>xz���;�u��7�7���mَ틁q�    IEND�B`�PK
    x�H��\f  a    _020_/resource/admin.png  a      f      a���PNG

   IHDR          }Jb   tEXtSoftware Adobe ImageReadyq�e<  IDATXíWP�U�����6tƔ�'hf8k�琥�C$5�ŠQPkK������UTRWYD�l�m'PX�Z`_��K����������?Ɲ9��=��s����BW������ɚG^[���/�f5�y��kfp��� �(����m_�g� L���Ŵ9pZ4�t��/Q�s
���oN�p��p�����E�k�+��y#�Yiii��X,�����fCUU�F��e֏�W���"�O�\�B�W1���<�i:	��|����#S����;ͧ�;��o�wVx~�P���r�XL�Tv�`[�N�0}1�WV�B�2�o�
��t�֞"���q@mm-���x,�z=
�����l�� {�@lD��P�)c��H�˒��5N�8j� %b$$`��qYs�n���p.���/�7w$�X���`#�kh�A�s����y����5H�ᗗ@x�����ꆵ[�
�ν<���2b�j�<Z1�+
3c��V��sV�+�i�^��g�b*�ʏ�n��v;�Xϳ��RБ2I�4�ε��RUQQ�+//��Y�.t�$eee�Bo�������a����i�� 0#�<9)lx1��B*
v�B��[��8eb��D2�bx�e�OpYrA�%$a�m���m�w�u��TȎ�2+�6�ꀧ2���QsHz��}�@��b:�V?�%�@�'3%]���Ѣ�dr��Ϙ���Ȉ��B��@��k>�~�9�n��p�c1Q-$N|�Bĭ�=��Y������"pF��H#t��C�h��Um����ր��H�ʙWb���$�k8���mu�!�O���lQ<�	yC'O�:̀�2��䤷�H���I岜���o����R&('���A�Fߺ����%a���Í$B_�� ٦q��;4슍!�H����T+�~J��K`�o�4�8'e���ჱ{�.t���@�3	��9!>���Y�k�;T8����,!<g���e9�~p:��o�n�q�k��e�&:�8�DfYƝc�JNM�'����	q��yl�Kp7�ʘ�*w��&�ׁ��ȁ��s��FN��?�[1�0oh��?uԪ�@��+ZY�,N��	�v-}�-��w*�Q��8j2xX+tX*��K� �#��?�G�P�8*��gT�����g`�,�?����t5o�CG�m��4����l�>��^Au�~#	���H����qkP^]���W��{ҋ\7|�S�^�g"�n�KB�!:�Ȍ��:k�{�y�v<_X�R�(h���,@���vခB86�9Ѡba���� ٴ�ߑD����=���I��9_����Sn0�%/��ȗo�"9��-M��}J���P��!n\>������C��J�}�-��:��e�#e�7��(^�>F�:%"S���T^���b�}��H�4	����'!���w��d,�=K�޿b6�D�Fzg����G�r���V�Ϛ�0Քr]�V�ٺ�:����n�!GU��93��E;I`��!݆�_e_��3R��    IEND�B`�PK
    x�H��4��  �    _020_/resource/logo_16.png  �      �      ���PNG

   IHDR         ��a  �IDAT8���Kh]e����Ϲ���D�4�U�"6A�]���Eq�ŭQ����Jw�KATR� ��|��T�hJc�)VB��[���}�s�\��nt����̓��)�o��}2�o?�Fʲ�fk��k��f�����b�Бg��hY����� A���6Jzf���?�xj��ƕۀ��{�C��=�U���t��!*2�&'��b�hw�!��?�,/��66��y�N{ki�F'�$�YF0%X��&�u���١���}������ȑ�}��l������5���DO�u���)c�DE~,�E�jwP��UCupApw$&�F5�I�WVL��aY�g!C�0T�����p�kC���JPͫ�lUP�Հ�a�a��������"�� ��ڹ��;�7�
��ɦ�e�Ŋ��� �fFO���������Rnf�T��1���bM�1&"	�������S���/���$�'���?Vp||� ��=U�t�z��s������oW�?9c�#���_J>��э���_^����v�]������������I����k�R}?+�e���y��Q���!��ˊ�`@��BΜ>}o��;�b��<N�� R�̢����z�Z]��f�����߽������lNL0(�h�H�6P��n�߿�n���q+��q�    IEND�B`�PK
    x�H�p�'  "    _020_/resource/logo_24.png  "      '      "���PNG

   IHDR         �w=�  �IDAT��_��u��������?�_�̍rL�jJ�Qt)�\e"H�]��.����.ꪐ��xa�ltUb.1�t��̩m'�����9���o��������	#���'����o`v�^�v����<�a�k����c���/⿌-l�_�
7�~��gv\=���έ����1k������?VzO�|썿��<��k/r%q����.��ݓsc��p��Ѽua�no �T2�#�LO�sݶ�F��/�yq���'_>��<@]�E���pǏ�`a����ώ?z����}(*!a�d(Ù�Z[GÚ9{ո>�E.���j�?>H��K��;��s��Lt�rf9�J��d E:#A�R*G�Y�&��ڶ���g�5Jx������wP>|�7����lt���V��4*�I�xDBI)�-��VZ"%��J,wT��֏�Ns}'�=3��1��ىk�g��9>֑d$B*��L��	���Lgf�&�J*��͡wn_`������}��Kt:఍d��$�)L�EB�JgԚ*��*�%�EM���Z����M����_b7Y�m�LH�$$`d r�G "
aI�iۖ����f0l��P,p��d�$��`�ِ���(YU��H)(��ԢwDq���f���r�HY$#Y���Rnl7ނ�b�,��dI)ɒ�R��~�� �)�B�Pc\Dccl
���,2E��N�Τ4��Ed��ӧ��]�[i7r1vI�A)�HId���	"���hm����������N�]3Tmo�JZ��tq��)�@ʈ$%���H�����c����O����}}?�ӯ~olv�N�%��8�2	X�����w�2>�5��=O�GFK�7~��V/�ھ�G��.�[,�RʄȄLeBf�F%آ�;cu����y���9�e�ƀ-�
����Y��K�n"	ID���&�y12O�8Ai��_8��7�啣?�^�s���n��A>v���A�h��&�qȭ��|������~� �n2�_��|���N�^�k�6n����Rln<�Q.�NMP_�t��\n<1����RY=���=J�	M�P��kئ�J��e0��vYZZB�~��f���5D�"'M�rV������@r) sY}I=� }�'�+i�����ͰmgJ��M�{%_�35bNvpD��fK$Dm�MD`��^���@OҲ�%�T`�������4���DDc[�#b�6�l�fd#Fl��vee��m�v�,--��~FU�
�    IEND�B`�PK
    x�H5��~  y    _020_/resource/logo_32.png  y      ~      y���PNG

   IHDR           szz�  @IDATX��k�]U�k�s�̝�ә�L;��h�J�4�	B��
>�C4!�`bS|DQ> &|AM�	$�F��i�D@� 5Ŕ��(0��L_3�;��}������N)J��/�{Ϲ眽���_���������*�k�t	�m�o�z�F�!S03 B����T�=<��������{�s YO�}�&��K��@�� �.��>�[)o�*eg�K�LPm�y��
�Z�תs��ȓf�='�-Ɵy��>���ϿW ��d���Vm���֍ܘ��Gw�f8>���Z�V��%5zzJ��VX�bf
�>19����s���۱����2��+�`�%��[�,aм�st���km^z�0�<�*��.�Dp"1B$Cģ�\p�+W,c������i��}�>��w��N ��6[��Ncf��]�c���7�`��L�bB,&K$FA$�Q��{�<g��6��W�S���~��8�o��I ��>��[i��gˆ5�v�}�@������*�$�3�#"B��KD�$ �q�<Z�6W\<����.=2>�_��kp��n�����O.Z��;O?���(YVU�$m� $��(8� �$t�x��gj��b����O,Ԯ���۲�z��ظfh�/����� "��a&����$�$��1��J"��fơ�*�Ysd�x��I��/�f����|�=�h�iA2KDsA�qWT}		c����=��N�'��V��9�LLΖ���7�v�֛-�,�Z:LU70��E*1̀(�E|�X�
C�uHB��f4Z9!�3G�n4#�V���@R<�L;4����X'W{a�
�D��U1��T*�e"�h��D"�$��*��$�	#^��M� A!&�4G\AB��9��H��B;�e���v�"����'�"��d�ࡘO'L*��(U4�
&J��Ϩ�<�*��i��#�,�,=/�y�QIMk�⮈:*����8�{T���]�;)�(��q�|1Ŋ�K�uk������ɓu��ο�:�������t�­`Z )6�3����цS���J��R�>,����w��V��`W�)����Y��/�}��RQ
!�BҌ�"�@�XW׊O�֚;N������%��E�59��Y���� *x�CD��(�D�ŉ�a��B��q�� �]�{~�=y�辧��&��н�n^��f%������X����P)�x�B�SAb�BF����˛�q���^���  |���V�u�_�ۘ�����P�Q(H#)~��b�< �'�҉YL}8��{�o�y��?�:<�3wD=C���w2|����~�}p�#wiW�g�Q�{��1�����;@m���T�%^g�ҒPH�&!� @�	�C��I��vek��ru�%�?���u����W�~?+/��Ь�	���_��j�:yD��߰�9�Қ��`��S��1�/{#o,����4x6?s~�&B��C���^�����봫>��Բ��?r?/���{/8t=[����U[�o���VY�|&�v���n��t{��,ZO�i���Xg9u*4)�+�zzѥ��P�V��j���V���u��:���LNN266�<���h��Y=xwD�J4A�2<3�ݨ��3E��S �8��H�~�Q� ̉HCUD�nfy��P� �������婒je�'䝜y���wr1�!f�9`x�7�T*�<�c|��W�{?�ˁ0�i�8��}���	`�x6�@[DfoL��aU�˕W^ɦM����ghh����J��_}	m�ZLOOcf9r���y����'GD��N���    IEND�B`�PK
    x�Hұ'�:  5    _020_/resource/logo_48.png  5      :      5��PNG

   IHDR   0   0   W��  �IDATh��{�]Wu����ޙ;3���qlb'N�����$PT��٢�T�-mi+��PyU�T����6(@!
⑤Hcp�1��8�3�3�=w�g���Ϲs�v�����:��s�>k���o=��/�_���i��0#[ϥ/��{1�!�����_�����yl��r6��?~'C#c��)R� ��[:�^�N��S�n�����O���{���K��l��g��׿���_D�F��d�����N�N���<b[�ٜL���e�;�Nw�[�ǒ�`���f��{�(��g�wb�G���<���nf��ϳ���?Rk��~��l{�n���}�d��n�|ٖ��ל�u��i��N�����N�^���j5���N�t8tl�C���u����Z76��������#p�>��߸��7�����?�u�*�����yቕշ]�c��/<w�^�CG�����]:����V��C�rp���[7���6����3K�5��t�W~p������Ů�<}�{��=,޿�G7`b�<�-�Ȇ1��x��J���3.߹ut������Gf @��̰��;<�q,�9��Q�e�+K�Lnઋw0>�����óK�}���۫�[���o��޿{�7���K_�Fb��9�t�߯�rד���7�`�Dۛ)�T@ '����zg���������\��f�p�^e��W_v����I����v���&F?9�ˉ�9n����'�l�%��V.xޫ�.sK'o����<�����7����	*�d.*��6 PmC�[��P���B��n�E�ݽ��aa���/�n��[��m�^�������Et��p�o��'��6�����G�~�y��|��i�d"����X�^���`���q7̜p�-��=sܡ����	�����K�:|����{��J4���	ـ�������������_uߡN�{s(��B��3�I³���k�$0w3�r6@�{V�e�
D���l�"»�@�^vݓ�̭ߞ�<>v�J�\Z����w��p��?G�U�O���O��}g|zvɆ�
2�03#RH�L�L�0fff�d��X�oA�03E��fX�aaY�0�3�B	"��������+F�=��+6��>�C譶I�^�r�_�L(�Oݶy����]�f*0�a�0L�ARV�$d��v`f��,b@6�¨vz�j��VQ�a������;t�g?�����d��p��s/F���4�p������&�w�7S�&���"�)&��t3K^ѧ��f�|��\2s���f�ܔ�"�we(�����<_�ﻅ�,���SLs޶�o��zOHE���0�N�%��|܎;�=�p�!˓�e,d9L��<�o�,Ur��T��S�����,��&L���g
!����G�:9��J�}C��
�n���N��#��6[a.�[����3f��p/�k+Y�G�%#��VU�
#Ly5�W�pYx�!�;2go��� &6����Y��TyT�HH�=�i-��c�_�������*8�aU�@a�XX<��Ct{�s���Y$f��ZQ$"��K��dfD�)S��L��S�("g �ޡ R"����J�2�H��.�EM�"�K�ND(D�L'���"L�W�%fxdb�|���jQA�L��IU���^�#*?P�ó����"ˑ��E�G�]'��-��
"XY�:X���#3�"GA[͂锨$��\<Ⱦ��\9!��N%�gz]sT�fp��
��pX`$E�heej�Tʇ��U�|YeB�
F2����d�}�TB�*!��Zq��9��v��8,�c��Y��#��I�2W��g��>�+Qs�P�BT�p��/,\��0�A(�~J��_+�K��S��tsDXD���D�aT1���0պ��yKfd^?÷B�����K�) ĭB$�@� ����LEفe�O�		KI뜠L�e�d�ǩ�\����%ɔ�	�Pd�E_ɰP|L!tb�AP�:ķ*s���eTx(W(���yan�vXi�s���V��Xs�;qVy\-�E�Dx@#!�Vd�{��>��&����bQ-{@��jE�395U�M���ZT��o�,��8�[6D��c�����4ۮx#�[����^*e�7�:r��}k��V���x�p��,�LXVe���mg�mqˡb��3�8aD|��C������)��W��r�Z|��v^;���"2�rj�)r$iF�>�-en�W�W��j�~IΫ�5�	<�g��x�?Ah/ҳ��1|��,?4Ui��r�;_Mk�f@��A�~Q#�J��`X/�3IV9���8����$8͙��C~-�e�9���������v��_~�Kټ�>p-�:��N����	�����Yb-�R�Z� ��Y��ˇ��?}홍��o���K�^��P�Al0�S�W5�~�������yq%��3�+^;��z���ēe��g��W?�m�����Ӫ	�S���l�~>�.}�������̞;s�Q{.�I_�f�[DS�$���~�T�=����3s4�7�����#Q���/���_������a�N~���fr���+1�{͸����d&��vԅ,W�	P�`�DYV��D��O�a�Ľ�?¾�yL�d��y=��ד���Wʜr����R��K%9~�z�{�2�!�Q7�5"nB��F��Qc���<�}�����ɪ��y��L^�$��n�٣f6a��ʉ噖��\���r������y	���(�CHS��5�J�f������"����}w��%�3���\��`h|���I����&�"�|�j(�����w%�4�6B.�^v���V�������}w��8���B3~�..�ͷ����h/.@�)��f�*ϕ9f�\����r�?��@GRs�Ň��?|x�g��s?z'��	��L��H�͘}��L4��pX$�]~K�I�w�KF�ÆT27��e7�6a鱷������ѣG��X]sss;v���n�O��k��)W\�ƫ�������r��=�7�1)ӱ����#-+���CQ�Q��t�GI�-:�ҡIIQ�����W2ׂ�49r)I�ݯ�����㤔8p� ����ݻ۽{7�n�v��j$zN�p	ha�x#"F19%Q��7I�Q�y�W�����K�:��wत��Е�͜`=IaU�R�XYY����UyN�o6��
��	I��CR��TC/r�� &�A�i�ϙa@X���"��0&�g���������,��v�3EU��xU�Q�L4Q6h`JP����dN�p�cȞ��?^m\���ڒ:�1���nn/rp�{������7�$���$А��}��Qw���}�~D؜*������@_ '$ͻ{YAh��O�f��(p��j,�e� �-���=g�f�Ja�@�(#?!��K}t�)�����TyJ)jc���RJ\y啜}��lٲ�V��9�SŌή]�~n�!������Hbvv���y���y�Gسg��6�vŤ�    IEND�B`�PK
    x�H���.  )    _020_/resource/logo_64.png  )      .      )��PNG

   IHDR   @   @   �iq�  �IDATx��Z	tUչ��E�X�R},��U��"N�o�9!Bpª`�Z,�e�!�<�{s3�@�<ݐ�L$�ŧ��|
���~��g�{ϝ"
�t-�Z�����������������������~<��0s6M������kR�׿ߡ`��$���}"ݵ
X�H�q���14-`���5v��M�g�Ρ��VR~��'������v
+�(C-)�w�ѣ�����C��aZ������v����(��0��(����p�.���3��+�Ln;j!���Gc&L�ד�t����+���@��?��B��)��2��b�=Tv�������m}�/�!G��P	4��6���ַ����t��U@�.�>q��}MT�9����3�������.�,0S@f3yg4�gf;=��.��ĸ�G��+��-�i�����|3--������5'8�u�Wr}=f�Xc[Y5�ֵ�b�z�c����������9+{�KV񗯘	�Ʒ?c�o|̒�|�6v���Ԟ`��0��v�֪�ީuY���1�7��c�C� Fz#yf�i��
�v�����1t��?P���|�Z)4��u������N�3�����>�2����Nζ���^h:��3�b�:�c�y��Z���A	��#�d�XTA;�f�ej�}����K����f���l�A�ͫ��t]������Z	."��f&S}�\X�7ēwZ� ��FKK�1��Wc^��P}3�����{��4�"�R���Q�{R�L�g^) �{s�50��F���;E9����� ��g���gO�cĄ�<_���b@���!U�F�����G�kn������3����|s�	�F��~�.�!�xm����c�O3$.6��Z摤��Ikd:��H ��z�I1p_�!\����E�a���	���ʪ#,��β���avϟ��n��BD�!q�Ԋи�M�3�ݵ��G�/���;(���3��辣�������-l�	{`�����7��7M"����\\�c'�E��z;!j���w�V�ܰ��嵰���@�3,2��ݷe_gdA��E����ܓ�h�J��<���%�<F	��)F�qۼ�5���7$�z����3�Ӑ�~M-�/��1y�N+
�I��Iu.��9�3!�0{`{��R�'!�|��3��EE��BI5� �8k޹����X>	&0��)O<,�ǭ�� bUg!-	Kr��-�?�h�4�s��4�{YŐ�p*��\���}[�J03b�� ٽ���E�]g���>D����y��C���Q���x�3k���@��:��g�2�,�����?���T�N�p�<�Ȥ���v�=���M6��=g���nF	%��+�����?�ż��PP6�}����P�r^�噻юx���YI*0����,��s�EQ���B�r�Z=F������؊}�l�b��ʯ��o�@�t�nɵ4����l���H��J���E�N>�e�����D�+�>q��Yf��̖��q&��x�!�p�	�AT�K�{$QD�j�1$�	�Bݳ��*�}�"��V���j�12����n��"!���m�+�����{����8�F+��S!Z��nЄĈ" ��g����w؜?��0,�y�?z��F��It��( ����649�x�K�7j��嬻 nC����`��~.��QgBغ����P#D��>����xe?����p�	<<���f�J ?�~4f�ש��Ʌ���Ń3Z5�Ͷ��I2�,$od�s�9r9�a�l�D��Y"��ENز�m�< �.���?���' ҁ|pN�_�#���9��4H�fkg= �݁8��J����.���?G9WęvnȐcr&�MbT]�E�IN@� ����S��{N�d7�{b5Hk�p,a�ѽ��-a}ސ8�Wg��a,x�B�ѩق�S�+窂t8
��nq÷�`S\�4L+������{'�!���i����V�?+5ِ�6t�u❶����P;�i!\`é6n0�(�R"�>�Y(��Ķ*���0�����'C��VB��ežaQ��D�;���κJ<$ߖ4'�v�] �8i�]�;�ybDԜ��H�O��K�PP]0+��w��(�n#d���J��$<G�"�kI��`�E�{���9a1Tw��Y��ؤi�4� �o�U,@����Oj���% ���ţ��M��y�仅}Ōk�K����i�'-��b8��<Õڜ�K$�B��z�\0/� ���wp��/l�z^mv�l�ļ�<OX��nG܎p���E��m��i�����E���Q%1*%�K>����lswAhn3/��)�� .�@���y��-1�!gC�Wg��q���߂Hc�6�m�1~���"�;A���@��6.p�ds��{�z,���� ���˳̾��6	ϖ����*qA�0��HATQ����z\�"�{l��:16����.P�	�/@Ux��H�[����ok}m�qY�H>�ֶ����F�d��,��B��p!B^�&1JhB���.�Y\�4G^�,%����v�W���Jmf_c}k��1oO^3�8F�X�鈂";���~�*D���S�l�:�r�6�*�"Ⱦ�[��k�k8y�\�~���a2Nm�㯘ul�VI/,�L�X;,���
�L�,��|`	��\ +�YW�PygP���� �Dh�,�)���X�ǒ�,�/�κ$.Ȃ\l�0�I�m�O�� ��ߚ峕����
�z�'PJ�:�@����s��~�'�p��˄g�=f�J^!��b����E�GY,�X��p,F
��q��g�,�B�]�"*a�$^�����f�T��ăD��+)0��F?���Z��>'�ƼiБ<���l1�_\v�-�6�'�p&��	RX{�Yr�*�!M�-a����r��m�>H��hҬ�j� pBnǟ������K�ǘ��-�����lI�q|[�t�Ny�\`�eW����y��e��.�wZ��J�A��ه�'B�l�!�������l�yI�;`�q��pB��Ǐ9�0�xEa�-��n�>��i�@�C��Ri^�{�����+\=yE���a@��D����v����r��󸎕�,��N�%�'����|��A�	�\`��UV�`�<`)��;t��#�+��|2��X�4E���b�#־�qo-}J�gk�!��U�s���񝯳�]
�6�gA�8�k)�|,�y@����-�����_�G�n���݀����!@7!�nC��=\�6�O&?������8�V3��N���7�R�-)WBC8"p�hÀ�[�jIT��Cg���!y�� ~y]4y^��o�t	�(��O���x�k��m���5>V��Ɏǻ�i�:'��� ߎ�"��.���Z��V ����S t�k����?���xhݷ?�K8@��!
�N(<Lxxٿ� g�އ<@�(<nY�ԹC|��hᮓ��KH�Y�e�?�o��-�Q	�����!���ݾ�o&��CQ�8�h�0��B�7bp�\lI0�g�uC�_�.J!��n��h��������r1�V�IQFa�#n,����ER���/�/w�P@^������wB�o���7�R�i� 1�o�7B�����L���x��Y��(~�v�?�(#Q����s+\z��p~�QT���S�(Y=e-U+r��t��?q��K�����e1�H%mYae(��Z�����%��� ��@y�,���@8F�'��4�����0r4�&��#
z	��t�\���RX�VJ��*�w3�g��m:rf ܗ�x�q����a�.=Fw�@E�{W'�t�5���W�\Y��z�g4f���!�s�P�'b?�<Z��t�i���6��y���yOS0+���5)43�1�����+�I?��a�7�7cm0��Q �=�c���ί�LB�ρ�X��XN���*NҤ��\����	Ȟ/Qp>O*H.�|i�|q�����_������x#c:�q��H>�]$,Q|�"�S0Bi�.�������SP�	
�>Ŀ-���v�<���o-/GP�!B�hL��!B�~�E��{��y��q�EfZeh�g��PM[��)]_B�z=򩼤�***����{�n2�n�:Z�~�6l�@k֬���
�����o���M�F3f�p$Lp�J�VPF�����n}Z��5����n��~�=C�y�������%��<\к�1}��o&?o����jZ��O/��	������/�<��� m0z	�y����%L&����`�ΝT^^.�E߳gmݺ��/_N���H2��H)�Ŵ�����w� �������%�K��/�"[o��/�:��0!��xm��x]��0� (4�'��$�A?dof�b���ր{p/�$��)0�
��1p�#�˝�X\\L��
W����~
?������R�A�)��E;���6 ہ, �<�%�������0�b���c4D:��̒bN��q�.��U& ��������hz�!`X�$�.�>����3�Y�����w�X�qɱ�ȱ�\�$��I�T���e@&PtG�S�;�_���`>�������|�C����o4��J���y_ʱ|*�vF���r�$�N�-Sr�/S�cf:0� Vk��@���e�T��נ0�vn9_�{��3�Ϭ�c)ь/G�y��Zr���K�$����Q��8i����3eb���)[nv� ��K/��=�3쟫��/5�s��u��8�m��F��h�ڵ�,�QVVf)��ؗM�\�a��7���Bb���(϶dzN�~�*���R�������~`�ԩ4{�l


"???Z�r%=��s����3�<#;.Jp�۶mc�c�x���ח��ݝ�L�Bcǎ���Z�l����    IEND�B`�PK
    x�HI�,  
    _020_/resource/user.png  
            
���PNG

   IHDR          }Jb   tEXtSoftware Adobe ImageReadyq�e<  �IDATXíWMLSy��{^�=x1i<{���Wu�f��hz��6�1�5�*�l������Pڂ�
�C�Z@��~@[k}}������Y*-��L^������3��<��{���򧥥�s�p����Mu����q����UO��5W�h	�K�6���i���n��d2(F;��u6� �L>F�؊�z���'(4㖇�K��I�ҭM+�|ޞH$��D�J����w�LU�F��z�fڇ�>G�J�]X[y-�c����)�b�G2��ݶ�f�a��F<��n�EM[���7�P�m�ߦ��CLMM�5|��^`�6�޻Z��(���4v�{�8��e�#����� ��b�G���Y-�Z��r_���6��2P�t(��Z�-�{L黃T��˜�#G� ��s��E��q�r9)��g�?�M>�uJ�^]��ݻ��X��������8{�<�OC�m�����U�{�N{��d�VWW��f�|�M�n�|n|����^�s�,,,����}�Ⱥ��(g���ëW�����3G�y�/x����p!y��`q�J1� K�N^����'z%6�WHTy\HR�T���}d��3v6sW����ᣒ}>�c;F�=uF@��%ܥR�^� 7�ρ��7i �~��K?m�J9k6���?k�o#�%Ui�Z��I�w>��\��
�Ү�L�&�	�-6��8uxXkee����,�#/fY={V��%�L����l�$���Ɔ�>G�:sF~3�h�(���U�077Wj��n|MJu����h@���8l� 0_���K���������^����������ݳհ�H�oe, ��񀱀U�6bh�P�=C^3�}�3�uz�t����4S�YI͆F7y<.ez�!8�btc��(�������tq磡A�1[<�%�=���~�CV÷��ߌw	6, Ʊ̇���e�T����,��`h�b� �����6S?0	3	�;�X���a&c�db�.p��庱aG@AX$�Z�7A|Q��t*���1�E����jim�s�PF 9���gq�4#*No�c��<������5����mǎCSS�
<a���L�0����&,�+��={d�'ʏ:o�]�8��YB������. z���v�`�������ۧg��#؏=*<�R(��,��~A��SH]��e����B9 �n����3�ꜤK��e�*�,D#�<�F����M ���O���3�\/򙰐@�X�~'����K�G�Z�AM���C>���ڵk�����j 4Ʉ���=B.�����T�hyy�>}����4��'z���q��U0I�j�D�Fҙ�+�EE&>Ya3�w�W�O�~s��!?�H'�X/
K����P�9��r�}����Т�v���Ifj83�Q�沶�Z�h�]����J�<    IEND�B`�PK
     	x�H               META-INF/services/PK
    	x�Hj�R�0   .     META-INF/services/module.Server  .       0       ��/)-�J-���K��	��Ћ��,��**LKM�-�O��M�p��� PK
     x�H                      �A    KOtupZesZNNfLlSPIX/PK
     x�H            +          �A1   KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/PK
     x�H            	         �Az   META-INF/��  PK
     x�H                      �A�   _020_/PK
     x�H                      �A�   _020_/resource/PK
    x�H3i6_  �  4           ���   KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/AUX.classPK
    x�H�I,9a  �  4           ���  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/AUx.classPK
    x�HZ��t_  �  4           ���  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/AuX.classPK
    x�H��7 _  �  4           ��G  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/CON.classPK
    x�H%�k�^  �  4           ��  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/COn.classPK
    x�HHY��_  �  4           ���	  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/CoN.classPK
    x�HL+Љ]  �  4           ���  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/Con.classPK
    x�H}���Z  �  4           ��X  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/NUL.classPK
    x�H=`�^�  �@  4           ��  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/NUl.classPK
    x�H�+��]  �  4           ��"  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/Nul.classPK
    x�H��-�_  �  4           ���#  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/Prn.classPK
    x�H��3^  �  4           ���%  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/aUX.classPK
    x�Hx�8�`  �  4           ��O'  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/aUx.classPK
    x�Hb���_  �  4           ��)  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/auX.classPK
    x�H�d��`  �  4           ���*  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/aux.classPK
    x�H|Tx�Y  �  4           ���,  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/cON.classPK
    x�H���^  �  4           ��_.  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/cOn.classPK
    x�H�*�_  �  4           ��#0  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/coN.classPK
    x�H�1��  *  4           ���1  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/con.classPK
    x�HQ<�^  �  4           ��A6  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/nUL.classPK
    x�H1�2��    4           ��8  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/nUl.classPK
    x�H�J	�^  �  4           ��:  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/nuL.classPK
    x�H��^  �  4           ���;  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/nul.classPK
    x�H���\_  �  4           ���=  KOtupZesZNNfLlSPIX/ZyYvkkRrqfefSmwkWfZMexC/prn.classPK
    x�H��ؤG  B             ��]?  _020_/resource/1.pngPK
    x�H[���w	  r	             ���G  _020_/resource/10.pngPK
    x�H#o���  �             ���Q  _020_/resource/11.pngPK
    x�Hw�B	  =	             ���Z  _020_/resource/12.pngPK
    x�H��Z�{	  v	             ��$d  _020_/resource/13.pngPK
    x�H��i6	  1	             ���m  _020_/resource/14.pngPK
    x�H�5>/	  
	             ��cw  _020_/resource/15.pngPK
    x�HD3��  �             ����  _020_/resource/16.pngPK
    x�H�d���  �             ���  _020_/resource/17.pngPK
    x�HO�0               ��ݒ  _020_/resource/18.pngPK
    x�H�%��  �             ��>�  _020_/resource/19.pngPK
    x�HSZX	  S	             ����  _020_/resource/2.pngPK
    x�H:��  �             ��!�  _020_/resource/20.pngPK
    x�H�m.	  )	             ���  _020_/resource/3.pngPK
    x�Hl�4��  �             ����  _020_/resource/4.pngPK
    x�H��]3�  �             ����  _020_/resource/5.pngPK
    x�H�4��)	  $	             ����  _020_/resource/6.pngPK
    x�H�5��g	  b	             ��M�  _020_/resource/7.pngPK
    x�H�?	  �             ����  _020_/resource/8.pngPK
    x�Hbȩ$O	  J	             ��D�  _020_/resource/9.pngPK
    x�H��\f  a             ����  _020_/resource/admin.pngPK
    x�H��4��  �             ����  _020_/resource/logo_16.pngPK
    x�H�p�'  "             ����  _020_/resource/logo_24.pngPK
    x�H5��~  y             ��5 _020_/resource/logo_32.pngPK
    x�Hұ'�:  5             ��� _020_/resource/logo_48.pngPK
    x�H���.  )             ��� _020_/resource/logo_64.pngPK
    x�HI�,  
             ���. _020_/resource/user.pngPK
     	x�H                      �AW5 META-INF/services/PK
    	x�Hj�R�0   .              ���5 META-INF/services/module.ServerPK    : : )  6   