PK
     +Q�H               ACvqqLVUSwkYm/PK
     +Q�H            (   ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/PK
     +Q�H            	  META-INF/��  PK
     +Q�H               _004_/PK
     +Q�H               com/PK
     +Q�H            
   com/smaxe/PK
     +Q�H               com/smaxe/bridj/PK
     +Q�H               com/smaxe/bridj/linux/PK
     +Q�H               com/smaxe/bridj/linux/lib/PK
     +Q�H               com/smaxe/bridj/mac/PK
     +Q�H               com/smaxe/bridj/mac/core/PK
     +Q�H               com/smaxe/bridj/mac/core/ns/PK
     +Q�H               com/smaxe/bridj/mac/core/qt/PK
     +Q�H               com/smaxe/bridj/mac/delegate/PK
     +Q�H               com/smaxe/bridj/mac/lib/PK
     +Q�H               com/smaxe/bridj/win/PK
     +Q�H               com/smaxe/bridj/win/lib/PK
     +Q�H               com/smaxe/uv/PK
     +Q�H               com/smaxe/uv/media/PK
     +Q�H               com/smaxe/uv/media/core/PK
     +Q�H               com/smaxe/uv/media/java/PK
     +Q�H               com/smaxe/uv/media/java/swing/PK
     +Q�H               com/smaxe/uv/media/java/video/PK
     +Q�H               com/smaxe/uv/na/PK
     +Q�H               com/smaxe/uv/na/lib/PK
     +Q�H               com/smaxe/uv/na/webcam/PK
     +Q�H               module/PK
     +Q�H               net/PK
     +Q�H            	   net/java/PK
     +Q�H               net/java/sip/PK
     +Q�H               net/java/sip/communicator/PK
     +Q�H               net/java/sip/communicator/impl/PK
     +Q�H            (   net/java/sip/communicator/impl/neomedia/PK
     +Q�H            3   net/java/sip/communicator/impl/neomedia/directshow/PK
     +Q�H               org/PK
     +Q�H            
   org/bridj/PK
     +Q�H               org/bridj/ann/PK
     +Q�H               org/bridj/cpp/PK
     +Q�H               org/bridj/cpp/com/PK
     +Q�H               org/bridj/demangling/PK
     +Q�H               org/bridj/dyncall/PK
     +Q�H               org/bridj/func/PK
     +Q�H               org/bridj/jawt/PK
     +Q�H               org/bridj/lib/PK
     +Q�H               org/bridj/lib/darwin_universal/PK
     +Q�H               org/bridj/lib/linux_armhf/PK
     +Q�H               org/bridj/lib/linux_x64/PK
     +Q�H               org/bridj/lib/linux_x86/PK
     +Q�H               org/bridj/lib/sunos_x64/PK
     +Q�H               org/bridj/lib/sunos_x86/PK
     +Q�H               org/bridj/lib/win32/PK
     +Q�H               org/bridj/lib/win64/PK
     +Q�H               org/bridj/objc/PK
     +Q�H               org/bridj/relocated/PK
     +Q�H               org/bridj/relocated/org/PK
     +Q�H            "   org/bridj/relocated/org/objectweb/PK
     +Q�H            &   org/bridj/relocated/org/objectweb/asm/PK
     +Q�H            0   org/bridj/relocated/org/objectweb/asm/signature/PK
     +Q�H               org/bridj/util/PK
     +Q�H               w/PK
    +Q�Hc=��  ]  1  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/AUX.class  ]      �      �T[S�@=�@ ��MEl)�QK,X(�T�LHw �dK���C��O>X�q|�G��/(��C����|�����3T�2���[��M20�(#���C�&���e���w<�Z:/	?or� �W��4C��>�6���|��<��m�(z�.�p�����"��X��y<���7k�P��"m{�[��Mm��������KW<+kywT[�(w�����%�
)�U�*�SP��A�y�ޤ)l͵�=������L��Z��p1�7l�Cɓ�E	9Ȯc�?;���a��9>�����mnz�t��ޏ.c�g	'�����Hx܎�P�T�JJ�D��&t�8��*jХ�
Wjq3�A4�a-��%tK�pUB_��Њ^	7�h�u��.2����0�l��[�F�/K`��b��S}��I������غ��o膭��<Wp'���&��cZU�����2��B�1����L�,wҶ��-͇Ÿ�<�2��܅�����>���N�,���U�_�)�i�$5�L��^T�m���g�e�e�)��uQ����	��i#���=�7姿�c]{CSIQ�zHM-�8�(S�Re�����#�U��0п�<����#�(�[��df��L��zTS8V�(�׈���^��h]��K�(A[�|K�d�����|sxx�������>���m���hn�W��Ms����n>�����*a�W]-��y�Y��0.�PK
    +Q�Hܧ��!  y  1  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/AUx.class  y      !      �S�n�@=�K�$��--Z�rkn���@
!�T܂�&$y�8K�؍c'�O�xF
E���n$�@[���̙9{V3�|��1�әC$�������>e`��s�n��m����y�Y��k�>��i�6�v�G\�M����͎���#��p�+��qlg�ǻ)��̠���u������>2�٧ࡂ
�+��`^A�!��?}�a#��A>v51����U�(U��=N�Uס"�WS�@HE�1���P�!��1,"�.��R˸L�X�;�$�mk�r˭�G�ҟ���6x����{�H.k��+Ct��aG/�G��^�U�o�}mpl���h�}���Vލ�{��aM�y��P��RmBy�ҁ�����1��[��^~ie�N ���'i��ԭ*���\ ��$7 �����آ�Z�%SH#�k҂�\���GH'��"�	a´'��V�3ֿ`��7hݤC9d|_��j�vy��_j+�R*����b}��)�L���8��HD���G̿G��Sl��[=�'��?�b�I1�PK
    +Q�H�:�k]  (  1  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/AuX.class  (      ]      �TkOA=��ˢ�QD�*����Z[�`ʷ�2��vvg[�_� M���Q�;[I$J7�ٹ��{�kf����^2$��"C��빊d�L�`�&���;��AUn�����T|O2���ê8�<�q2��;~ y�ݖ~>U�@{�&xM��A���Zw�b��A�r+��9QHOq�����L�y/w$i�2�ч<���.ϔC[&N���*��[��6�=,Hxa������l���i�	���>�u{G���+.k���aN�cD�=ـTձZޓ����9�
���|�ЗY��ЂL�Իa��t+�.<O�ϒ�������H����A��!���4�ά�Jx�(*�=箕�#*E����������]��@(���k��*?��W���\���1��·��Q}w)���l���j�/m��+��@��9`����U/���Zx��t.�謮4��"�@S�M����q����5Du��aFK��խ;[ɏ�2M�"�:f���?c�S�Hd�O�hL`�1�c��v�`�.�٘�CgTˤk�o�zKS�?��c�9���}�}��D��y�{"4<�w>�A�����PK
    +Q�H�]O�*  �  1  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/Aux.class  �      *      ��MO�@����"*^L<x���5&�Vb�^�*�6�XZ>
�+O� �qZL��0���Lf�����	v�J�%d*Wqʝy���	$ؓsOv�b&L)S�d��{/�Q�+�J�	���A�l,&J�()��p�=e9a����̎�i�5��"�G�<V��sXaW����v�'ھlƁp�Ԭ�h�w��50G��s��f����ͥ��zu�ڬM�܄ڄ� ��+<i|RE����&)�z:�zxE�5a�cy�c[	�#��i����O�=x��j,M�PK
    +Q�HqpCo'  �  2  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/COM1.class  �      '      �S�nA=�Е��@mU��jE�ڑ��5!
ؤ�J�۵���ewaѧ�L0��� >����&t7ٹ�g�=�ٙ?�~P�c�@�^϶���������W0,
���ڮb��U9"�ː�u���+|8��ҕ���nd��NبBUj�(,�ĉ�17�v��]�2H���2,��u!;��#ᑄ�H�/A�pYB�!՘�\b���\쮔=dX�4���-������U�y�ٷ�iF_��=� '�G�� �egv5�yl��b��AD�B�BXB"��3�+���0_�5����!}���w@]��0z��W���auV�����bP���F�2��{����'zK~nW��;���٬U���;��\֛�%/�W�"T2�$���t��2�2l�7ۮ�*Ep[�\�Œ#u�)��P�b�C��!���'r��u:`KtU|ј�u@4A�.�ᶃ"L+�b��[�<��V�p!w����R����)�0�r.�Q2w�ǆK�ʔ�E��G1�� 9��	V'���N��7�1gX��u~���Wwν�i�N�~PK
    +Q�H�H?�  Y  1  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/CON.class  Y            �R�NQ]�ޤ-iA
Z��"�FN|FMj-,`Rl>�N���Μv�S��/��K���f��G��&bDf_��{��O�����C(_8f��6mS�e`��	��0����y�Kvm3�1�#G2���%&����ܓmCX|�x"�Jݐ}ih��ђ����͐퉱�p�3�.��]�X%�cȜ.�V��V��$2z�-���zC9�1$bH2,����dX���H7��ʑ�iv��r�%�1�8��4�cik�s��o��D����{tf�Іvh���|��5�$�`I�0��4����4R(�1��8�p%�4.�&���=�LUٮ�n����}P���)�}y����e����t�� �F�R��棆����Þ�7�{������@�{[�g^w���W�i�I��E������k��ty��p��0���ق
��U�Qva���q���a�R�dW�8�(XQ����0��Td~QՉ֧Z+���[�>!}����V�=V^R��*C��M�1�~�:��PK
    +Q�H�9��a  -  2  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/COm2.class  -      a      �SkOA=��KQ�(�@Y^��[�����#����t�bwf�-��L�&���(㝭�$m7ٙ{�{�c������9�dH8;���E/�4�l�~�pM���M��B��]����rH���<�ű�*�cOp7T��].+��_:U��t�L�Bu�к/5�t�h�L�[QJ����3��F�I��eȠ�yT�}�)EZ[&N����.x�W*�6��,,YX��`ᅅ+�:,�f�MD^`�p���Âi�S�5�eՐ�3�9F�9�uHYP��j
��\�niEE����B7J�,��H��M#��K�����$��,�<�ы�f�я�����Q6ܥ��̆A�E��\!}�_E3��CW�By��g�,��W�4vQ�P*���L�zt�/�ݪ�/��� \w_�r���C�-�Nj�+��T�ڼqtMFY�9�˛��fR�n�����3�ըצZ�����:=�F��L3�57Mi"*c43���Z��0�VP4��jW��I|B�!:�&m	:�_�[�:��)���&���3�sL$��wg���Pt��=Ў���N�,���o�%����13�3�	���C0'f�QL`�vJ��R���PK
    +Q�H}w���  �  1  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/COn.class  �      �      �UkS�F=�6gK�4--!I*�%M�CI���0�4m���X���&��_ҿЙĴe&? ?�ӻ2h���sw�={���#��?� p���6SRז{�"��˱��
N^�)H���/��#h�(�6-��vN|J�SA�tmݷ���ön������߱����dՄ�fzB8
�ΐ�wD�䶾�Y#�\��qG(P�Q�6�&�����]�&<�?q�@��+�\ȭ��T�lr��X��+^�Z�W��49��j�똡���:\�2�ldVE]��G)��;[����-n���y!5�mu�pA�y�rM�Ŗ�x`�D��q�ƫ·��j���a��%˷ȯ�UᨰU4U\R�T\V�R1�bLś*����y���_Q�>���W�������v��u��ޠ���SQі;��^Ĺ��#���ԝG��㺢�Z��q���~���tv�uh���R3ġ0LH���wcxW��exs*>f���n1��6�$>aħ�x�,	�aL�!���5�$�%\�|7�Y��	�%�~�o���H����𥄯$|-ᎄ{�p��snM��pM�,qϒ�[�i����s��H�m�5M��=���$��$��%߿9#�k������n���v܂��ɇ�KO��_Y�?�4�r�BhP�I��Y�+J!?��ڨ/MK9��a�����ŷ���Rc�����.@8���+Ҕ��z;��oЅ��ȅم���žr��{�nj|0>9��t�TI2�@jTv�����3����)�I�,���<��lg�c�9�0� ��-�i
� I��F0Li�h���2ݕh.��N�� ����P0ҙ�v��ϐ�t��T�rk��I��.�$�c{��.��[]<���(r�/��w����Z9}��.�?�t�Rޒӥ.ֻ(��r��I�,UD���/PK
    +Q�H�}"�*  �  2  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/CoM1.class  �      *      ���N�@ƿ��"E��x��X9kLH��X��U�lH���Y��V�4| ʸ[L�w��of�7�v?>��԰K�*U��W�Tʜ��/�e�}A���X,,�ࡰ�����>�>#�々���>&���Ds?(H��+���O��	dBG*�5�9䐗>��	E7��c3�u�VA��k ���c�n/�S׻mţ�ؚ���E�<�O�D̛��24�kˎ�51����Y�W�T���.�� Q@���R�d4WM��H���7p"��YM�ܿb�)���VL�J(�9_PK
    +Q�H�����  ^  1  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/CoN.class  ^      �      �TMSA}C+q��|���	W�Oj�!Z���i�L�Bv'dw���п����*˳?J�YPQ(�ü���~��5߾�`O�h��Cøi����J/HZfhZ�n�h�I��.C#��W68C��Ž-��j:�͕UwNx��\Wؤ\�+��W]-)�������K�+��|�DA/����y�5U�=ۥmSs�����>%�4�m���a^��,���Ւ!�*8�tVEU�c3
TM
�(hV��0�1��9���5��Y�`�!�\˙.�˺���1�9\X<����=`�����/,1�E�{7�:U�ty�.%���Ye�pMaǣ(ge;�.��*0�B�Sъn�qA�)�����F�Ŵ�Tm�
��C8�>	�.I�B�4t`@µ:q�z��������2Q�G����fVw�
Ow��|��-wB��I��t��)#���˦�\���$Ǧ��C#2�I$+�܋��z��6�D֘�����7����M�^WWf�O4�i��.DN�p����̌�PI
I%`�n3L���=��9��Iqt��C�uo��)?}M�,��N!�~�v�d�Z�25@;��5a����Ҍ�Ӿ��04Q����@�-��±����O}��t�qc,8�\�A[g0��l���{����˯8�a���F>�1��Q'�� _
�>�	��>�q	��<4��*����ۈ��Gf�3x��R�|)H�Q�PK
    +Q�H�w\�i  �  2  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/Com2.class  �      i      �TmOA~��rRhQA���V ~�
��Ԅ�Jkb�=Vrл��]��*Ml0���Q��+����v��ٝ�gf_~����2V��|�A7��we��=s<'|���:���<př�Q��������W��o6�+̿6y��e�./��q�l9A(=�dp��,-�Y�H�o�I;dW�3�2�(�:'td�`��u^+:�u�:n���`����w�aъG�V=;j6�r��c����IV[�3��UM3�뚶#���Z1�S"e����%�KYa1�a��"��,Fp�A+���˷E�"�����C&�NT3D?��iҋ\�%k��:=�*{;���O������F���i�$^mn|ln�^yw�*K{��pf&�+���Z�n$;�����s�k�����،�������j��n��M�1˰�C�V{خ�a�nl�x���U>���	�`�\?�P�]S4�&d���WL|&���F���J��/��-E8x��j�x���0���q��H��kee"��e�}�4f
�Z���������~5�U��`�x���u�I����8��2T!�5�jLŕ��Y�zфz�X��Y[��~EQ�R~PK
    +Q�Hb��K(  �  2  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/Com3.class  �      (      �S�NQ]�J�Q
jo�ӂ���I3h	I��};�����N[�S��M*&>�~�q���1�L2�̾���:����߾(�C0�n1�R�t�a�a�Kv@/g��k�ֱp�ڎ):�m3dt�T&?�p�����)qu06��zP7:®�õ�p�����^�w�2�|�Zj\�8J��2Ø><��I�#؍`6�C�ru�"�Z����U�HX�zIV��E�zi��ㄮ�!��(��8
�X��:v��C>����G.�ܔ˭q��Q�;�$k�5p���yoH�������y����{�D.+�;+Cx0<�v�����J�um��i��S�H5.O�?���Au��~���Uݮ�H�.O����.��?��$5���6��\��9*JЖ?�f�P)��/�54j��2~T�H���>4�*n�A}�H�H$IV��%1/oԋ�#C��^PN��x.��~��W�&����b�!����|m�.�¸�ҴT�Jh�g&X�`e�;$�0.p�#�f��	�o��f�k���/�Ē��9O,)�_PK
    +Q�HS	R��  2  1  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/Con.class  2      �      �Q[/Q�F��[�����'IEҬ�x@���v�,��Vw��W�����Qb�ă�dΜ��7��7����`˄Xv�H�ڱ��%��W"tU�a��[ޙ�o
G��,����0y-�R��f�t<qi9e7ȗe�3o	=A;֘�r*
�,*XPХ@!�����3Y����ϭ�� ��	J ����M ��$z���F���2���]CV��֒��yV�?o���B%�z^k��z��,���E��=1���~�P�y����}P9Ў�v��"������ >��(}N|=��>LǷӘC/a-QЧQ�<O���fBi�u��םa��-�8��WkO|��c��(����^�����]�j���[h��Ä�,���,c��'PK
    +Q�HmzK|Q  �  1  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/NUL.class  �      Q      �T]SI=#f�#��$d����(k26���]v��`2��n����_`�O�`����W��9��z{0~���9���{����/����ݑh:�U��K�c{��"�Z_gP	s�f�-ϭ3,sϨإ���;C/�9ׯ�8�D����d�7��o��<�{���amY���tí�\��9Fޒ|�=P$֭��iE�c��V��m�Ѵ���xͭ��%����;r�]�=�7(���"ȂS�R�۔���"#'ㆌ�2��X���8(㐌�2��^"���Ӣv�����i���"ѽ��E�^.n�g��ӵ�I�<�u��w�E�v��ո
LE� E@7�T���	_a\E�T�׽8���,)0$ ,`X�&`
FqZ�g��	�"��Qp�TQ�]��p6�/��W��ƣRGצ�ϯ�7yѰ���_�2�(H�*]�O��nT�-Y�U�n[�
_�p����ݙ�$�����j>׼kV��7[�k�����R5��4���Y^0��ƲC�MG:�Se�N���3�L�Û*�3C��WڏtUqFE
��/���:�.�����J's/;D'�۝D��dI����������x�+^���&B�-z�ę��=�r���W2��r�~����`W���,`�^��Zv�O�������$f���!/cf�_n���C��͛�/��ϫW�q�o<�Ř����]h�-�`N��|���m�&�֤.�bP���t��b�-��Ӂ ��=��� |�M�乀�ڤ��Y(��X�������������%��/H�H�AŠ7��7%8'Z��I3�S;8��^y�WH?/��PK
    +Q�HCQ�$  �  1  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/NUl.class  �      $      �S�NA����� mԊ�(b/����jRkK�k5���tYI��K�ҭ>��`RC���g�&�`jv��9s�;��Ι�_��������F��b�<��]�{I�`���5�����05�����bh���P�΀낻jGo��3Cq2`�n
M���2Gb ��r��!�t,ۤ�?/ì��g��Ix(၄�$	$Dr���e��欺ra�a9/{�pm�T���j�]���0F���m�T	��%Âg]�b����fs�Q$�C�c�G&��0��Ɓ�0S5t���=��K�0�eC��0���Sw��s��D'm9Ǫɰ!W��~_n�n���M�[sv�>Վm�u���=ܪ���]ًS<A�����CJ0�r��T}��A�erd?����;Zwq��@i � M�vd�����JfP�nx+ē)���,i�:����B4�GȎpm����@����p�]rH�	��a%��/�d�I��i"X����X#��c�䛢9�^�/}E���9_\%���"$��V���PK
    +Q�HQ#\Y�  
  1  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/NuL.class  
      �      �V[WW�I�����z)Ԇ@��V�V���! 4P�����0�I��[�G���G��VV]]}�C���/h��(.1�Μ=_�}��g��}�,~`D;�B�dR���e���/��H��';��|Uh^I��V�k�[��{9�c��y1b;y�")G�­싕͘(yV0(�I��i��e�sW8MK��5��&�rӮ#��5ǭ�6�j��k�C��u|aI�q�4�Y_ȑ��=#	�Vv�3s���>��Z���7y����2<���q�Λ�6�/�� ��TzU+�IU�6�l�[����7i�S�i���Tm�<����JA���{�#l(޳˻��b�e�v��
�R�/|� ��N��
�4(hTФ�YA��c
Z��gJ��&��w�<m.
;m8BX����W�(-�*D��^E�߬?�:�ꐹ5�,a�����N��B��DZ%}(:�??�;g	p�&�L��aܤn����0}��Ĳ{U���?�%��]>/�Z��l�����AU*ڠ��I�Qq�T�x_�kޖp}*��o༊>�𑊷p�'p�'�&aUBYB����)x��Ў�:0�����G��e	W$G��.�DЍ���|"aHB�:*a/R�5��s��1役Y��3��9JY�|oo߼F�J�|�\�
�D�AM�<���Y��A�Y)�#�E��ִ�¡~�&��������ќ.z9���`����OO��˙���d��+�a�����[^+gGש	e߆���:(,�fX�]�H��I��hU^�L��f�lFeX����<�ܫ]�Z�;���zU�ѣ�B\��%����W����`��*�Wl* ��$&���0��k��M����s�����G�l2�o)�7��{�֓ԝ�!X� s �J	�Wʎ�RZ�GM=}b����h0 �ۂ���xwl�kW�qm�u\���Cz��a1kh����:�!E�?)���%��)H~���M���&&�d��&n��#\�A{��]fn7��M���T&ֵ��m| qd�g�1[��؟p~���(���laaf��ۘa���nn`�H��mA�cw&��|P*e·Z�?�7�:w�v�΃�N[���TE�%�����i�L�-d����G����	��n?� ���ȬdM�a�	eCf�PK
    +Q�H�u���  �  1  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/Nul.class  �      �      �S]oQ=JWp-��/Z�jU>Z�>��i$����"Z}0�ˆ,������H���(�\��&>�;s�̜�9;w�����C<`��-��ǎ�;L��f�R�?G6�|`w�{b,���؊���{b`ׅ�w̰2;�?۫I{8�e��Ѿp�|�ݳe���z��h�m���s�`?��	IH�����خ�χ]��}��1lZ��T*��k�2Ò�{�������Y��Z&b`&�ڜ��$Ll%q�$�P�&�BWR��r
Y\bX���Y�������y*;�C�#/��ӷٶ*��hd�^�O|�S�tR��k��Y�O���\�oI�N>�d�x&�4m����[X5q�Q�U�(kRQ�WJZF�&��i(ܤ�eA�A,�ժ �$�~�X�!E1�z{B����fX�0����~�����	ק�	��J�gTt=4�C��.#��_�*H
����ޗN�v��ϸ1%蔺Aa���������8��Q~PK
    +Q�HB\�%�  I  1  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/PRN.class  I      �      �T�NQ]���"�p�mG���ZX.,�������i�����D����7���¸�@(x����=g������+�~$|�h��YRpfȴL9��&��ܐ�m�
g�v
"Gl��!f��X�BwK:�L���׋e�Z�'�fN��#���}�c��e�5xA�X���9/�"7!1a�Y����W���ǣ\i�uö�q�%u.�i�q�Ĳ ���덽t�٢t���WC�A�d�.d�Q{���(dܕ�8ϋkN�M�(J������>�����aTC\C������z�440���t<H�[�^D_�x���R%U�n�I���4G���^�dW�It�-r��s-�g��;�r�2/���#G��I��\��|`!4*FMgqQq���\�f�(�4�ъ�J\�ה�D��:	�<n��%���>a[�aK�yޥ���z�Д�i<i�%�Oqjn�p��	˥�b�L}�x����J��/����U{�xVN���5Y�K�)��'��s���}�TR�o�_�c���4N��{cz� .��]�'M�r�kv�:��L�|�F ����x?M�	�����%�D-���'Dwp��2S��Z��#S���*Z	{3~�?�r}U�g�h��z;�}�T����9ax@��Ch<-��`և+{aS���0�[��n#��X��^b^���(�	��Qa5��R}�PK
    +Q�H�Yq�  �  1  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/PrN.class  �      �      �UmWW~�$.�[(��-�V�$�����/E76X���.dwþ�cI�B��Жs���z:w��I>䙹3s���yn�����|		-S���;�"Ĺ��k��I��ZMB���E7� �.���dZ�ݚ�:�IU�Y����Þs=��^�������l��?,�5�X>箄�S�.�[�j1G_\���u�=�����%�d(2���8+k��ϯq�`/�(�0��.62;�.�*X�ns�M\l*E�˪J���Qh7t�s����d���c[�L,J|����)�u6��u%��ڡ��#j0p:�
�,�bQ#�7��/5��Bۣ�rU��^���SK?-W�P�
�e;��.Ó��pd4d���ʸ(#-cPƐ�K2.K7�ô�1�݃��	����������$�qU;�w:/0���'x턗�Nq/���V�i2�AÇA'f�/�;VB��c��V��Nv�4=�Λ>+��$$���O�GH��X�{W�!&Tȸ����0���T\�]��� >�� [�/A]���Qpc�aZ��S�)�����by�*Є��s_�R�W�p_���q�ēy�FܺuV�g]ѥ���{�:1"Ϝ<k��Ol4T@�~��,�(3��]�P8DM��RĘ�~ǘ�����'+���w���5ۚ�V^�5à0?��U_�?"�9St�3��=�T�w����~�
J�����u	���&�vRS�r*�aS@N,�4�F��md�?�۬�R�^z��S��Cr*����}=2�Fo��I<!^�З�$�u������|�h�=�>��@3�Q4���F�|��W���($r�T�lc� 7(`������3C�`��GIs���Ǟ���ƓN�F��>���� c���.�m����4ž��T����*I�)0��ƃ���![����le#���1��x���El��j^���O��PK
    +Q�H�b�Y�    1  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/Prn.class        �      �T[OA��-,�"
D�m��w�"Zk!`AB���M�.vwa�ۢ�
�&�Ml4�����W�,$�"��=��̜�93���� n�!�?�34���3�i�8C;��2焽dن(Z�OcHh��V�.T��RH��
�r�R��eu:�����l!L�s��\����uj��ĳ,��(��)G���9�ZxiNԃ�:zY�,Ssm[�����55�y�$�C�\��SN�Xql�%��е78������Zgh�8�v��������w�
(hQЪ�����6'��3�2D�G&ln��c�򚣊�,|����G��Gb��n�ϊ+t�1ۃλ�ɋe�m���96�y�����{P��|>�ڥ�t�I�ߊ�I1D'F���Bݸ(�� ��=�+A��C m�hmiˤs5�</���vYK��<�u����%9-wUؤ5I@|�t��0�+�l*]][���j�
���b�jOjwa�Mfթ�Ld^ז'�O�9ۤT�c�ڐ=�B�?�ul����zg8�!�ƙ��Q�u��XMmү���	�ý�?���C8|Jr����i�*y-�ÉO�µo�*�|G��b�BC�DH�Gt�,$�z�:bun!�A�n��&:J�f�<+@e1����]�����ċdbh��ZGr7K�����=/���"-�fj��Yj��PK
    +Q�H�ms�'  �  1  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/aUX.class  �      '      �S�NA����� mԊ�(�8�=��`mIuh���.+)vw�^��/_ɤ����S�$ƳKH45�ɞ�s�w�s������ ��'�B�Ql1L<��]�9{E�`���5�����05u����bh��ıʝ�wՎ"4���W��x�R��Z'Fa3d�@s���|�c�&%]��2LY�}���X�#	%<� I�(!ʐ��g�0��0竫�
�W"��Ձ��������xs�!z�ZزM��	���a��]�b����j��Q$�CWb�A&��2��ƾ�0Y5t���=�������PD�%̮���mO0̏��N�r�T�aE^��}���r߷5�?46��n��^�X;��7���`���o4e/N�

'����(ѿ�HwNI �B���M���	Ԫ#�Aw�T����K� -@S���PnG�"]�z*�dE\ �MOC<���{�e�� ��˥��dO��L*�-�9� �e�|[D��]K>Us#�Mz�!Z�!�C\b~�kߑn�B�����E�_���Y���0"/��<O�ɇ?PK
    +Q�H�9_+a  z  1  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/aUx.class  z      a      �TmOA~����+�����p����O�@OLx����c%�=����_��#�?�e�=�_�~������>3��ˏ�߾����5Sc0�j�mU[��\����Ѥ�0�w|��8�<�pO;~[�#����$��G�<�MGx��&ѓU�B�d���U_�"Գ���j��n�I'dծ#�.97��
ݖ�2`0}u���c�W��3L���w�a�NG�L�ʉ�m�B.B�s���u�^�����V\��˾�)%�-�b"�E��>���GZp-�1��<q#�F��M�쒿C��}G�j��j�M-rAt�;���P3Z\�ڵ��x����=�y/G��������xwu�%_�lb��*��(3lX�w������M���]�*4���PM��T'����!sr�fML���)\51����TdwMea�nj	�h�)��@���&�ꠏ%[��4*5N3��;i�\i��'2�G!9|�F3@be	��������Q�S�˕�����A. 
��!�	8Czj��hT�1z��'�w��r��]�d��z�ܥ�.��hW�
�M���#�,��ĳ'ai�g� �H��_~�h�9iCR�/PK
    +Q�H���  �  1  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/auX.class  �      �      �T�R�@���J�r+Q��R�x-mA���۰B�$��-�&>3�:2��P�gC�2�LOv�s��~{�?�}0�����:C�n��[�?gh㚣�ƪ�>�־�&4�м#�Un	áZgD^h�؞��A��E����6�n��؉��Z�S�~	E�N`,g;��\&��Z碬�5M[X��p�K't�(M�ᚽk�2�(:ϛ;>���C�� �`YAJ���f~-
T��P�m���h��?0�<5���ֺ�놰�kRD�£�}'�n*i�H�*@I�?v��
�`<W�t�z2�E:��LE�4�Яұ��h���)���5�����?:pǏn��Dȏܒ��rۇainKsW�o�ܦ;k�#������ڏ\�ҿCW�(��(b�&l{C�4���/�d��x)S��un�R�5i$x	��.ȉ�i�Q��T,^<<L��ϔ>f���{fZK�����O��^�K�v��Kt�iʟՕpمЫ��C��D�1DIE�f�ރ��{��mϩx���t����d���Us҅|��kѤn��=ɾ܄ӈ����h� �~����E�<4 �	!�h��$,��/[��r8�u�`$���X���
��x|��)F�+��g�N6"e<����'{��l��[A��h�O��4� �Qa"���x1F��U�_�gK$�5��
�.0���Ǭ[@��D�]y)���PK
    +Q�H.�גy  �  1  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/aux.class  �      y      �R�.Q]�Ucjк�]"i�4rO�D�DZ�>5����̴ә�JB��ę�����g��ʾ���' k�Sу�8bH�1�i�
�
�	#zeee��
®�x��]�I��2m��&�2��K���S�a�1x��]�W����%�&�=�[2\��c���/�;�5�3�q��uE�*�ЇQB��;�5�}�N�uax����@Tn����O�f��p	�������߆������JX�wr�VK/�����Zu����~q�:���G{���|?wȸ)�N\�`�@��4��������s�~�D2���G$ץ�l����H_*g�@���Ȉ�/mꭂqL �פT ��0��_���.݂��~��tU�e�PK
    +Q�H�eN�  U  1  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/cON.class  U      �      �S�R�P]�-1(���Ƚ�@@QQ�p��f�V
�iz�ڤ$i��_��	�Kqd����q�	���<d���>�z~����$��,Cc|��5����1�5�8Yy���F�6��H�#a1$4���e~(�jM)��Ε=^���FQY��anj�CԷp�QM� �?2�C����,�d)�
��B�pV,^-t<����Z��1ϗ�+�;%���}�������b.�P-AH���%�j�%?K?ȌW~,����Y�47xQX����UԄ�(����D�pJ�*�t,*�׏\�U�r�4��w#�'4��2`2nxp2dt�h�Aܕq]2���=�{���>�%D�BB;�=��WB�;�M�U�5�U5�ᆓ�*�C�e�����;11���y��U^q��⡄G ��Uz�N�/e��{c̜ͲɮV��by��ԂZ;8He�l����r�g�kK�r5�z�\q����[\U_)��:]0�+�9&2�k�^m9���2$�z�j�_�My�f��G�bnZj�����cWO���`��V�4>��u�)�0AR�HCգ�4
i\H$�\x!�H�`���vn+w��:�s[u~�Tçh'm"VGs;�:����3�<�H�>+^��/4�vPP��x��&<&~PK
    +Q�H���9'  }  2  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/cOm1.class  }      '      �S�nQ]�@��hik�bk[�å��Ԅ 4��6�"�vN�Թ�� �O�|6�����Q�=��Mәd�>g�ך}f�� ��3���j1��V��0�\�t�%ۣ�3�s��m�P8Ƕc��m��f��k�S��*�:WO����H���^]���9BXD}l�=�xWx�U�eH����b��*N�"�>�Jx"᱄G�$����K֕���G�*����s���/�/O#N�5�!�e��dD1##��(�b'�y�H`;�dcX�u��nR�%�#��l����չ1����>hkܨsG�mC���E��q=��|��j�4�����������O��ը<8��X�y�~��a��-�V5{�(ፙ���L�7I��x�a��l��AA�l��>ڗR�_k`���רe�T$�Jf��)���&���Lb��A ��K	�ᎏB&0҄l�|!��l�����o��BG�{�n��Q[g��`1�/������j�S�Q͐ͥ�Xcu�[c$�:���'���f�3�ޅ�����譜�Jj2�9R�O>�PK
    +Q�HO:��)  �  2  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/cOm3.class  �      )      �S�NA�N)][
� ��P��X��jBjK�咀E�7]VR����E�J&5DM| ��'1�Y�H���&;�̙�}�33�~� �Ǆ�L���"OV�{F��K¨Խ�mm��1�C��	3�m
הg�h��%EǨ���=�r��ˎ4�23J�0u,��L���u$����k�����.e��ix�ᡆV5h�h�R��;"���
��l��$
���6,O\�+)���6��hJ.a�s����Ä�E1��(F��b"��b���15�$n�E�� m�����d����~
cU[�͚t��4vՠ�h�v['�CX��ۧ��ګ���}S�ۛ��N�����t��һ��z���ԕ"B1����-�I�2Wq��!,�7j���A���5��⾂^%,$��CXPL r3�9�`��TB�)�g �;j��DR��_�s�$����?��t���.nu1��ͯ�O�>��_'�������>r*�.��0D���41y��S��Z�,|��9R�	R��|�EX�^��/PK
    +Q�H� �  u  1  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/cOn.class  u            �S�n�@=�$�IM[Z ���[q�?��I*S�҆$oǍ\;�%)|
?�3R(| ��u#!Bؒw�v����|����;x���;�\'�d8�شM�)ۥ�3,p�7���:��葵�PН�����c��&W���+�Ĵ��n��NCwæԇ�9dH��NR��}��?��W���Q5�J`�Ix(၄��I���f(i�O]a��i��O|����rԄ\'^�EX��ߥ$d����Ĝ�V�8��I,��D��XD)�%\���q�Ω:=���؞�m�ɭ���U���9:���5y�2��"��Đ����2lkUu<i̓��m{����=����Ｏ}�e��n��Q_({��� �g�H��]��� ��]�q����h;�Q-)��ԩ2��y�b�B#D��D�V��4lQ-� �e��!��B��Y�zhV�B�-�Z3G{�0��kS\�"��r�+���ۭ����['��D�봮��i��蕑�50b�!?cyB,1�ӥB���_��+�&�M!L $�
e�����'PK
    +Q�Hϐ�=#  �  2  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/coM1.class  �      #      �SmOA~�Ζ��jE(��7X�o�Ʀ�-H���8I�wG�-��Lj����5���A"��z������3���~��������:a�q�jzO	�I���״�-�yk;�q��aN�M��������]�b}�ׄ���Ū#M�ʈ�#$�dW��״E��z-�u	��]����ᡆ�k��A�pIC����\$��?b.�+f�	�隢(d�Fװ<qƮ�좚��yDKr۞Ý�!���V֕Ʊ�
LBD�r	\�b
�Q�q�.�a�l[�'-�.[^�b@H�l]���i�F��QB9���'�v���R+���v��z��n��#{Sޫtv�>T�=w�Zy�;\+�����uňPN���`��)�cXB����Y[Φ�����JepW�^&䃐�J�h&�Y�_�)~*�X���Za4W��w�\1�;7y��U��R���>n�1����H���Yx�M?X�b�3B��ȡ��,g��0���6��"��CȞ�?a���|v?�	s�H�H���� �a~�[a�Q� PK
    +Q�H��ߤm  �  2  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/coM2.class  �      m      �T]S�F=dT��C �!m���8D@h��$��j������ʲ�ؖ�$;�?iAg�����t����s����\gh�i����{��{�v���~��L�@4����0�l5,�>�ɤW*2�f6����-�Ѫ�5�x��^�e��f{-�"	4/��C�r6��7k{���s]�A�}��+z�UT�޴&�yi4�dP|E��7]�v�ɛj��I�{�8�QU����̚���i��q˵j�k��T�!�*L�Pp��E�EDl�����!�q^�c�K4�z�t����)߫�&����0��5��Η�M�M0��t�j��kٍD�_�5^v�5�	"��� �����2��5A�+c��"��0�u	�8Lr��0�!�!�%\��>�p�C\�w� �!�ᆄ�����v��C(cz���,�\3790\���Qs[�}"��������Ҟ��,�z]���LI	��^���t�j�I�0�X�^�PB��#��j�!�k�5�I�탃LaK�<-Օ�};g<줼���RM�ɮ���TW�G�z+G:Vf�yf�agI4h~R�##��Գ������?y�����3G��oB�����@tJf���@�����`�}��؝�)ibiXX��A/�plhzLb����m}'�/ĭ�ݐV҂أE��r��H���뻡�F��&F�Ifc��G���7d�p�V���(͖�?c�K�9�N�<X�#��	��~������'�R���v��O��ݏ����^�8½���1fJ��sW�;�DX�.K���#�����rX�	]�=ƥ���v��r�|ǘ�����gO�=_���>�7�}��o���y���b�7\�w�1}�t�x�'/[pB-X�E�PK
    +Q�H�B)  �  1  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/coN.class  �      )      �S�NQ�N)]{�"��(�x�{R5�ڒ�ZL�b�w����ݥ{�oeRC���i|���DM�n�gf��f�9�����;�u<f��7�C�IW����KzÌP쮡�Q�w����vC�&NT��.��v��ƞo��	+uShj�2
�!s$�[nW?䕎e�T���e��T�{�G�#	%<�p_�$ႄ(CV_������WW.�3,�eO"��Ձ���L]������F����m�:!<�X1�yޥ(�p/�i�G1Ek1�q9�Yd�H�
C�j�SUC�l��-�s�{a���l(��fWtzꎷx�_�h�-�X5�*^�5�R��rkw�}��x��h*/ܚ����vl[����f�o������R�V�f9�<
A��[:�p;P���ݡ}PuGK�..2�(���`SCAr;2����U	%S��d�z� �E���A�<!�	٢K"�+�8ĵ!����v�=�ߦ��S,}�r{���p����0D�����X��!Gɟ6A6�Z�/}��)�d}U1���!���¸��PK
    +Q�Hw��  

  2  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/com1.class  

      �      �V�VU�6Ic�P-�b�a
VԂ���h�0lҁd&L&	Գ����%�@��t-��W�|������b���?���'���3 =���l�c��Q�V���a`�L���tX�Gg��[i%��6���+�������輻2�NWh��4���#1���)����8�f�$g��#m���[k\�n3\\��bXʤm�Nܱ���$MifR�l�<���8�N,�r�.�;M�LS[J���B"4��P�H-�ێ0�7���:\Q�1R�n�zζ��(�c�]t�i��I�?��P�bU�&\�&5��4}8K��cp
�ע�Sr��,e��)q�s���GV� PÆ���r��l'�e��M�U�U�D����$TI��𪄀�Z	u.J��� ᒄF�N������)����܊�6�f?C�zz�I�A}I�Hޥ�GүW_��[I$n�'3�/J�>خϫ�'xR*ԇ����r�o_<���M�`9�g�FU�J��k`W�%����r���?w���}��(a+��L�G��;O���ф�2<`2��A��x[��[2^pE@3ޑQ�>��]>�'�}��v5Z����!�  _���������o!��u����h/����~tY'>���M| `P����Z�Z���~�p�B�l�4���A]�,�J:�s�TK�Rs�m�J�)�J��r�Z�;-'+2V��<���e�H�Q�d�����#ϊe�n���չ�xa-�V�W��>\��fFG2Nv|$�YH���)��1r�`Y?8��˙e��(|F�>��dI9�1yA���=8����4PԺ#c=2V��H�[F������܁�c4�ϫM-�[���[�ɖ*#�r�r�b�
_�'��g`j�J�'�SÁ�L���B=�6�Qw�R#2�Ԋ  �R4ܕ��"��Q`�L���U�H��>:;H���S��hKԲ����Z�C���}\M�:v0���������T 1���G;��z���rF�T��	C���+b���u_Nw&b����)��k����]��ەGy��x�*��X�%�ߏ��5_���a�\�&w���'��SD;����G��X�"���;������i�Vr^�S�(��Ja���F#���-,vu�:�1�u��1���-z[b�E�4R3����)��I�
wWI��;/���PK
    +Q�HA�  5  2  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/com3.class  5      �      �T[S�P�����MQT@�6\B�;��RP0å����XMBӆ�������O>����"3�c��C�����M����@K�h,��0i9Vq��=�Ǡg����tm�`�\��4�g,C3]�ki+��ϰ9�zi��3�B�r��\��bz�;T0ˋTp�[�-2Z*ĜA���mn���Ե�;������_�rT�1}��NQ3��m�Z�r,�ל�&���?�_�Y�k�;$�󅌂��HX��KV��%aQ]�$�Q�9	������Oc�a�,�_�A�a=@k���"Cl�=�/%��鍥�)� �LA��6�(��WA+�"hǼ��:0'�������7����T�%���MW�э[������]�ȥ�{^=^v���r�aDO$��y=��R�Y�����hN�R�����n��0�zS��&絤k�Qka`���v�։�.������K��CN-$O�`XX���I�pU�&�u����8�8�z�����d�袳`���?v.���U�
�I��糮��^cx@��!D��W�)c�U�(C;�mra��8�4:>�S=��Fߣ����C����u�$���yE�#�����q��G*��P�SF�xL2ə��K L��!u���F�}ӫ=fhB��Z���#�X��5u�PK
    +Q�HִLn�  �  1  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/con.class  �      �      �T�R�@���%@�CA/�B1�]@���@A��ʿ%�%X��-�&>3�:2��P�gCQ�v�'{��~gw�����3Ԇ#�7&�p�����5
"���q6Ķ����9C3�]�2W��Ѳ��Y���p[�.E�:%�Bw�ά��/pͰ�35�Ynf��][p���C�)d�m;�Mmb^'���Y#�kY������l<c��Ҳ���]���1c�a�s\n�u���*XV�� �`QA@A�UA#CW8���EW�[��I�'"����E��r��C��Q�p�z������
	����"��{{�|ț&߮x:.zR�MT�]E�����SQ��*��Wф���X�oh�P ]������ BR��)�Iq_�0�/n���i�ģ��l���� ]6ІC��(bhMZ:Ϯsې[^�B/U����я&c�B.�\_K?���ܞ����չω�Y�M3s�E-��)�t	�a:\U�U�ә׫@�	@�)�*f�a��d�E�tV�^W���6'T�����k�*�uy[�M�VM���z�� �]�`������%�"9�<���y���������M��xi8�u��hz3ݺ��eh%<;A�#%�����7�%<���'}���p���e����1L�줶T�^�����S�	0j_�X��+�XK߆����WD�x��� ���
ȕB;`ު�R��oPK
    +Q�H@���  �  1  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/nUL.class  �            �R�NA=Ӳ���m
��-�1^x�1�k%�@�ۖI�u�K�[
<�>��H^� >��L�Q�za&�}3��s�|3����� ��H���a�L>�/~, ��s�5Xj�X�`���#���e��]��f,�b���J��m�ȵ���[���E[��ZV��=���vx }���u;�4�'�qR�E�F]��vc�d�Nӱ�#���1-Pp�޾K���6Yy��͚���y����'��k��.�� ��2��8��TX�`�Y��
7؈���0�b7��ߗ�����u��_����iQ�P����@��<�5�ju�N}w��U��Ý��A���yZ;���g��Ak�~a�Ά��(cN��D>��Y �O)>�/(1�y��`�U
yhy���Md�X�y�\9��G��2΍P�
0�i���PL�n��	��XI�Ø@��@���S���0f�K���� ��4�CbJ6W)��ϸ�=�a��U{#W5�x�53�R"f�Q�>�-��c֙�5�PK
    +Q�HL��}�  �  1  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/nUl.class  �      �      �S�n�@=�45&����r/�K��OEQH*��M���X�S_�IZ�*R
�>��B̺BP����3�ggΜ�������'x̐,����lώ����������G��kum��b,���Z>o+��k5�����a9>�}�r�~$�Ad�C.F���^�oɈa�/�v�y��X�A`{�~$�a3��d0�|=c���4p�4ljHiXԠi���n�G����[󏼆�(�i�,r�R�@̀��E\�a`C�%TtdPR��F����jy\aX��]�g���p�"�U��ӶS�h`�f�6�vkrx��a�#_L����� 
_7�Ǔ�Nm�4y�>E.����Z�m�*t��Aa��:V�Žy�W[�TRY�e���爖j��M�p��,�$ry�@�����1��tz�vU��$��(�X9��	־�֔ F4��$�2x��1��Ѱx�$bE�����9Q'��3�}�au��׿����Y���S�	[�a:�`�H��T�PK
    +Q�HR����  0  1  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/nuL.class  0      �      �T�R�P]�RBc�&�(* J.�
��8\�NH%�&4M�~���3�|��)Ef��������k���>I�����^0���Cݘe[�8��e�ڠe2��NN+�}��{Z��-C3�k)+͝)��q�Ҷ�gh���3�l��l���T0�=*�ŭ�M%b� ���67��r�Z�m���R������,շM�u��i���,S���%���k���'��2kws����Q2�	��p`��-	�$�K�$�K8'A�p^BC���i�2�E��<�>�W���������鿏�h��鍥�)� �LA��t)��[A3z"h�.`6�6����"�$#h��2&<�q	}2:pS�D�dt��F�I����Ȧ���r|�Ⴟ�]�iO�(�������r������΂9$����]�0?�|d�s���O�D�J�t��˰}�d�l0�AL%$OgX��|�G'�⪂1<��jƳ@���Pfh�q��}�U��
6�V������0\FMS����Z�?gM��(�����!D_�W�*b�U]/B;�]r�v#�h��v��7|�~��_������k�7Hd?T�(�xG�sL,���ˏT��1�B��j1A2�/��#L��u�U���}½��.
34�N���0��JV-uK��PK
    +Q�H�W�  �  1  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/nul.class  �            �RMo�@}��1M\b�����B�p�����)�P�rh�7;]E�����/��O�P$*T������Ԫh����y������	�1,��Qk���Px懾x��^�riy��r���m��CѠ�L�6xG�ݖ�}U"�g��s�]+~`���/H���S?�Z/C�#dj3��C������Et����x����(�lo�0���XSQR���b��G����z=b�3��"hƨ������OT�״1.]s4��4�Ӡ�:�
V�Y)b%L�4w��Zd���0n(7H��!긁�}���4��GJ���!�I >z��v���λ�����5�E[��i3��8j�x�U�0�n�o�0	�5����Y��iX*� ���LL����(]�I=@�Hq���Hy��#(�߰t�{_(bxHV��@A��4l��XO	��^����wO�x�����YJӰ� �#O��L��\&�Fg�H���*�Ќ+=�0ɽ�j�}�qK���X��xL�t)P"�G#�I�����X<kY�h�PK
    +Q�H��7�  5  1  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/pRN.class  5      �      �R�N"A=������U/���>m�ل �H��b|l���`F��M0�}���h|0��Cץ�Ω��~x���&	}��!�m;���@�O�6��gR�[^M^Y����U6eM�v5!y!�R��V�r|qj;7�Udݷ��x����f;�~h��aACD�F�5>�����eg�J1�@1�AQD1���(��Gb1���n��I~DE5\SVK�i�r�:Q�'�ꪓ5#�o7F�����&n��	
����B��w���^�@5�L���	������b6�)L�M����?�o2:�YE1DX�l��a��Wa��I��[�a � |a�'���r��u0z�I�_��7���q�c�Z}��|
�|a��;��/���b�o��+^��i��	PK
    +Q�H����  t  1  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/prn.class  t      �      �S�R�P�mI�A�PPE((��?�f��)���iz���$i��O���Mad����q�qp�.�e�=�gwϏ_߾��C 6�c���_�n��K����w��Hh�p�w��q��-��)��m��ꈴ��6C\��1��P�5�E��ۼ�U��͒��Ӌ�Z�l!L�h��=W��좰�|ߪ��}�4dN�e�D%V���v�;osC0��x���V8�/��	+��e�����×��f%$$�H�%\a��ϩW�l�6
m���K�-�$e���$�w��WԄ��������9]jŵ�n�șؤeT,���p��Bs��  �@�����[�U�(�WAn*�pKF�}���}�'#��2:��Àwet���Q��V�zך�L�妛��*�C�U��IF;hsڷ&&��Tژ$7���Vm!ᑌǾw�"g��-��s���qfOfr��X�a<�H�vwӹ�o'o���֒6祪م�T�u2�}���|�Vl���S���K�^lC�ټb��ɉյK�����fp)"I}���LIz�-�P�d(�=��!��z�!0< �	��B�G7Y&��A&X��#s�@��芯���P��kua���ct�u,��o��1~��1㣇 �����c諟�;))�i� �Oɇ�PK
    +Q�Hq�l�  J
    ExNativeAccessWebcam.class  J
      �      �U�WW�$��l�J�kX�VjE��E��HH[:$Lf`fB���R��ڽ�������x�.��c�����f��i9�����o�����w �R_� ���/^_�����;�o�/e�5]�O
�\�Wmm�u�b̲.���� �t���!���q#�,����#f$+�.0%5�����1�0l�bv��I�Pu&@"�ձ�Ϩ󪢦m��0����F�P��s[Us^u��ђL�4CP�B�&ȯe{�M���\��Y�ѭ�Ǟ��a���b�5"�t�l�+��#9at��𽦚dkɐ:�kI9�M��	'`%�����"I
��Y5vQ@���d�{ؤ�J؁�a�s��Tݨ�Z>�rڇ�8Y5mL6�L���K̕iv�W��#��M$�Q��"��"6��Q-�FD��:�Dԋh�Y�[4��C�k�)`�/��L���5�����U]�"+.ݵJ���(�7�Q�_VrJ8h��G�o(����hq��e���%��]v>_����w��P��N��),W�-����[��䬡S����H{�v/k^���N	<T�򮡝�K~�(� ������R���!�;q�s2�8HxP��8ʹ�8tr8.�>���'eT�a�8�]�`X�^tK؇s�cH��?6�,�A	-Jh土�HP�N�����=Nsx�C�CX���/��8��p��|��R�]��i@çam�S��."̂24mi�i[B
�*i��ԤC��cw���Y^L�$���4��kf���w�Ǧ|+�.���p�z�_�g�4��Q	� �i�P-�-�y\�*Wi�k��L�~__��XG�� 7^�K��iz؆+��*?��ktn��S������,�����%\�[��V�.��(d��w��=�y����g>��X���h�'���QM��n�U<T��)a7nR͋�

Lgi_�c�]�������`�b$������t05t�Rpֶ½������YEO� n���#|�>p���q�J���Ѿr|C�ln��E��;��*\V�i[]uU����J��V��AvSo���
���ԭ�����䐊d1��%ϡhW�X���R�W2x=��uO�[��)[�m�Z�����DF�=����1:�������+��.����p��{k�v¥��Í7@���z���@B�WK�o'y��D㍻�p-��⣟�I7eZ�ar����ϰ�`v;;�ے���k�d�)T`�������dwrP(r5�C;��p�(��"�D������EJ��rƢ�dad�̡�O⚒+\����gp1������6>v&��JQ�9���0�=���H��-��,�$Y%{*y0�iO�3x������6��#�����)Y\�`:��#��a_+������AJ$�X��;���i��1m�?PK
    +Q�H�~��  �	    _004_/SendCapture.class  �	      �      �U]SW~N�V�V(UAE�6,��ֶ
�*!�� - 1�-n�,fw�� `ۙ���U/:�L��2��^�W�'�Ծg7@�̞����y����׿���C����у�-4[ˏŬ.�S!�[Ѝ+b�GC�ъ�V|�k>���H�r7p3���rT�8�0.�/$d�'L�è�[qB���		��f��eM��:��tt�f��uK�,.�;�Uϝvm���ɖ,Cum��޲jjj�K��fr��#������{��Fr?��Ah}���U��Y��Uf5[׊>#�������9u���Vu=��2�'_�6xY�ԒesuV/sk����َpd��7m[[}-�޷�b����ʹ��[��NPE]��U�JTaJ'�����b(�Go���Pe�	_1(�W��7�lCse|EƔ�cZ32��KQ��5�R�U�B���]�S�VIB^F�$|#�[|'cNDw��IE�d��ny ��d�.T�	)c^h�v�J���"�Pf8�f�1�޿@Ѻ^v���\_Xti#��[չW�|fZUNM�'�qs�:���ш۾��w����嬏��B-:5�jL+����pĵF��yn�r���أow�v^)��S_A�rL�W�����IQz[w�M&�:��|!��sj�n.�]���H;Z�Xa�R2[�����m��PX�&�`�/~t��9ĈVǵ��ēW�������vo�Q�R��0���A6ǫr[�m��#���y�6�&��k�H�FQ��}�� ��^pV��s2�'��7S˵Zv��t�A�PkK���h=�͌?LW]gb,�Z_O�R5o�<0����Y�r��'+�	@ �.0I��+_�7:K��%��W-���Ч<C�O��8�G�J��/p���]�	�_v1<��I��5z�`����N�!������{�X.�D�>�S߲��ߌu��uNT���DXa���H�7�6����?<���st(��u}�(�c����t�>�M>(��=�ßUq�t�H[��!��<.4��
	Q����B�E�����눬!*��D,ORz�C�h�@|�ye��9K������r"�\��m�B�[2ۏS�j(�gU҆�Y���V�w��:e"����7??�O�u�3DϬ�����&��m��Z�X�a�� =������m�?M���B?	�{[u`~[|�����?��Du��F��8S�7�^��m���V��PK
    +Q�Hh��aj  5    _004_/WebCamCapture.class  5      j      �V�Sg���IN���r)� M���(��̐�@CZ]=MN�@rNMN�n�6+^��t8/(N��N�:&M�N�n����ǟ��@?��9I,i����y��}���=���>�>�ͅF��?f�#=.Hy�e���x���*����w!��,	�H�2z]��a&o`��y�For�æ��8sN�k��9�(�~�foa��L���]�2�\؁G��[��ęh2�e�����qJ�6tJW	#�;tJ��A},k3Ӛ�jشDڛ5�W��Y3���XkB�{����x�:ff�q�	=av
�zo��f����n#�	�CFLM���:�Ԏ3��F��n5��y��>d�G�2���Xo�+�V�#A](f���:���]LhC15F��T֖?�m��Gm��~��n��8j+����(��>��Q�x��m���Lƴ13a���~��Ʉ����+m(5�(R��{yV[n����
�H)�a(�ۨ������V��� �q�B�����I��Kr(�HƵ���܏�
ގw(x'P� )x���2�(x�[E�
g�>���
>�*x�
�^K�{L��Щ��\�5ejN8�U�	c��M�`�$������9�M���w ���m�exthD3�j�\�%ԗ����-�1Xꛗ�"��#j�4���<�Y�;�F����2��5k,�>��@��o0me�o���O�H�lR#�ǵ��3��&���+)��=��e����C#8	�o�D�t�iEgo|�	TM����НP�mt�؇��̨@�/V�ìh��wN�,��=>dIM�o�D7������(�
�g)�4X��������?x���*C�T����LM���M��&��xq܋chL�wD�G\x�	,"����i5Fh���ܢ�'��4ݤ��c�8���B��M��O�B���a�]�4>��Yܛ�}T3G�x��ga��sT愞�8K�7x{��t)���l��L"d'��#樂�1�_&VlTMw�i�zԭ�\`�W��ށ��>�.�Μg	A=�a�L�k]����?Ϲ����3�4�n����s��3+ �����=f�|!J��% ۆb�=C���ѵ	�ѯ�H�C� h��0=�6W�M��<�}���I���W��أ`J�sKK�׉��'i�B��ќ޵��]�����훽��>�'~E���ݹJ��;��inlk!�?�^��Wt8�'�d`��޺ƶ�]N�ۨB��3)U�9�Zp@��9Z+8^ҰWWr�x-���J8i}zg��x":���pN�7�Ó���`Oو|)��h_���c�1�NJSv�ۧ|$��`��'��@{�Y�4K��hG�}��1�.�G�՞d�k5�MD��Ξ�=��{d_m��4�T,��Dr������K�������@3Q�V��p��5����,���D��C�Kp�(�!����NUF�W�%fG���)l�{��Z���E�c.��"����#����ƶq-�:qW�jy^OV�A��@g>�EB��Z�,V�ϣ�Z=���e\�ݑsX����e̐ƚ�Fܿ$�<<����ֻM�6�p��[�P����59l䃾�%�r��a�r�L�W�����5�.�*��h�vG�25��ϖ��sxWFn��c���JC
6R��ub{�}w�`'wc�Z��3��¹����O/<f��e�
�����K�]�w*h��?��c7��
����%�KV��b��9��+�mD���l�6��h��}�`
V�{�&��8M�;H �HM�J�[;��Q{DGH���呣��3pp��R�ITJ���ָ��^��b�a�lv�7Ϫ_�nj��A�lK�Enl��*ͮ�v�h�+��PK
    +Q�H=�;/Q  K    a.class  K      Q      �Ti[W~G �ID�&�b������kj�FS�m]�n��c`�A�.�{�s��}��?�Oϝ�ȇ���眙s�r����� ��o
���ج\B�Yoe��R0�.�S�M�t(P8��|^A�i��a�]a	G��]��E^zeG���*�9^��9�vv��nҶ��]��P��۔l���O�N^8ߵ+���/}��ꐜ6��*�������)P\-�-pkSO�r��z��Cv>�%rmÚ^��D>����48�&�b֞�k����ˤ����2)ON��Q2�XOK�xJ}��)�.�M�'yZ<啂�,�e1_��#���<g��["$.8�p�_4���]2݂L?�+f��c�gx��-�7*�i�3��>�(C?�Y��A�s��F����Pp.f�,фl��G4~�s���%�׎h�u�~��<����W�Eסz�`~�Wlt��oyT\���wxl+�vy&sn;���v;x��dЪ�_A�`4v4aŒm�!'F:�
����7j��0d�7:6����on�lsz��SP4�&�"��6 !��
Bz���!�)��4\�Ѝ�5��w$����$Lh���.�}a<Р��x(aR�5����e70�b�*nbI�-��ቄE#H��\\B*ƥ4��T�Rґ�0-ᑄ%�T�FZ�KqV�c	K�'���c�JL#sp�Ѝu�S���M��4�;b2���1TT��kj��I׆a�xa�;&�]�@���I�DU�W�a�L�lo+ˋ�g����e�s��Te��^���fR���G�'��l���d��
����+X/8ta���Po��L�Qv�����A��������+�X �O4��i:��tEY���a�B�J����H7��� � �=M�g�M贊�&�d�%���L�6w��L0�F�H؃�Zخ�nb$A꾮}�����Ql��߿@�yl��Rbl���Db��M\�D$��x�d��g�?K]k�*���l��I��&Q�g�xf#�k|=D/�c�<�x�č8=�r٪㩧�rum���1R��q��h`����$����JW�ve���tɩ�/%�&NJ@h���+B�'��PK
    +Q�H���  r  -  com/smaxe/bridj/linux/lib/VideoForLinux.class  r            �T�RA=Kra��K�*",H��$1
I_7ɘ*٥6��^xA�0僯V�Q�=�� 	%��93��ݧ{v��ߟ� <�G�WbT������mn-!6-!��X.|�l�܎�-V](:��t8[0KL�x�,FJE��E2��F(�|@��l�3�M+),�,�0�?e�@)��N��Z��6�gI��t��1����ir�f�q3+ºv�}=RЍ|d� ��lnP�ndvY�Һ�E}��ˆ\��=F'�M+_��@�� T�\��Y����9�4��q�^L�7�T�bzNA��e�,:i�����+���M��2y=�-n�JN�N�m^�x��ŀ�^�R0K�%�
vZ�����騸��d�����zkl2N���n��D�����i2*�!*v��磊����ˁg�8d5�a��m�6��^�O�)�u8�]��uz��S��n�F�k�����)ſ0�g�Fs�?ZgQ�v�"�KU��,PE�*:�V�G�]ݘQя'*�x�����/��*��cx ����WLീEo,0��  .ୀw��-�9zm��ʆ͋l��x���ôu�a(����yC��#Yc�PH%)&ޡ]�]�<���I�{& y���w�=,�@���*G���[�¬�1����OiOS��ۈJ�r+�%w�gYp1�}���o�g��~<�j��M�6YAj�����n��7�##p�d�w��͝�A�t+q⍝!�#q���ϻ�E4د|G���`S�A�)�����r{�P�r�ۄ-���+A�PK
    +Q�H��\�+  �  )  com/smaxe/bridj/mac/core/ns/NSArray.class  �      +      }��j1���o�u�j��ejC�A\U��
��$�I �>VWB}�>T���Ei ��|��$�����=.	�vg����SZ�>�&6I�&b#��U�U��8����N����Z�F����<_����Yk��d��r��Hh��]����pl���l�:��(�e�:z�~:�/k >ҙU�GΗ��2N}9#�f!9��7W���T�_�@k�SF���}6V$����S��­������?��9�j��Z�nQ{��l�Κc-uﶨ�x�g'�?��/<g�p�����SE�5�~ PK
    +Q�H*}b�$    3  com/smaxe/bridj/mac/core/ns/NSAutoreleasePool.class        $      �QMK�@}ӴMZc����@�熂
�h��U�d)[�,lR�oy�x����٤�βo>ޛa���z� p�.���	��d,�1��P��d�o�e���A�J/N����&�x%�DL�Z���?̗"L	�H2&c��D�+�����-Z,d�
m�h�d�!�{�ɯp�d������)���{0θ�}��ɿ��G.,����*�4pT��/x�"A���"ҍ8�ፕ@���	g�,��`���L`�
�b_`_�h��)��T��CV�y����Qg?�ȭ��NލoPK
    +Q�HicK�  �  (  com/smaxe/bridj/mac/core/ns/NSData.class  �            }P�J�@�M���Vm�E����ϖ�ԓ�o�%niv!ق~���?��ߦ<v��f��v��?>\c�ЈF���Die�~�fe�p�����x�<)�r�s�����?,������L-_K�ٗ~��a07E�Z���������d�����i]2��4�j�=g5�����t�h���Csf��b�mU.cU�d-o�6VXe4�Hk�2-즐8���i��y��T���?ޢ�^��%����q0�ڢ��t=0Z������j؉����PK
    +Q�HSہ  �  .  com/smaxe/bridj/mac/core/ns/NSDictionary.class  �            ���J�@��IҤ���h�.i\�	/+)*ܧ�!L1	L"�c����|(q&)�"�g�s��?�9�o� �pH�{�{�~Dx������G�<���+��u�'4��`AQ7�+Nk^�x&8�[z�Z3Z8鯞a)���B�k�	�2^�LX0,�,XSo��ޕ��<$�y�j���q�λ�E���ơ�E_9F�M�`L`\�)#��<+��Q0Ö\�����j�d@��`�(<����������~��հKl�p�����7���Z3^1m��PK
    +Q�H��@�     )  com/smaxe/bridj/mac/core/ns/NSError.class        �       }��
�@�g5&�_�,E��am�;QA���NH���U���Ļh).��.߰�|� fh��Ɂ`�"ق0e��Ip��DtbI�P*��3��WJIE�Om�'f�,Bo��*�wR�Ws����B�J #N6\#5���'�{�AvQT42��E�z�P�r�oE�`G��]�%�7����Vq�
�PK
    +Q�H�U`�  �  )  com/smaxe/bridj/mac/core/ns/NSEvent.class  �      �      }P]K#1=�~��~ow���V$��EPY��łPSgȤ���I�����LeWa0C��=��s�y~y|��_���%C�DJ+w�P�6E�F�Q�b쉱�o�vI_��J�Q_$�;�;7�粽+��H�=����<�ŭ�U��"������f�����c��i��MpD�b�H%NZ�ҍ�&��r�
�����Bk>pv���5�8�C��I���;r`�&���s�^� �:gy]9��fF�p�ji(�UGiX����&�t���v*��*Q~$�6N8et°��+bI�D��i�&Vb34 ]E�t<}ߩ��N@�{��L��-x=G٣\�n��۔_��a���j���z?(�Pw�v=A	?	�yT}������ma��hO]�
PK
    +Q�H�:X=  P  )  com/smaxe/bridj/mac/core/ns/NSImage.class  P      =      �R�N1=�)���4j��h�!!$Q	������ִE�-W$.� ?�xg`������{Ͻm�����
5�t�b�H%]��ֿ������fh���b:�c8����X�֣TζNqyK�}#�sy�\Y~?N8�~�z��I��.D�<r��6�M�����Ҵi�܍o�P�0´�շ �f7�zۊ�vt1x�~H��~���醬�X�JE���L_O��ꣅr2i���R�yNje
c9S�[��PY��`1�C�*�d�+T^��.��p�l�l�y�Bu���Pf�G�K�:���UI��PK
    +Q�H�_��  5  5  com/smaxe/bridj/mac/core/ns/NSMutableDictionary.class  5      �      �P�n1=��HJK�gW@V�	Bj�M�$EEJ�fp�cWS5��U�,������D�J���:������' G8d��W�V4RZ�6C�5ꑉy������y,"+�N�e����2Z�[��֋�����Q�ϒk徝��"R��ucS�d�H���8i��t_zC9��Y||c�gy{̐�!Fc"""d�:�K'��gOjsU�F�+G�c<V��5���Q�F���������l�ا�l������6	h,�D_�i��22`e�ɠRB/�����W�Sӗ�ԯc�T,�T�H�{��^c���9�VĒ<k*v�@7��X�~���xڻ�m�U��x}�6x�� �������f��	�Ŋ���`�oc�|��։�����b��
atV����L�&+�����PK
    +Q�HR��  �  *  com/smaxe/bridj/mac/core/ns/NSNumber.class  �            ���N�@��
-���U�&.Z� �!,tU�T�&�:�idH��Z�j\� >�qݐ�̹����9�_� �pF�O��0}f�U��˴��2�_�����y��i!��K�Zn�?ewɆ���k�#���\��Bd��k�o��XYQa��б`�'���Wy_0.�-�j��zQ͢�i��?�Q�@q�UN�k��@���	��bM	z+���
��$Wf��nyƲ���v8z�
��j<�Q���f;7�T^���T7u_�F�;@c�N�.|PK
    +Q�H���;  �  *  com/smaxe/bridj/mac/core/ns/NSObject.class  �      ;      mPMK1}���v��j?�$���<���i�b���6�,�	dwK�Y^,x����d��`of������O ��"(���XH�Nj�*�K�
%	
,!�	TL��m8��X�4f��T&t6�C�m�W��i_����JȔk���M�a@�v�ӗ�,ʸ������A��70)�'|���Ȍ�{��G�G��x8ɹ۾�5��+:�X��l\@lh�(�Y����qfC��4UKn&�d21_�D��R����s��,�4�5l�=�5A�ܚy��[��r����h*�޵P���_�enuj�=S�M>1�&(� PK
    +Q�H,5-4�  ,  6  com/smaxe/bridj/mac/core/ns/NSRunningApplication.class  ,      �      �R�N�@=BnM��K/ !�gL$�)"�}6뭙(^��!��'�>�|b�	P�@%V�9�=3gF3���{�V�����(��G�lK��?Ve{i\*��P���@z21�өw�9<�*i��v�ךt�}~�#XJ�@������҅�Rz�LL:�*��%2�ѕ
���Zb����=�5*��*#�f^��E���$R�i;T��or���>�P1^D������g�4Kn
�5گ#��F~��q��*��ۃk�A�6[\sod3��9�Ll�=�t�a)ί"�\Ug򘩠�g�*��"ov7	y_�E�ʾQXA�yw�.��7�&�x���� G�p���s������e�9̊2&0������I1��X��G~���?�<���%�=�S������ PK
    +Q�H����  �  *  com/smaxe/bridj/mac/core/ns/NSString.class  �      �      �Q�NA=��ºZ�bQ)--�I;�	�ILL�6�>.�f���Կj�@�>��Q���	��p��s�={��퟿ >���Ê[=���t3P�i1�6�}�;�w���P���F���:��Hx���*�'����̓��n�E�O�H2d}i�la �
���{�BG���)�P*�\2�B�Ϭ?��2R3��ԲwsE#2&�OH]��u����Uk�J��[n��
��i��<�J��/��o�l���Gw�w6j�H�q���v�8Ha�A+�(8�bׁ��,�(��᥍M�l<�+[x͐l�}Z�s����"�o���ZS˾��2�s�<I�� ���-G�S�_x�c�g�D���.�	���^�d�� ب���'ʛ�7*c��G��ڄy�Z=��PK
    +Q�H]QToo  �  -  com/smaxe/bridj/mac/core/ns/NSWorkspace.class  �      o      �Q�N1=�� �KP|,LL\L\3!�;c�H��ah�8Ӓ�`��\a\�~���Ȃ��M���{n{����	���z�ǰa9��"h3���q�(��=���}-#ӳ�Q���7o���w���iJ?�c��y����W�V����z"����x�
���>�����%���Nx�4�i�j���?r�.w�bJ�*��z���^��W��9�V V�=ìUd����w��_[m�y����É"�8X�P�Q� ��PT3�D�!q�4���D��=ዾ�;R��w�FW�L4�rT�$X�L{���̢hs���YB��%�1ҩ���~@'�"3` OV䗱O:K�[t2>FN	l�P"/��[@��E��PK
    +Q�H^�9_  �  5  com/smaxe/bridj/mac/core/qt/QTCaptureConnection.class  �            }�MK�@��I�������G�C��\"��A�{��e٭��[�
��(q7�$�]ffg�w��ϯ� �x�HdB
��*U��._9�k�X���X�4g�a7����W����=v�P�k�y���r�$!zR�.�%o*-֮��#œ��˟AwJH�uJ8�;�nٓ�%yˮ��e��׽��Z��#x ��!9�G�j�	�L,e龈S��\���6���O6�k�����8H�78��Ț�!�ر�m�|PK
    +Q�H9�#��  �  B  com/smaxe/bridj/mac/core/qt/QTCaptureDecompressedVideoOutput.class  �      �      �R�N�@=BLBZ呴�%�E�k�H�RP
T�l����l��[�,VT]�|T�;6�EPa$��;��s�x|�����Xg�ho�y������[��P��t*��K�gFE�Ȁ�ṯU��Gr(�'�#�2x���4�g�=�r�Íx�J�Ը_����dZ���-�T����$�a�|R�mu3"gQ�;��F�<�s���w��G7R�wy&����D�1Zg�:��b$SjgXO������T�P��`X����~D������Yko��(i����c��-5�^��s�qb�����ޡ/#U���V�{���t�p0Qǌ5,bņw5,�-]ݎ���Q̭ZX ޮi0�Mq��9BF8ٹ�������rz��DX�l^b��?�SB�UQ�2U�F?��%�#,�|���|����;FS�������V��9�b��U��?PK
    +Q�Hf�ےp     1  com/smaxe/bridj/mac/core/qt/QTCaptureDevice.class         p      �T�RA큄p�r��Q��_�T�CAH�������.3�h|�|����,{�V\,�*�j��Lw��9;�߾�
 ���A~�Ҷ{����*��bw�ޮ�BC��-,�A��M�^8u�ޡ���J8R;�խ��p)}�ܴ#�l��yh"%��]"���>�|S�ad:�o���Z+��1�=[2Fa=2B3��z���"Q)��~���8��04H��p���i����L��끔�%�1�E]��Z��J20B���G��6$�P�`�\���Q�>om�&q��vt4P��&kd_��J4P�h�v�>�~$2���`��l�Vr)��+�Z+��؛ %���t>a�~�� ��\B�XXm���b�
�>+%�xke�Z�Hy]+���r<�G���l���$꺓�Ŀ7�T��wG�w�����R���u���ERЗ�ikR079X�fif�@g=����v"i�)�Pc�%Iw�wo�P�[V��Tk�q`����E�|�p�>�lx�lx�|����	<�ė��y6Cp��;8Ox��
�z�.��X�!���&?˻G8�K�+p���������ȏw�D�_��,��c���c�yR���O��!����? PK
    +Q�Hb�:��  T  6  com/smaxe/bridj/mac/core/qt/QTCaptureDeviceInput.class  T      �      �Q�R�@�/A|����x����R��|Pz��E6�,�~�_�	˃�GYΆ�r�rS��L�twv?>���c�!Q�^1L5쾐B5ҍh�:�
Űg{���#7��pnMײM��y���Αu�>o�a�cy7��ڟF���2�_�k�nZQ}V/�y~/">�xB�}���>�~���A*�t9���o�%��]���$X��ag���@�R%����4j�kő5�^�IڕX�X��qn&����'�X�:$P�a�:�s��
C��s�����˯D �}~ ��,%<0d/EOZ�;��Y��`���������6h� #����C��!�F��YS(R�(/1�LH7ʗ(ώ��m���c���X�VݤHKC>@�PK
    +Q�H6�\��   $  0  com/smaxe/bridj/mac/core/qt/QTCaptureInput.class  $      �       ;�o�>C~Ff�0F6�̼�;F���\���ĊT���̔,���d����T��b}�`�����F-��
K�C�JJ�R=�
JK���X�4|�ҡ��3�JR��AvKb��Ѳ��0010�v.VN����✟����������A��(@�`����	�Y�Z��7���ف$-���4���v�<� PK
    +Q�HV�@5�   %  1  com/smaxe/bridj/mac/core/qt/QTCaptureOutput.class  %      �       u��
�@E��H|���`��X�[�A�>�EVHV��[V���G���R���2���? Q'd{���X�	�ʈ�����V�݁EA�B�8��l�/�j����j=�:Q|��c�]d]���L��׿�"�\�lx�{�*Ȁ��%�Q�R"�r�	E_����� [Ɵ6�j�F�y��55X욶�if�L��P��Z�� �PK
    +Q�HC$���    2  com/smaxe/bridj/mac/core/qt/QTCaptureSession.class        �      �S�n1=N�\�Z�B�$ �xm�HP�PTQhP_�fcE��v�����ᩈ>��B�w�%B�T��<��ό��|��	:K��~"�*�p"��=�Rw���ᾜƖae���Z+��P����&�F���[��|�?�b8�� �C��/���8�N>�c�;�~�Lm�y�#��K�9��r�P���[b��hv��D[�0�k���:�$�Ԛ�������ƪif-����Q-�V�������`�}>���aXo�����t;�o�r�]��9�n�������T�$ϝf��a�e89��h�n���ΫE^y�%?�	� �3��=���KX}:���;-E<\t��f���Ľ6p�~ɮrj8jl+"~,�L�S)�,���O�#8���:�u��I>$k�4#��9���$�����k��K�G�����4�ƪ�p��S�&���[�J��h�.�B�A��w~�P�3Az�̑���X�o���X�^K�U��%�@:�_� 募PK
    +Q�H?��~  P  5  com/smaxe/bridj/mac/core/qt/QTFormatDescription.class  P      ~      �RKO�@�E��/��"^L< � 	MH���񾔕,v���&��D����2ζ�R<ؤ��o���L��?>�N	�Uk�(>�hr���sW
+��Y}�#KP�r�b�Xw�}�\M�ZY6�֣s+����W���'Py^ε�V�j�Ǫ33'<����sd�Oɓ.��Ģ
AՔ@N��s�I���fS1�؂C�3�&pX���Ώ� ���j�5!m�,���	B�ފ�F�W����ܡ�6Zx�����k�3�<���a�f�a��M�������S��k�2���-(�pD`�Zpc9�}�C���Q2O���x���H���GF.`���S����c��o
�p����#�+�,������������PK
    +Q�Hb�� I  M  0  com/smaxe/bridj/mac/core/qt/QTSampleBuffer.class  M      I      }Q�N1���(�� M<�zh<CHPC�!�b�w��%�-vK���ă�Gg����&�ɛ7�uھ���)��ͫU1ȶ�V�à�?;����PD�P���8O��V�g<��\��zx��d�x�=:~{��;[L&�2(M�����q`��)�TB������9�� �\��闯К�m1�6������T�'��^�Z#AAop�@����D������a��*@R�[���2��s3�8��B;ɑ��ʮ��	��j��[X	G@2Z`䇱����Q�[B�e�@t�.cNa�z'K�_��S��p(`�� �}�{�7W�5�c�&�'PK
    +Q�H
5;�  �  K  com/smaxe/bridj/mac/delegate/QTCaptureDecompressedVideoOutputDelegate.class  �      �      �T�N1�$!<ʫ<�]�.Ұ��&QI`%U�����!c�[�"��+>���*$fd���ܣ�3Ws��� v�����.�\����\�H�q��H�{��x�k)t���P1+�\��0?b#��PUzJ�M)��KQ!��K"��$�͕>}v��Q�P��ԕ
��Q��*��4��C�3����fRJ/P���e$��D�6�0�<�	�R�ǂ���c����J`��<�\hTUki1���1V(�/�sǵ4����Fjz��z���Z�S-?�+���)<���%0.a�(��އ���?�R��b��y(���>�mJ�tk�4����!w��/��̦���:�/�U��`��b�̻ev�qdN�#ظ�	�4��L�1k��3��	n������1�X6Q�_�m�.�l;�B��	+O��?	Y�GPK
    +Q�H1�捥  �  ,  com/smaxe/bridj/mac/lib/CoreFoundation.class  �      �      �X�C��b�a06v��!��4M�Ђ@���lS��JĂ���V�J��H�����L���I���&�Ӧ���L�7��i�6��f���yoޛcG<�吏p���		��c	!煼$�5<ϛ��tN�5kJB����ŧMS-�Ŭ�Q�-	�Uͅr�%f%VU��\�M[	=îJ��g#�T�5	]�(�gY1mjK3t	�l��o�E��gUK��L��^�|����U�Z�)[��h�Vg ���%�)9�$ӳֺ?��y@�,��R5�x��CA'���Z��5j�H�t��� ubm�dE��ɱ��}%5'�;'�t.g�U�0En�Xf|RN�.�rC���w��uQ�u�
�˱���rL�a��O1� X{4�E�O�̸�U%��:�;c�eF+]�~��Y�)��["����l��:��y%힨e�R,a(N�fT{�H��G.��R�`�ˌ��\fk�#Mo|D�~ծaig�8i�P�j���[�F>Z̫WY4ej��h^MGsZ*3L�ۗ�w�3E
F���]%�uR�Mc��ϔ�лɰ�e��p��zE�jFt�0��<ф6��٨��8�ڠ%ݣr��U͔�\��{���(F�&bwoͲ5��#����|�����vz%����3$V�'�2�:5u�5�l�U�ڱ:�"�J���H0��Q,����s�x!~�v	��3sMɹ�Νm0��ن�Ν�����k�aA�jz��*��l�9U�af�]9C�.�fɠ-�Ww�Q��`������U9*r�ɲZQ�e�;���2ۮ�g�u+�Z���}�	���D�s��a��up��E/\�b�D�_/dDe�D��2^*�/�1.�Id\�2&N�ݢ�j±e��<����Z��h�����'��I�l���=�U���c��#�c����9N��#'��%�����m`P�@�a�aJ��p�����t����3���áh|5'\����)��8����� �dd*�:��\zՍ�N=򑰝K��T�:5Y��@~��;�`�nlb�Л�]�&�3A%K��̢N�8�,x�����v�ŰS�D��9� �|���v��{��V�ى~v�b�=��Q'��6��/��O�n�Q��[�@��>�d��m<�����|���a{!�l�.$���SXG=�4dPy�S��N$����M�o[<j�	5���FAө�4����V����	�̣E��g��Ѫ`��Wr!�M�m��`����RpW�BY�I��)oTp#ު��ŭ�V���(�	R0��*�_��7:��GC����:Oq���CXõ��n�x,�a��6����\TB���!��-.�����x���s�t<��'�������h���+b���^Ҋ���u�kz��k[RM5Ϩ�{H�+ZVW��ɨr�f�`S��S��Zp�p/�Ӈ_E��>�j>|/�}x��]>�Z¯����������	�|��g}�u��|X%��a�/�%m�#�G�Dm[�:~yM<�:q+>�o"j�#�9)����ه���&U�m�~����o+��F�E����2��K�D��9���G ���+����S�du�˧v������xz���W��fx����;��d�����!�};�G�1��PlYzݻ0x��V�c��w�(��N���l���@��?-DNR�OB?�:��p$����[I�~�u{�Mtڞ!W2�'L�Ôo!u�o"�σ�n%�B�)��W�{Ƀ=�����-�2��om7��Ѿ,h]�1�{�E���+�k����J�>���M�4�xKݴ����A�5� �3��!|��y�9�0�:�7·�t�x�>��������H��ݟ���U�3�ه�/�#�|B���m��Cdɛ�>%�#��ho���R���'E�"�C�/v���~i����������5'�煭E�1�wҸ�PK
    +Q�Ha���  R  &  com/smaxe/bridj/win/lib/Avicap32.class  R      �      uR]kA=c�n�m�6M�6ժi�cC�nA*�@�f7�0a3f'��|R|����;�؈nf�ν��{�|�����x*��:�(w�XieO�:s���~ �Q��H�_l���9�C��'S�:oȞ��9�42jlU��Q2�ӑ�L~hT�O��c�gתC�I?�z��Y������l�
�,2Rk?HtFz�botسW1�	Tj��2O�C�C�C��M5���B#�0����v�I3�\
��2����B#�U����u��>Q�7~R�;�$p\D�O�*�+z�*�s�;���4[��\�r+5܂�b��Ğ�j���	jZ�	b���
4��T�
c:�:��]c��h�~?W~�8�:K��
���<�h3��R�+��8\T����<��p�q���O�L�E���W3���>��3�v�v�a��C��=<bR�û��'��PK
    +Q�H��>��  �  -  com/smaxe/bridj/win/lib/MediaFoundation.class  �      �      �Uko�D��+n)��n˾����q��ew���M�*i����\%�p����ć�@��w�]�D�/瞙{ν����_�� %�5a���LX4�c>1�Sn�pۀ���#V]���Qb1? ��I�sQK�w�,��< �I�Ȁ�(*s�m�~�<aK�y���ĵ%V��F�2�f�P��XMx!a�ǵB:%d�/n;A
%�<�����lL��K�8*iX�#j{((+��O�C�O�D�E,�Y��2�p6s��I�t�Ҁ��Ye�E�+�]�~ ��$$u��(/���r����q��'Ԧ�g/E���yM�<�I�7�[I=��I.�^�����rӀ�5)�a�'�ik��c��lrq��;�3Ѥ�Jtx ��^��z�ܥ5<��d5�+�yp���g4��K��ߢ�Q�3��d�@��Տxq}��a�P����w�]��j��ft(��7��kע�j�5��ݷ�6�;�Z�n�ߍJ�'y�>+^�Y����;��a֎i/3��Y|;qvZ�;9KZ��?p�����q�Y/;O�KˣI����]���y�b��(�/
� O
� ��w�W~V���l�R�T�O&&/{�d�_�jz����1���sU5!���իsh�4;�Rߕ�����4$����6*�c��س����1��NH�W�������^����g���"W�V��S|n5�"�k��W��`E�g
(x��&�+(���*��
���l)�^�5�f6?{3���[�Xɲ$g���W�����=J��I'�Y�軎��Fz�Ńa�.��8����O��qTd�jF���(.���(>�:΀���������a�$`��]�q���)pp}�uG������y|����
TsSs����474�����s�3ͧ4���j.�h��-�cl�X��i���"	xߢh�����PK
    +Q�H��хN    5  com/smaxe/bridj/win/lib/MediaFoundationPlatform.class        N      �T�NA���,��BA��uQ�H��&�V5%��L�C��%��TE_�n��x��PƳKM�	��sf�w��|{v����S�����¤�)9�X�T�d+���ZhJnH%�&�M�Q�h���2F�v`�ϐnT��q��bH��pm����z�۬m�g��Ʃp�eX�x=�����nk��}�lW��p$�z�r������r�����O�
��ii��!?��U��n��a��>h���.9&{�G��!��� �k�o���]�ԱP�=,�����$;�EW�Fh���G]☻��0ma��M��f��h�݀��D��P���ő�y�2{��.ۚ�K�a���Ў'uP�&f�X�Wq��K���_g�2S���ʛtS�RHf0���XN#��4�QJc�4��!j'�W�T�V�&C����QI���U��/�o)�h:K5eWqh:��x�]�2O_�u�I��n�t�*��M�)Ҍtb�Gx�P�5�_�R.v�'{9v�G_aſ!+� ����PN��N#�x�۔<v���5B�G��yF�;T�Yo��AGiѡ������/ Q���*�PK
    +Q�HdU=�  �  6  com/smaxe/bridj/win/lib/MediaFoundationReadWrite.class  �      �      �Q[k�0��&�r��nٺdwڇ�/ڞ!PH؈!{�m5(����Y{�a?`?���	t&�����s��7�Ox�ppv>gh�Vn�p2�V
'��HΤ��[�Ne��d��"I>F&�Y*n$���|�4OT�K���:N]}�ʑ�p)V�'B/��p)#��N�hh��
^�إ	��o�J�"���>�4p�����Hr���ᡇ&Cwr��g9�S9`�O���~/��D��$Za7�����_�7���v���%���'k]F��J�P���G4��`-t���曘��s���~"�Lf�ݫ�*Sa"�hm\�j⚁Zh�r[l��/|@�ҊC��ESwTV@��'�<k� ]_���t�T�#�)���E�'8,
I)5�HԢ�1����PK
    +Q�H�ا}�  .  $  com/smaxe/bridj/win/lib/User32.class  .      �      ���w����d�%Qv�ĩc+��PN[�q�V݀�HX�a -�`!r-��  u�Gz%=��Mz����J���}�w���@���������,Ap��z�����fgggwgw�'��� p�,������)e^�HͶe[�I	�.���n�ٶ_t��m	&su��SU���`�����^StA\��39˻h����<s�I�/ow6r̻�;��r�<�GʐⅬZm�l�,A�z	-�;F7V�<�LTTʺ!���{���1�F�BNN6��C���ƞ(0?�6=Ou�5rHh1��Xӗ`9�fI*Š%؏�E�ek�ӱ[=�$j��c+�9�KKlG�M�Ѽ��y�w<�m���ZM�k��CCN�����~�]��gwJ	�t����Q
88��%YUq�>�NV�l5y�7��^u���6�S�rCV�E\�ճ��-�W�_�"��	��2v!��d�����!:ݱ��Y��.3[Bײ�^1����1Z�I��ȞѳZ>_h�GI��X�h�|I)+%�,��8��J.O��FI>�9�Vq$L]��]�b��I�r�E��u2P���U�U���rE��2z��2��l��m���P��P���ǌ�|��[�,�=}P�]�Z��a.T������GC\�>���5�f�C�w�����fCdo�n�J�-�h�[q�1֭0}��k�^?�G������z?ℕ�|�����f�c�p���C��*�@��|����5��,�M׋����Z����
}N�z�Q��k� ms����*�(5�L�0*�n[���vB�T��%s-j��ͧ�=i2djM�u��pV�jEWJ���J�W��l�M.�UY˗q����F��0�YzյZ��[��n[�����x����M3�6�te�<�fw-�Π<%��}�i��co�g�>4�����M0��g�����	�4���ҥK!�W#�w� �O�"��=�	���=$FI���Kb����8�IS$�I$I̒�Gb�Ľ($r/�{��J�t�t#��!G�a&p�9Z�����8��úW����j\�vO�:l��qnhcw��䚈�j�����-�#-U�`ߏ���Tu��d�	z�c)u+�L^�H��}W͸:����A��d��,�B�5�(Ǳ��GO�@Z�8�:	��	%=�v�@�y�sx0\���ޥ�F�;�����|[憶�{n2��o,Z���3�>��$y�F��XwU�.��#�w3xJ,<�\���'{;�AmZ�!Kv�����m��:uũw�.]��a�~|�i�uSj��nM�0~�%�y���Sw	B��[�Đ[zZ���`S��Zj�����2�=w�W���\�d���S�^b��!t�?���1�`��w�/���~�e���S�>y�i���~�C��6s�7�n<�5�W�l�~��c�m7^�V5]s�ᘗ�tk�6������7��0�;� ����-���3��oxyJ������g���	� _%����E������@xy"oL�W"�����|*��r���xd�;"���^�"��x��߃�<�_��|�w�O�j䅈�D�?)�+�_Y��#�#��~=�.���_�\�5����.���g~#��oBn�f�	��� �Y�D~��oE~��oC~��oG6~'���@n
|f�Dg�C��y?}�|�~aK1�?E�y��!��!y�;�	�\ȟG~|1�/!__�~�����@P^_�~�||!�!?K�;��?@�>�
���y>��7D��_	��ȷ�Ǹ]*(��A�,�Vh�C�g��C�r�/��6�t���1�:����2闁Ǳ������d����-�·y�B��'xY��@^�Or}��K%����T�S�,���~�"����g��������c�k�h�{��q�@���Q�	��Q���a	~G_Y��C��PK
    +Q�HRA�3/    (  com/smaxe/uv/media/core/VideoFrame.class        /      ��oo�P��--]�Q��Pg��:���hb!��C|����@X7��4H���P��*n���=��}~��s/|���+�MȈɸ&ㆌU��^:d�z��D�
*Yo�,6
�]���{�N������9�<��"����hN�f(���y�Y�yvnz��Zf�?t��B������K�ֹe�X������i�Tj6������3��v�z�9"��C�w=�Է����S�n�ε�.E���pS�2�ּzJ�A���G��H�3�	�N���e�Լz::�����[�ƿ�e}~Ͽ�*4,�HsIAU��uI�R�@�"qYS����%��r���2X�r��Υ��PH6��dq_An*��\r�d^�m��~� q��8O�:�"g<�D��<�>}�[ O��GlѨ�ئ�3��@�R��+�G�U#�Ki�]��B��q��1����c�G�����0B�H�#l�(�f룿Ni~J&��v�(<�QRH%���d˗�B&E�H�0i�7�~�:��y�3ro&x�-��g�s���	Ӻ�k6��c<�"T�Q{�PK
    +Q�H��͘�    A  com/smaxe/uv/media/java/swing/JVideoScreen$AnimationOverlay.class        �      �RQOA��k{PN�ӪU��Eڥz�+�ć6$�`���r��Kz{�w�$�M�h|����&�<�%�}73���N����)�u<w0����i�{�J����+�U���u�(��>Y���$�X|���8�e�Dp �"H�����d�)5���nnj�L%zw,�H3�F2��d���d�/
��w�d���;N33Lk����
*�QCe+���Ŭ�Ŝ�y��Zq�����Ƈ?1i(����@u�G'��K3CW��2-�:���U�t�i��{�F�C��<̠���{X���2�԰hᑅ��%�U���*��1����K�ID+�ZK�=i*Sz,5R��.�.��i��v��i�);��6v�{A~������r�x'�S�賏9E���x����-�&j��q�7.�o��$߱�%^�?�� X�͓��?=Q�}�m�|FX%��6�P� PK
    +Q�H3��S  <  =  com/smaxe/uv/media/java/swing/JVideoScreen$ImageOverlay.class  <      S      �Q�J1=��i;���j�.�Q	�\(�vU)T(tgҒҙ��i��`\�~�x3
�b �$7��׷� G�fH�=���U|�`;��#O�J>�pO�J�M�?��=�ʠ�R����<1���G��te��&V�d�>d(&�#A���tb�X��"M.�qH�R�ҷ�1��U����ag^JL�Ÿߗ�t�|���C*V��������ȿ�=9,Z�b�B���0Qְ��R��U�t3p���/e�|_�͑�"ї�$R(i7Z�k��)���i�7h�K�4q�~B�ޟ�j̰fΰ� =�(~�u#�؏��o�M�M��PK
    +Q�H�,���  �"  0  com/smaxe/uv/media/java/swing/JVideoScreen.class  �"      �      �XxTյ^;3�3sr� d C&
Dd�AS�M�H01H�4����Ir�<������Vk_B�"�d�R�Z[���^������������>�̜L��������k���Zk��;�y� �`8�c� 8��]7,`�,k���q�-�2p�hPh�3�l���5Ӱ��Qé-���5{n��]�nk1�l���&�V�D���\��բ��[����S��8B3�������-�o�>�X���*Z�v'�׍Z���d<���{���DT�jS�j�ZXWk{�V�Ek�fC�j�y�v�����n=�W���v��c�����1�Gդ���Ҍ������bvKT��23��x,�Œ��x"ɠeԤv����=���&aK<�+F4>�A�I�4����6��$wg����
y�[L��ߑ4�C�KۙR#��^<�^=٤���ވ>���I%��5}�pZE����zB�SIܞ��c���~/�(F�Z�g�ψ�bh�\7i�j*��������ڌ+6GT\��F�6-��+D�JW��rͺx�W�K��,��kz_?��v/'Lk�tÈٕ���jO2�����1�#խ��s�S'�?�_Mܦ�"�~���MBZ�c�ԈƳAY=qst0�����xT�ہ���Pw'k��#D,����K�g����q�Es2d[�̢�l�/+��4K�%�d�.�1�Ӣ�B��!��۫Ǵ͆K��LF��=P�6�۫ZX���nR��)�B�/�e�!wJ[<�Exs$�H��;0�#�F}H�lĠ��jt0�	-�f�d��눊�ڦ�I�e	V��I{І�uj)TTے9ߒ,�U��^�%`����~pO{��Wk4u�);�d����.��4r�;���?�Tcthl ?ܥ3��R<�i�����G�15߬S2;c<�YE��G���~P�^�[��l'~�$�&DF��BC� ZQ��tb0#���G�hfjn4t\���"��Px���j*qc_䄔0k�I%����c$K4��8�ʑ�Q9H�u��mS��h*j�8���	�#Y�/
I=I{���#z_,��Tf#�]��H�nd�l�zw����erl2�'�IR�Exa)<�ԠYS�.�K�İ����b�~�fvoᢦ_o}떏?��J	�J�`��$�`�wH�E�N	>#A�[%�&���%���#�v	T	�%� ,�&A�}�K�Ů�uf�j@��ή`H.m�Q�f��ǁ�9�9eh�/DH�����%.k�X1B��\�l!ן˵��|�g���5�ldw�)Hj�!�n�o��5���O��~SrmK���<��WX6;�ri$:�.j����|tS{N��z�D�r��|�-:߾v�F�����xY�PM�3e��l߶�tE`Vty�}�����޺��҂W�o�KE����K�,���%�.\$����
�1֝��3�Y��&��@�]�
UXzxڵw������T��3�.����Kߒ�N;��y�<�>#�g�l�b/��"~�r���t�+9�8s,ޢ(yͬ$hi�D,࡬�_.^�7�Z��ri;:.ع������<�^M�s���YZ���e_�6�y�rH�	
�@�W�_�[	"Q��^���I��(�SO|.W�z�{>�^S EP	�+PC���Q�I��#��WÛ
$	|�=��-���I=�3���YV�9	Z�
�N�\
4�'�	����@-�*���%X��	���H��	>�1(V`1���2�	'��(� �|('����PA=����
|�U��	��S`A��	�B�U�/��
�H�
��wh��U���3���_"��ߧ�(p��������_ЦA�?V`9���R�k�W
|��,�sVl��T�F�[>G���z�&��W�*��&��������B�o�N��Mp�������E �	<2A�BPBPF0���`.A��`�|`�8hB�^`N"K��/�?�+�������FF�.'XH��`	�r�O��"���z�z���kn$h$XG�Dp3A3AA+A��_/�!"h��0��.��(�wX5�2�Ȯ"���Z�6l&�"�2��6�*�ˤ�i~��	�$X*�Qv�gd8Ʈ��8��'X�'�
N��n"X+�8[F�!ͪd8MJ_5��`eL��ۊ`�]AЁ�����r��BŠ��ŹE��p����%ӌu5�������ɔ�a�>��i����j`�] (�gq�E��>�ko�6p,F��^�X�x�����?��v���vy�����vP�M�1�3�b	��1orO��o����)n�6�bu�m��c�v)�XC����AΓL?�{�j��V�,⻃S�k�������+�B�烓��A��!K'�]�i8�5�ޚ`�������&�'x�%'X��۱��	և�ʝ���Iv`���7�&X��T�nF�;p���I}�l�`�ԏCi�X04��L����n���
��l߻8��Fr�6KL;"������7e�kg��.���6����.��
3���c�]��g��"�Ψ�L����*:(<�o���l��N<�pfR8�$��Ĥ�����B2d铣4k)E�5��0ɾn�|���#���YN�y_��+M�/[���I+Ĥ%�� ��ٝ�hv��5;����l4͞��>��b�e��9�`��3�QdI��d������w�/���PJF���6�6;L���݀'GnZA�쾪�@�z���^�s��?^̃C]U�I��/y��R���PU.,sQ����L�kp)��{L�A��u��r�:0��b�B�a(�����n��w���>B%}�����
XBR�s��h�ۺ`����doW���O�7������=b�J���x�TR��}Ө��c�_��5��wF�I����t��C�j�s�?�j*9��)�?(��H�������W�]m~Uv�4;S����n�;��9��������B�u8P��ud�`�_���F���&�Y����FmG�f�<!ħ��/�%��۟�;���F�C��^�ހ�]^'f��p�>Z��4����p���l̇\oa��i��0l�D1�ބ��|
��4{�s�$2�>W'����"�l���|�fs?2dS�p�+y�^�WN���TJO�w��K>�4;���l��^���>�8�s\c�E�{y�C��8s�}^�_@�G:��O�%q����/�;���VI&����<b���e��>y��e\>y��f�ri7[K���,E�e�|ҙ��ﰏ�;i���<��E'�D��^w���/����F�3�sR��t��FI�E��3u����[�U�u�"o�����+I��u�hl��
oi����z��%��{{��b6v��<rQ��^Bkd��wƠ��ˣm���x�YS?�0Lz��f����W�[b��沙d�A+%���֐�f����T��Eb�NL�Y5���dCUf]�t�M1�ٛ.����3����n��i8څR;�3��XW(tf�M�d�)v��&Yښ�$�fxϞ�>J7�(:�P�����3�U���10̝-!�>a��Ɉ��}��c��.!6(�����b��{�kh
�<�+:�dvi�a��Қ�m�É`r�Q��3O�l=@o��FZ;t�+��߀�m��_�S�zR�8)�%MG�^源x�GO�1�(�xDt�b/h<z;?�=6�\ߘ�ۖ�,�� ��`/�}��c���m�<W���Q�`���vy�=J����;���1��\O�3l����]��d�q�����(w�w9�ڻ
����.W9k�d���$�����	�QV�t���n�<�Z��4������.��\%U�i6^���� ��\8�
�L���L/�N�A�}2�xI��jx����J��\���}��|.�f7���~i�\G�3����O1}�w�-,w����1�N��i8��pL��X́O�S,)�V���U�O��遼��|�PK
    +Q�Hf�i5  �  5  com/smaxe/uv/media/java/video/VideoFrameFactory.class  �      5      �V�wU�M�L2�PB�P��Y(A����M!%�J�5��4��S&��L�������}�+���~��x�LҦ�*=朹���~��o&���m ��Wp.z�C�Q�`(a�1�`"�\$nK~K�\�ڒ/8���I����ZA3�I�W�,h�dA!sJ��,f��"���aF7
����wg�|��W�he.�W���%5:�eUc���	]4��)�95A���i��UG��*�:^�LeJW�)eS-��i�R���r�yJ�r3� ��3j���ȓ��Z�$�w��`�R��舡H�}Y���T�DezZ-��D޲��TLņ$���VR3怡�3FV�t:��#��V��ꈶ��#J漚U�E]�[��Ќ��R�X1GM�L^���������67���BF-��Q��6�k�u���6��W���Y�o�jt���]��aw�)�٢�#�J�&�X���E)GS�.+sTi?����bnYa����j٤j�h��Ȧ�<\����,�Ƽ�v�<͌*�~[D��S�.�E��-�!�xDDPDHDXDD�^�)���I�	ؖt�l�ϴ�MW�	Xl,��(L67+6���kE�ܐ�uCɦj�%r�l�2|8���-���0�KF�3s���:�t[WbcV��*��&`_K�w9nn�}Sb�5T���3��n�7�Կ����hi�9��]Iu�k��[M�ƹ�����+��GO)�kϊp��j�����K;��-Mu� �Al��$��h��+�IF�28#c<2`�^�1��dD&>&~&�{��|�,K)&#2��)���8��e<�q���H�x2z1��9�=/�/�ËL^b�0��&Y��y&��&sL��"�f%�Ce2��5	GaH8����u	'�K@I� ^�G��)a3L4	�������a�3yU�iЛ�=@�����g�L��#<�F�ڑ��I\�����iu"a�P�7\�}KJ2wE\��K���X���@��*޾
���luc��$`����u�YÉ��q�����v�Riw@H�=�p'U��5e�,�U|r���K����O��.x-�VH7�=
�%�T�[8u�ra�!���!�g��=�!���t��+��k����7�U_�q��z�N͏Ӂ_�q�&N��ᙺ���"u������$���-X���'�i�F�n��/?-��a ]�`:���*���(��{�������
B��+�vD��!�l<��.����8IN�(Ƹ���~��8�CT��Vq��z�:f��Q���"Kx�Z��ZX�Z�6���nm"�E����hH�{I������w��D����9�vQi>����I�PK
    +Q�H¶t��  �
  #  com/smaxe/uv/na/WebcamFactory.class  �
      �      �V�wU��d&�)ДR(��M�-�RZ���E�ɴ����̤��*���;.u�Z�ԞӃ_��?��w���M��%G�9���~�����勵����Ȋ(Q&b���"n�[D���Eq�88|�[ll�񨍽x_���h,�Al��4]�9��N![%%JI$T�\�E8TE�xȌ+�j(5ҕP��Q����e$�8T.�Ǵ�PX�o����V�25�&���c�S9�1��c!I��QʹL�T���4b)K�T�A%�t&����(�D�\*d,*f�:j��4KM*�ϐ2���+�l���ꤗmR3B�T�mL�B�#�*:��׹��!5b-�����й�R�RZ,�&����PnS)K����I�oZ��m��b�)���m��p�����7K����C�̌g2�Ֆ�i啕����"�]&G"�ܘ�����J�J%�nSM(����j������!��۴��evk̋�L���B��)=�$#���b)��UٔY�|�x�Tw�T��A#N��a%�R;�)��u�	����@N�̉XN��+G4=j��Aʐ:���e�
�4��iD���N@����	�	�.�/  �F@�������4	�'�Y������^��z��/�zv���z������-�ssDt�o9��,6/����[�_β+^���̻Y4X�ȳH����m�cE�,v���,d�+fY<٭�Q��"��]����L�R�jo(`�~S���8��:n�-�U.4��L6l�Is�F�4����#��j�=����iO����˸	�eT1����Je�c���X%�f��c���xD�=8!�N(2*�'�Dd�e�ȠQf�ʨC��-���2*���I�"&c��N��S<� )c,7Z�b0�FF$Z=���J8��%R�1x���^�Ўg$t�1	�ep��^�p�)��7%܏�$t1���� �Ѓ�$��	��<�'<[��x���t�<����j���^�fC�T������.m@WثK���c�8��gh��W.طО�Ak�5���3؄�~���p�E��Y���m8���8����vw'f����2�l[fq�g_z�,��`�"޵�,a_M����q��3�0�R&?p����g�^w�c�>��%�'���*�<)?�q��6��⇶YtQ�o��W�4��,&�kfp��.r`�f�#�4��j���s�΢��뼈s��~VP�k��N�}��Ҙp���R�BTC���������ݸjި�$3r�/��[-��˫;�+fs�W8����s����f�ѱ���Σ����Y��:Age^�t2�"'?y��&���,8�;7��#�ܔ?���h��pm�����s�	����E�8ȷ�m�:�>��<�햺<ܔ���ةS
~������^O��$CŃ{��i��|��_yG+ص_V�i|���OA���٧z~�(�	��7ϊܜ]�YWh �PK
    +Q�Hiv[�  V    com/smaxe/uv/na/lib/Lib.class  V      �      }�MOQ����t�0��R@�@�--~��h"I�
Q�Iu5-N3tHg��?0qC\���#��D�0��+�sKk�Vgq�;�y�wΝo?>��=w8�A
?�I�"�ߊ�w:g�!�g�.�� �L���9kM�״-]-m�M5���6�����M�����9�$��b���uUwfMͶzI�]�E��kk~�Ot�*sz��M5,u�����兒�^r��F��u��o�R�h����6�ªZ?��In��uǰ
=M����9�A�����E��%x%���-�G�OB��� C(���%��v�J�n����8-��@���$wG��t�QP��6�6��)��L�ă�C\
���t�"W�(QЅ�qE�p��q��B\� Fy���ja�2����+����Z�:��AzhP�$�jӁ�D�о^��\{�
ѽ���w�%�C�gʌUq�wU\O�)1wǏ*��L��]t����O��N����1�X7�bH8FWH��6��XJ�e,$���ƹ+�𴺤�\�y�{4�9��1�aY�D�M8ؤ���xU�;��y���o��.�a���A��8���E
����
��$��L.~�u��� 1ZEr�V�ҤYK�t"��b�#&NL�PK
    +Q�H��:1�       com/smaxe/uv/na/lib/jitsia32.dll        1�      �|U�0>I��L��������)E)��&t�W�laqmK�4�NY�]ݽ���ʲ�Ww��˽W��+&۲�Baݺv�S�j]�)��y�$i�z|>���/��9g���s���:?[��]���8~��q�������(���xe,�B�+:ˏ\�*�����[�g�]���������`�"�g��}��;|�{�_�����<G��<S�|�l��X�ܳ���s�Y3�O?����|v�_}v*��w����8[��7$�]��+�ww�h�z8n����mE*��3^1Ɛ�q��D����b�X�eI{6r\g`�;�Π3��vX!�^D�뷽wz|�h�Ϙ	(V���y���emt����a����a]��0v���[��%��q;�8�r���2���u0��������5���[6l��n���@�7�F��p��������_��2��,}�����??��+���5P�R���_�q�A�t��u��?R���Y尬$鋗,��cq�~�C�<���O4r��Fy�By%�+xe��z�u�G��ԓq�E���s:�+��0��Dx�����&��e�9����ېQ�[�i��#Iʙ���8��yP-w�k�&�r���Dr�pj(hS6"`%
�c�4ym}G��k�������+��,��g%�|^���Z;��[Urȵ�q����`\��V   �s�n��,wW�*+|�N�O�t�%�w�c���a�?��*+�}nb���QyY����φ5M9(���\���@n5mI�N�j��� w%�~*W��,wL0$��Ƒl�5C��j�v�s��qүJGx@l}�'3�_*[��C���ڙT���4��z̪lin |�*��a嶭�Z��ղ��Ur�I����S�8�Q���F+$5�@Ĝ]mzk%��&ɱ@9h6�I�4��xXe�{���3�f 
���c[�x�MV��s�����λfm}��3J���j��Ŗ����W�
�u�W�	 ��Cn2%���#t��x���D�Ç�/�8>�<D�_�����+v��1�մ�p"�|/�,��� ��aȏvYm��v"@�韦3����E�r�xD~��x�I��z�����!@�~xm��<>%���^6i�B|��7p�aO�ӿ�4!� �_;�~������3�$Nx������a�&'Iv r6ٵ���lk5�[�,/��P�;+�T�"zy�~���͵��L��XG�����;��%P�k_`Z�Z!�
Wڂ�@8�s0��k��z w v�a��J<QW�`+����8�b�W��+���t�EM�T%��z@�N#J�CH+RdG9uM��,g!��'��|A@(tK;ʨ�ִ2�"*����q;�>X�R���nB����	��Q�U�������v,R������:�dgT������j���gU+�j��������i����J��C�J?�bv�
H��H.����t����O
u񅖼����K�O������]G�Y������U�ؑ;�+��ڭyA� 8����S��k*�B*yluA�b	�%=aI&а��!O����͊)����|@(ͮli�@�{�t�T&����1�P@�R��`Ps�Xu�U�B+�39�9k�/͙�;�.�B����L~���H��T��(0�i�88%y����9��x�}+����}m���Z9��r�S�ݪ���>�$~{���U7Zc|I���5i�����t2�r���/���d+H���5,�gt�r��P��Qm�����I;5M�|�/c�����F� >�Q����u��3��	��"��2X.��(9�,4�J. �%h��� �+�>��y�L�����<+hC��#:���K����7S�z�w$`*-�dHpK����z�<�	<�T���r�M�B1� P�H�V���:W�4~6�ՓS�3,ɬr� �~M��+���ӿOBVR΂9��6q}Qȍ������DZ�v�\��,���N7_�����E���/K{/K��,m�,m�,��{���{/K��,����������e�7e��A���F�cKE;|��oFM� �|(�z���R1�ޕ��%,�1��M�{gt��c�,� h?�L`S��8�|v.���a�/03��E5 ^H�n��2e�41�2��"~T�uO��%�B��:3�+g,h���W?8a��E�iS1������+Ⱥ��	�DF{1���rn��+-q�'B�2��5����d8R%��1�!�ϟԋ��T�fs�
���I�J���+M����T`(T]!�����A0���fg���B{�q�(�俎1ÿ�����
;b�� ��|�=n+D��L��_"1D�>�vT�,Z>��틼����0y_(}x�tK��iYbwuIח>\(]���������q��m�k#�$>{���u^��ymc&��}�Mf�� �bӠᱎ�l�`��������&��̝��XOMr̍�wp�qZ�J�n�1>�Z� �����d�,�s�XWe�d^�5t��ٵB ����DI�\�h��W>�49�5@$ƈ/m_��z��q���r�f�
ƚ k�����Y�&M�ƕf�ROL��U���#�m>�Ƣ����s���+'�BuI%DV��5t��ԧH� uG΂�;�:�!W�Z����-��$��eZ�9�]נ�נ�b��l�� �p��,�KRS.�z.��.�G�B�C�F� �n@`n�Ӊn���	i�g^�,�wc!/����uo�sn��W7��j#����9�����2��H�I�Q����d{�ɛt>��;�WX�u\�ʐ�����E����q�:e���D�ϸd�TH�q��HET� T���W�G:w"�WϭW�ZH�_2�0`|���S�ԛiS��ĥ%j��rQB4��Yc�t�O��ev[��V�ު����B�ޮ���j�l����,�`�bYl�n���ׂ�2���L/�}c���)��bs�%_@dvj�=�MV�����ޔ̤�J,�`b-�L+f=�qyVi�liL�� v�Ms1=w$���c$mǴ}$môm$mŴ5�&�`T�_�@��P�0�\!@D�6�]�4�m�T��$ȟϽ��d�j����O9S����}�!�y?�A�Q���g.i���O��Y�W�i�l����uJ�����&Y��#�
�s��1�������]Y�H�KȲb��:�^�6� 1�x��(��b�-�T	�4��[�܎E*��!����#ʱ�zT�E��fu)�O��bB���^P$?�%2���ւ �uU���r���`��ھM�P�3,Vo����P]�٠٨��Р|tP�H��&G;=C�6vK;��x<(��?�iN-�?������`,���S*Rsze��4S���Q�`�DYȉ�.� �E��d�����,�[>2͆�d"dq�f��-0�c֌��D�����$��v�3qd�.f��py��cL��4����N����5�~x�  ̼O��^�c��0y:��|I�l�C�*y�T!'��w�t<HT9��V���Z�}����`�4�qHz7�%�b��������@#��2��,����Ї{e��Ƽ6�t��-��ٿ�[8u�*�B�@�� ]�sr.Bn��sztԞ&z;�$Y:+��sƦ��v�3H�8���('v���?n�@X��@7Ú4A ��l�P:dP�d}�eOX<nVb2z@����d����L#���L��)�{e���B����Cv�md�:��ot��_��w��W���ߣ��9?��o������n���߿�����g����������T�T��f�ôf8LX�`m!cؠ43ɯ����$9BԴ���yw+���o�>������&3'ekV<��"?�,��Ҝ�rq֑��]��H>
Q!�<���R�`W��rC8���3w�o4K�I�\ o��a�_!������*����i�^p�x��4�G�tB�n����"���yWT��K_H�t��T�`S�����#��cH���� tΞ�M���uq��2h[wR��9h�]I� ��w�x䶆��c�+�����8�W���ؒ�8"0�W��m�EI�����l��Ҹ�� ླ�=�m��,��k�C�porl���Z{	1 0װ�`?d����<�C���G ZE�
�A�M�J�$Z��j�M��E	�s �{� �s]_J���Gi�Mk�J��f�� ڹ���x�ډ��\R�*�� ��	��KK� jT�R+�}H�H��������P͓n.	��q�<C�!�(I���Z�Ṏ�A�a���/���������~��?�捊?��o�?>�͠�?�I�����.{���>�����T��&Mz��é��_�7� �Ҥ�z3�qd�h�H��P�
��^����_�w��Ol��Bg�#�Ć���U�d%��1/�����v�� l�6d����̢�b����w�/A@`�{��<ũ�ei+���Lg�ե�3�����\���O8�}M���Ҵ�����3�������p|��9>�K�=>~�������@p69l�?[����V�>�;[�0�	��%}
���~WcAz�@�m~Ť��/�4�9&�ˬ�/䄯��5�i������16ȳ��n��vI�� |zg�%,N���]��)�1ד@e1PX� ��r2���{�\�q2��:/�Cr�[���̅<`L������]#3�E8m��>�1�2ذ5�y�2�D�ɛ���v�h`i��~��q}�#�0��d��8�e���.f�%B`LT��@�����?ؐ ��s�.Ϲ�8��g��'��3d��!Cg�S��V?����L � ����r�j%���:{��H9��/�:]�0��t~�>���?k�9���t�86�ԹT0ԯտt47	���m�龱��y��B��A����S�ٕ���+��>�1%ͨ�, �ai�xǐ�)x!?���+x�v�e�����aD�䇎�!+ŕ&�2��<M}8���.C���svi^��u��X��J,�Z��z�P���ک�Zw�}]����#x͕�fQ6����0~t0`��TY��@+7u���	�A�g��[.4��*e=s!8�&��_E��5\�V��M��w�
7��3*6)�-ל}Vs<a)a�z_*}���c2uk���	�#b�׻��KH�*��:���o���출�
C�RC{�ж-5*�&��!?�F�{�A�N��eD�IC��a�N�Q���-G���w���~���6���Ê������������p?�sp�� ܇�>�#h�L���74��l�ïs<B��C�]Ha�^�d�8�#��lD�q(�P:�l�H�_:��|�7����N�9��7�&�6��m����	��s/�̐h�0�<޶Ԥ|Ƹ�9�޿g�Fڒ0#m�@�Vhˀܕ@#m��I�IA��{܂�����k�_"�ߞy�m
�ׅp���w+ܭp��ߛ�n�� w����G��Σ��� �ކ���6&�:�-Xzt;d�j��-�$�����G�11&_O|r(>�����^��G�/�U�YV��yɛ�e݄��?Aȣ�C`�p"U��BD�}x����Oqj�p��v4���P���D{�>�z�7�V����� 'H9�8����ܯɽ���u��Bc��|h;I��t7dr�j�`����-�e�,�3֚��~���@��v٘wu�"�k�>$�H�9���0ە7��P���]O�k��i�s���&q��6�x ò�n-1�|��8JV?-�yi-~�C����!k����qNMm�UO���G@��P��<��`#
Ɗl\��[Z"�n�mV$?TC4�kr�X��1��%�恘"�PZ#���6�LԤ隧71��Q��1�$z��W�)�A�Ű�"��Ԉ���i�{���>�f�H��QA��^	D�4���@�gX�x�����m
�l�T�O�����(ZS�XEy�kUOo
u.�P6� wJ=����;���O�u��(��E�]q�F�^[oJ��m��:��^J��F�j
�3�Ժ���f�|�>>	�5�h�28,M$�b_e�n����M�'z�,���;���"�����V�����̈�d����� ݎf�J�\��h3<*U�Zi]�<3@��K�#�ק�� U�AW���Ӆl	M��L�hr�)ˑ�x�g|7��?d=�s:p�r"��٘C:����'���ۃ�	@�C�_e�E_�"+4eu}�y�eě�bͯ��J̮�[.�`�4|�;@ȁ�`��Xg�����f>Y#�:%����P|18j(�p�`��P���貳�;@�6�E[�2�Y`�s�o��ex3|��)���옥��	z۲��5���)�v�V`SP_����Ak�D%j1���-�:<�x�J��Ջ��`5wŶ�(c���3k;4�f1D��Xq��%�l��(/X'$�0"?��5p`;
�I(�L=P.;��gNZR*�0�M����Y!�S�{z%*�� ��v�82�,d������2Y�'�t�&�l��r��!����&�H��u�q�W����J������HL�k��q��y=���9�dW�#�:3�w��=���A����x�֣�����<6� uy�X�� ��<�����N�̓&Ufu���1�uC�k��>�8D�\� (��g��� 6Ū��Q��˰�v�%8 �/)�=�Q�
�y�6~	����6��͌�X�m,��V8%Oʙ_K�04O�q�<0�gpF�}{�n8�uyNC>c]��3�zz����v)ND{@̀�~e�9(3�!N�pN�wP%P='#��:;�<�����0�XT�1��B�hnf�oG<�qɫV�ռ][�l��<�I���B�N��$��$��x��J5�2�RpV��� �g�J�F�(z�]n���OwbS"�o�6���ʮ:��#�گ]�k(!��<�1��%�r�?��I�{X_��B����|߮���F��0�_j!���s�aM΢�E8TmYA:���<C��|c��Rh����Z���	�,(�f��g�P��1l���y��mYt�HG�J�35��e�k�}T+xz�Խ���KW�AyDpU	Rp���uq�'ō^�p��b��qt
�W�j��A�K*y��Hb�v��������[��'��h�5t�!5'vpA�����ʺ�<g΁r�U���IѢ�%@�m��n�;�����I��H?X��w��Z
Q6f�Ӌ��oi�(�?��,����A7��/�3-V�h�Ǳ�g��[��2=M���D�^��T{z�<����p3��~%B>�C�[ �M��Ř�n�3��B�͢T���!�R}'�x�u �!�1ݚ�2�oj���Ni�ap< @?���J-�H�fB�����V�:�B���GP�5���| �u�lf"��Z��Z���܌��%���b�g�y��<3�*�O�(EX�`6d���
^K kw`��w�b�$��-`�jA!�_�q�3�c����;9�Ѩ�� +)������ht�(_���8��l馧Wi���֟r���G���ETlU�Ye��(�����>z�B��N ��ĺZ�L�,,|�
���?$�����L��F�&
$�[M�[��L��&�;��o`vR&�h�痠�
8&Pc�g�au����n�#�'��hk��QM�W�蹙��	'�Q �o3&�L�>��]h3g�[I�;�Pd\���S�ԕ��@�Ht:�kS��n+{��P�P+8�8w����C �A���SO�	��wD�����r�Y!s}i�l���|�������4
����p�'a��! �#31@03�=ܟ���awYr����5*��3�ϳP�����H�+��p��ү9(1�y�`h�(Y4%oj��s9in�$c�Hd�2�sb�Ȣ��ӥ��P�	����X��X���~�bwl��ް�
J��.LԤq��<�o���{X��fM��Ƥ�j��,�cQ�%^�����<�]�`U^@�����Ҭ[�2�W��J�b�r�"�<2��r�I��[��ze0��h|����%j��?��N���@�W`':}� n�~����r;���U%fL�1�h93��c�C��Z`��4+^�Y�Zf��Ɲ%�?�ݦ	�ų�U�]7�z걬"H�������p�x�=Ř�iZW�f 5pn7���TW���<��*do����B��"�y�x��r4�A V&������g�8�� �2���d�	"n��=�VP�]�x�t*="��P֎+�}�#mHd볿������.�E�9��v k�ZȺ�.�y�m\�6Ë{ o�����A�۱cs�E�"���6yH�2r<�)�?)�{;r"�,����ϕ�D�Ab�>��O&��"���~�|;z&)��*�.�ϯ�_[�`���jr 0�m��Q(*峵}c���<����� ]���C���u��k�j�b��$�?�w�]�iA�ϹY����>�2�擐�u��Z��A��$n���[Dv��vfjp���.d���1��wh6$�}��S�{�u:y���F�G�q�d��!;�=Cwg���|MV�}Ee�=:P�gP��@Yi�]w>}K��6{q{ʴ#�K p��������#=�=�4�:Y�<L�~49L�cC.`d3­��)@�K�2�|G=�855\�pw���k\ѽc|��l`q�<�^7lo	�0=�{q�>�@p[N'v{�}�B��k�{���K�C�.�O; g[�V�6_0JY�������i�M�e�������7-�\��vI��fzэѴ�O�r3!�>�35����Ylōc�͛ ǽ	:j��H�_��������V���<䊉�� �Js	#Ml�1�Z��i�V�U�s�)���Lp"j���0j��I������/䉏C�BH�lS�����
ڽ�m5�ڪ�T֕p!#��%n�Ǽ4z�>�x��7�a�Eq���G�� .�|������A �����h���Ԑ��y�=�>ݢ�ʊT��"���j��Z��Z��ۏ�ˠ �EXm�~����R��i˙���y FXaAi1��0�N�>,(����W��Q�2p��H;=��G!�7V!�ν��_c��0[`��F�
�%��2��)q�1���~j��\��<�o4nt1&��e��Ԙ�S�&��ګ���up!���с�@�Tʾ'>r��>�3ǶO�a�V��d�Z.��}��<��Y����ͯ��pjDG�*?���*��K(�o8�0A��+�ꪲl��>a�"�il��� �gttr��6���eX��q[�!�z�9����z��on�%�9g`��:ŝ�����0��ydT��4�F1|d4ѕ8o�,�h�)G����#�Kė&�>4��W��)�}H(�F�FX��ӰQ�׍�����*>c�:��5����5��pY͖b�ng����MUI��&�˨օd�\�	&�/�70�7Ū��+���yږ�s���@���'@!#D;'�$�����컄��i�Iׇb�ϒZ�����FZ�a�ob�d6�C@ׇ;�H��^�.ڐs'a���tI���-X{��>�ЊK�ht�*ϖ3!feG�W���MʫF�.�U_�TP��w&�yG�G�8	c�ĭI��7�����}Fcs��wF�+�+��ӓ���A3a��aJ��T�u��ִC�%E7,��bOeX�J���Ҋ49���{��v�5�$��-S�-I�#T ה8A���"tWwV�dF�l�#�//����=R�~� ������7��;f ���Ә�L��Sի�"s226bLP'����`0���G&�=�UYE��qP����?lL�|]51�ƻG�x<�7B�����Z�lVӣ>:�ʨi6��F}� �S��2�l��X�w2=U��U��@������k�T��Y�W�p�憸GY��� ���E�/q,^-	>#��)]6�`]R*�aG�[�R�Bx�`��_�G�� �~���aM��4A-��[��5��)��,��Z���R6y��F�R�&�>Z���1����s��jc��T�4�C��j*�1�lr����Dh�B��\:��]�{C6z��Ʒ]e�*֑�o�ʣ�9}�t�<��"��<)@�����HR�zcԅ�� ��˃R��q�z���,؈�5Sr�/����AOh]k��k�����{}�e���qQ���a��oNOj�ݍ�!��^u��A�J��z#�~}.N������utթ���?��hv���Ǳy��N��s�͋<l�i�|�u��t�K�S��Ya&����!�p���dE��P�7D��(�Zu�GZY�E�5d���H��\�N�gY�{�'8��v���8�~�*mn3� ٣I��$��H���2�鵋�.�{"UBK��[�푯Q�J�rN��N�*M-�ItBWB���2C]�dC�������Δ�H7��٤jP�4_N����Tm�4T�R�
~
Q5.��J}f��xH�}� i���6��51(Nv��^6���g�\�^�vCz視un��r��l��� ��]3A�n�~����v���9 k"֐�He�V+lj��'����lC߲�l�Z�ֽ&9�<2�{5����h�+M�ӷ{4�e�YCu�h�@啍W�1o�'_t<|�n��,�H�&u,��+x2֕/ ��x��
����r��b��uI���)�r"�H�h�-lrܛ��U��lą�8l��l���h`��-e+�m�}�f���h�,�V{��8���Ύk�:�8�]�~�t��C��PCvbN�I�țt��e!������ke����V�/�W;ީOM��n��?��Y���� �w4�#�_B<����i�fS���Ϯ�ٕ��1v�=�vÕ�$:�s�^1��|"��{/a �G¿�)�u�/�����*�n��O�Sk_����j��&���,6[��MB��T��3��q��BV�T���yj}��s�5,��O퓜��}�Y{����=�9\[O��� EK�W^�~��;��ս�{�~P��7���#�@��[cQH�rb�|�~J@������_| #�+��.�9Ƭ}�����1��C��=��
�K�)�$�W� ]UY)@Jo�5���B�g��>�l�[	�-�����_�n��毮��*q^oY�fH}i��4b�x�e�e�bX��ߏ���)��З@��a��z��him���<�ۇ'�0��DȰ�òL�i�*(�7�I�5��~DH����"ح��K�� �zs��R�[�����}nxn�Y0_�޼�P,۔.c�ls�l!�,p2��t�g结_� �z���x����)��[��wYl� ����x_-��!��<�mQ?�W|񀗮����Q�j�+I�-���&�=')����W\��	� ���]V׋��#��!�������2��_��$��j�	��bxg�+�҈nU}�W�ȫx�[k������)�	�Db;�]���Q��@�<�
E�>1��|M��F^�y#��&g��L��-(U#"�����9���<f�V��L®]��`%�Ɱ����&��Csbb�Հ�����럐�ė�y�X�H+�&x�l���]̼�Gڗ�1�.Ǣ�֩�GTLi5puJ.��<*��ƺ��qj�%+�(fT�S�3���{����O?���n��,>v�5�i��e���E����b6��=�e�>i�2x��'x7�>߬��+�������jj�3M3=�!Nq�!�J��bvɼ��Q�6��	AT�G�w�Oi�[��m�q>�Z&������}���bp0���{�uqb����l�"���W�����:<��>f���-X�ؔ��d���&�t�{��l��������!5��IWI��f�%�}Fg�>�@�D���sLg#����X/�`a�Ǩa�4����$��6�(	[[��*�y�l���;p�u�dc���z��Q�h������C�[��W��\����F���gN�j�ƶ0S�y:�����*�~�	2� ��[>�Z˂��1����]����A�"��d(���<�� \�Lӓ�O� M��1�"ڭ�ΟTNp�?�\RvA�|@e��T�w��9��0�{����2A�����+����J4fM����Z����?���P�u��O�bA>P.�6e�7�ƮH���Y�$�^X�
��~ϓ#G�K���Ɣ��k��ȝ�u�F��Q�F�Q��&~�����{��J�,k.�,7�~���_R^E-�7�!,$�9�t���.)Wo�����ĜĘ��8=a�ۏ-�a.{��=��"V������b�T��.d��z/��*�4�k;����������G"���˔-j���/�HL֑A�Yt;�>
ݩ+�2�GIR H��W�lo(��#�gP!nW:���͕g��li���R�α�fjA��'
���!k�D#�N�p}�R�*�X�A��vz߹�ы���&h,&����������sژ�n�A��v���9�~����a�n.q<��yd��8�E��w8��՜���R�Y6����?�\�z����^�@�r��'��l]�!WL0��}�Bײ_u�l��D��ʋ��.��婕&x���u�������2���^l�d�p�n9�l,��Dl���8�b�G�塻`��GH�0�>l0�K٨S��_�RH��d_�Z��w�H+��m�1I����5��Ѭ�sr:}p��q7pD�LG�(��-'�.^�D�/ل=95�-�5�p'� ���܁�A��	�`�f}ܨ��W>�A�b�Y�O�M��(�^�g��k���K���M������u���j�!�ņ:O������ܚ4��ݼ�oN<�Y���lf�V'�"Kؔ��pnbk#���aMZH��
G�ԅ������:��G�k4Is��D�ue��E��w�h�͵� N�E׮�?�!�d{�Q�mi���WD6���!N��k8tFr�Nw���8����g�fz�ૹZh��}^^;��g�?�LO_�Fu)��rQ�r|���8��,��s��p������܌�f�3��p�%}L���'�0Sr�	�	}��K�>ӫh�6�|b��"g���nvd�g���м>�3��G�x5�GpE�p��gY6��e��1�t�*�0ZΤ��82�/"�0���20Z��&���~�
�cC�k�o���O⹨?d���Ձf������`dmz2�T��h�m���r���^/��>�Ak�e�2�G��H)���E��oʅq�密�Y���qZl��{jtfL�
uq�keKز;�M4X���SY��,sj�ߟq��J�V�ͫ����c7�(5ނ�H��O���\]��Tm���vd��ƥg�@bI?}��m�A�\G+�g��'�������Jb:�0�"QsK=f鿉-�cY�v����R����˧���Lk��W�Bo\Eγ�楅{%������n��\�o�<��fm����/�F�L�Q��� ��d�p�����Gw��/�6���ң���q�Ksr�'Xx�	Y���b��F(tc�afA+@.x�:R��.��O�	w�y�?e�bN/���x=Ύ��Տ�u�ABT26|H2jǕN�%���I�����'�N8�i�<Ff��D����qg�n��p����[q� �Y:��n�.8�޹Ud6Ϩ����R�6~gm�45�Otu�K�����ť!{Ѝ͛L F�܈3�.�:6�!�������/p�?.��Ϡ�`Ka���..�9>%��1�1�6��֝VO*���캸�vZQwi��7H,�n�b�
����J-�!'S(J�N�Y����X�SwL��dXIݱį�<�n�AKc�r�mB�$#<�|�.O����J� �0 ]��8|�h��k�X�1�v�~�}�5���=��q:x�7+0��L�n逫v�?���*�B#[�H7ऀ>e�m�R�6����Ǟ��` ����h��	�a�Q0I.��݇9���V'n�����_?|��WC�Q��-��S� ��S��<��(�n¥&���)�Al��36����23.C[?����!�ݚ�[��� �V0#����7�%���A���y���۸g�,4�m 3��hdwF��#x:1�Y��dN�����w7�pU�]�~����q��s4d:~!x�y�祛�#
+`}5x2�#Y� �Ӽ$j�YmV��H��(h���v(�����t�>���:�s�Ц�uV�P�5i�3�n^ڶ3K \K�J���*�P�y��<��mu�wAfR~}z:'�v�M���E�V�H|6_g��$���!6i
(t�:�vy���Ztv]7�F�o��1�>��;� ��̍��}��Y�
ͷpҭl�IV<�g%�~W�F���6JY9��w��m�2H�ϱl�t��_��H�pe+�,�f�U�7[�'���ÞمH}���(ft���1�<1�m�2di��U�P�F�_-;x�ؑ-��*$Ld��ʽ�K5c)��Z�J߅vk�r=�7d��\F�HqL�{���+1��
ԭB�Ď׽CФO-:��M>C��s�(�Ef$���x2eP&2�d݊�m�@?��B�ҏ̙�{˜�^�p-%�'%�v�I��TZ[.س~2Y��\��B˅+�.OR�����q��"�͌�汸3�+�ېAΏY�����ܕd�B=��n�F��6ZxXKOb/F:����J�bj�'��Ѐ�:��x���GJ,�D�cM0�R��*g̮A9�JP�΄K�GS=�Js���A���v����"����($�^A�g�K��CdP�<�2c��t���J�F��Ίŕ��Q��݃��w�z�lե���1�:���}��v�]|�����@�ة�j�ai��`ZCs��g�h�#`���ь�H�z��9�tH��ֶ�"��^�����s�N@L�x���y�f��N�:F���~|G��YZ�mgR$ْ�dM.���ao�~|�E��j��~�9C?���-�|�	�4Gd+�Ҕ��;P�A��-ʆ�z\歶�G�d��w��i�k�M�����Ǆj��Y�}�wR
�<��jM�]�7⚧'�u��iu)�}�~t��-�no�� 3jd�czM[2�[�4�@/ �2&�c˘8�1iv(��9y:[gaӻ��p�@G�O���]���m��EO�5�hw*�rb�j�֒jAl�����<V�Yl]�YP9���|D�Ѭ�9O-�='H���i�褛�~�؊�	����!�ڠ]Ŭ��~1�Z>��|�hŅ�m�3�J�捩b����Og<��҃I`?�Q_���ʋaܠ�h4(]B �Ti�&��G�e�� ��J�$�#��1^ �V)�-z�+K%
��7ܘ�>�Ç�ՠ��$�E��I���cA6��}o]zݟ0�����Sl�ߢ�W�"u�Dηט#w�3�d�{����
Y*��rq���Hʯ/2¡�}�)��%l�7?�x�H׈ez�Cf�t�w�7�8ɂ
��N�5]��m�&¤�v�Ʈ��z��O; � CđG�>7��Ǎ�nfX0�W��1Q����S��;�䖅&&[g�:ω�hfg)5A*�R�2�źN��{�ku�7S�@TfW�O�t��v�����6e����荨Nr!C��Q{���fm`*\U���vr�"�ϹnnX��<�c1b�J�T����� p�u����[�
 �=�c�3M�@��UɅ�]�B�3���Zq��ܖ�k�֧�(g�#u6���p�JY�-CK�LP��Z��w{o.�:�ڂ҅b���'-�ߡ1�נ�VX]qi�n�0� �1ǳ��p6�;{.��Г��1.��)�1f`U �-+e|C?W������,�� m�P���]��h+4��Q��eYi'"������Y�g�X�9��e����֨|��T錦i Zd��n�8���D��+���cZ p��J\P���s��#Tb��3̓�?�C{�<�Y�����]F���A������CZ��G�d�����MDh]'�P?�QyA�[��^R5Y���Tk�H�s�clsC�LD?H�Ѧ-x޷�Y�㪢3�3S�VHL��s�)�/�L��)Z�%Ηz����VE�9PP��؟�%��$D��i�i��S��^�!Vu���D��x��.+����x�b5ښ9)/��� Oq	��-#�* ��x#>���(kb+�2�U�Y��6�V�V�%xA�N:n'N86:F��_��E��� Rgi~F��ֱJ[���su6�a3�mR(�5�O*��/C���;�4f�.����������,�ό�}ПQYa=>�� �a���cn'�\�ISZ����{<��|��֖��ݠ��:���(��-��.B��C�7Y���{K"�l���|��ݲRiei�|��Ŵeni�u�դ�����L_�~V�Bo����	�tb����xE����"�@���;X�Z�N��5i�v��̂]��Tm��ާ��^� �G��q/'GM�j�,;:�|��s�����^��q&5�!�kyGH�Ϡ|�=P��GS�N7U���e�(���MV�is����%����%]�g Q(���^r�E��
�)���V  ���1��p��n\��ڶMt�0i�����c�cԖ���w�#6�w��Y}9����҃X�c׊Ԯ�$�DE0��-߶�Ն�YY�S��^��D��e�s ����=bi;P;�;B�B��L�rb эl��L�q��E*�o��VDF*���T������=��S9z�\O]8�R�z*���,�f0���;�� M��&M�*�R�[4l1)'@�ρ������yG�c�M���� ��'9����:k�V4�f�Vw�|rF�Mg֧��7�3k��o�V�g3]�vz�3�q�v\�&_��k2oz�:NH5�wq��P�{V�ޔ�z���ߔ����LE0�	d�6nsͥ�C�Mhm�O���j����`������`KzBb	��w�2���<��T:i�R�����J���;vcu�ݨ{]YX���QD�GWXT�=I�����2^d�؊'9�yx*�<,N汝r��0Ibu�$��A�X���[iq7)C���Շ}O;�'eC�Sڳ����h����4g*j����k�ȐC�w�[�����o�������'2[q,���}S"��?�8�ŀ��;4f�,��юo!��f̲|�FZ�a;|Y�������W�>/z5�|��B��]��kڱ���u�WC-0���^FGTM QW��n|炸�M�slK�ۃK�I,��_�d�Ulkv\);�C��M,�?j1O8q�g�ы/(�K��?P�"R��=�OC�R�?a2�j�ޙ��:_�駏@��e����ʐ�G�OX��o�����X*�Y�t��9�[c�?�[U��GN���ʊ�ч���Z��.�A*1(|d?zS������q��g>gԯ搿C�ˀHJ=���{ <�N �7/�R�8������R|<ZY�Z8V�=�͸X�1�O_�{+�F�4098R/�A�ޞ�y�m�
<M���zJ�	���o�h���/�������hƳ������v�_�+gW$ήH|�^ca����� �� �i硄�bQ��;�H�,�'9�eb�T�K��yҟ�wF!F��~C����!i�2�q㝋�B��/�.ЂR�Q n_�+-�����Q/ Ϥ-W��o�~�Y���3R�D>�O�����1W�a�� 9�,}cY�W�_��
��>���<��NC	|||j(�~-e�Ms���8���^�����C�<Tb�M�<Dj�"�A��i<Gq��[��૷n��T��N���d0�Wc�]�-�����9q���I7���Х��=���_|n&��$p�n$RdG�kl3�s��![����R�d��uXZ$&��R����~���������C�����:�/��1� <�k��b�P�{�fܬ�B�C>���&Hgn�yd;r�^�Y��%���Vl���сP�9����\���o嬸��$(��S��#/㈪�k��-1����+�3�:y!(e���Dq�*K6+��$]w_/�0�_��[�N]��T�x�`�E���Z�t���T������o��0`}�9.*�vU���9�T�+���S⾲������e?I�Ø^QI��C�XX�X*�(��/�q*�����}�dOL�-{�9��!��m�C�v�VmZ���
Vc�~�&-��֬S��|���� O߉�H�ʡ��$���;�^[��w��?:����q)���=x(Ab�eV+�f��:�Q�u��(���h��̜sz�����r��; s�>+�Ig���뱌�W�N�����+�kA�>���rX�Q���������H���c��z�*��Cr�j��]s���f�2<,� G��հĻ����H�ȝ�a!c�J��0�ɇ�h�����J�{��|��%${�?Ǝ�P���f*<�c���ٟ�����ɂ����+x�i��QK��t���&�S���<#^�&�F{�P{��=0�$�o�>�)R�	�Sӎ�a��)��� ��
v*�)�!x�i����28������Y��.��RXY�I+ݗ��< 2}����l?����ө�q�ٮ�Q'9G�Z)�B <&� e7&pIAN�}�CГ�T���*�Z����y#X��,q���<6����"YJ�Cw�#�q�rڨ
1A�Cw��9�v������u�l�ű UR7�s��Km��'������h#nj�6�C�U�U���Di� >q`%T����6�Z�یN�f����b/�7HSI3&�cb�F�VdP�k��`X��?"��ߧ������a_�z�o��FM߂+�^I�3�,�yGUM�Jb>r���&��HU?Q��)��/�
�%7�+�I�v(��(��`���#��e�~p��Mκ���WVr��k�W����0�'��ن�XO�����+=�HT�N��#A-�0CԄ�oj��.y�~'�"�%nc-;TͼM�I�s '�}Y��ם��(���rЏ0�w|Fʋ�f�%\�V3���!k������74���'Y�Bj<�o����4��[�nӑzO����^;5RxLg�GF�ʓ��SQܿ�F^�� uzi������V9��7��9���$&Ӻ�/l�?��<z��iR�Cԅs3����<����'Q�tO��?6�����ݽ%��j'��;��a�}�SY��z�a�+k��G�D�T$��6j�>_YP�IE�Y�isސ,�$a�<�:�|�/&_h@+8�/�3g��'
h��*�U���;�����5ipfkF���$��#(?x���I!�O�(��#��~V/
��l�:I�brd�d����J�y^(����	ӓ��N"��^�"5mF�0v�땦1ܩ�4�Hy�9yT%Ψ�z�lN𑆃��U��L�r��kGUvT}��6�p2r-0�ZJ�<5�y��1|Yi?@ԍ��(��T.0u�/-����Kd;O"�z�Sq���캰%���}��-y���l׻[(���F��JfH���?ǿc���K�Ȇ�A��*�S��&�<N~z-sm8%�
������S��#Fg�?��RU{l�M��2牖R��QV�Qǐ}��u�W�+�K��/�+%�3��yp��ٕ�:�g��@���B��(xiS>�G�nS�x���d�}d�4Y~��_��#H�Vx��װ`���fq�!��<:�� o�|>ܶ�)��j'	ӯp	�6p= �a9�b��5+�x�\{�3 �c��QE��?�
�B��������91�7�x�;�t%�����/1(q#������	A!�����^\�DC�P;|��l�H�u 
��4v�my`(�m>b@��v9�o;=�\�<�yy�4K��,D��g`�� Q��ldX"��)��u}-�RgcW���36�k�3y��ֱ��t,��rq�y���N�D��|���1i�T��Y�N�[�zsKgj1���lY�9���_b�߳q�tp7��t�4Mٱ��&��l��N���8�Η�ӆXjp���*���m��Aɦ�3���qF?���?"��4H4�%�`3�C"��GGF!f��� `0�uZ���<�++���
( �8ē��K��L�^ I�R��0��'n~�e�`fC:G���QK��c��z}�ـ�(���$N_a�}����b�t���qׇF���1��k�F/�̛�!@�c�A��RX�3ɕ�~NkQ�=��u3�GCE�,)�{����O,�����VsiE�in�P����.�*�� �N�1�TX��s�� rtt�hyad����VM-۬��-�TT�ei�[��XVx)�l���Ṵ�)�9��9�;�p�v���������s�s��s���=xu�����]z-J��cxw^�'��W? �y{%����[��i�`��w{�k&<�Q��`�>0��ja���ǡ�����G͐p������ꅭ��9����I��	��ۯ65jE�hE�! tw�OZT+�n�!��)��a<�o`Ί�^��o,?��ᢗO	����E�P�<�{Η*`c�	P���"j˄|��UU�Ǫ��9��9zI�E���ܟv�S� �op���[��u8��Q�����}��!����u聧
�k�1)ĸJ{� ���%�F�d�������ž�?<S}�`�e�O�~�V��b��G�	_Jb|�F�����_�Vyf��g\C�A;���^�U������3�b��=PS�+�+�*\���Q��6X�l��PT��J�F�;A;���&F�=��lYC��^V�0˖5C�����v�}-͝��^@ƯG=��p�D�<i��-ێŹm��ċ�s�,�htŎ���$t��
B�9G:x�Ol���D�뜍��R_�1�������D��L��B[BAŊY�=�B�.�}�.�c�*_oV��8ј*�w���B/8�#�$�{{����	���^��_b�{f��'�-�N���0�,5�ZN�o)�3�q޻}K�q�kAu��]Q���vZ~��kP�n�b����a�����2ENP|= ���a8L�-�a�X��l"X�-�rz_��=fv�j�U�)1t�^x��'|K1��&��봫�'��!P۾�F�����E��x�1���~/0���hI;�3�7N�~����8ݓ�.Ce�4�Z�g���F����2���v.u�h�'q���L�F�.�A#X�Yطg&�ʐ�ڛ�ޱ�%�9:3�5�n�-�8�]��n'�
/?������V8�=�z`�U�sջ�y�4��୆��	��ۆ��G��+NC䱺�X�E�2����ｖ��{��|`�c���'3��u��f$�%4��a��ڙ�zh��Zm�_伺6�U�~W�r|yƅ��M"�X�i��&�=�t����c��sW�@<��7ל͈�v#�;���L+2�j��M��1�v�@~�����]�*�Ӆ���&1��K����sx	�9�������?r�K<��%����n�Lf�\ܲ�Yu������e¶�r��|�΂��;��.��\��S�?G��ѣ[�j$�k���N���z��ڟ��:�!NA�����ϗ�z�k�`��{NQ-�/�cb��_�^��Rzq���������8� ~#0_�'o�|鱯#SEД��?0�@~`�%�}*�v��}�fq�F��O�p�(:��n՟�/fׂ�ܛ��t���%|��n%_֏��ڃ7id�s��h����Q�-�y8E;�R;#�N	�4=8��W0����$��e�^��:7-R�qo�4���)��}�K�8�A:Gu���78�2�(�������h����o"}�5-!J~��)_NX����y��M��(F�o���E�(�����O���2p����|�`+l�%��~��s���z��`����#�ຜ�X�� �,��'g[�?!�w|}�?3C�����9�%���Apc������:�T�11����s�?
<ҳ�U�Q#�/��5��55�
#Q��N�x�l�^�8{��x0k'�t�ė�e���*?0��)}zTY4��^�,Q��Y�K��>�SX����b��k��
C/���,�6&ҳA�y��2~�^s���.k�/6�'5B/�;����g��XP�7��kqcFC[v~��r��eֶ=����:9��弇�����waPB{�6Ä��������Mر�������N߷���h���m,;��sRy8H�iK;���cx����u�5Cq���6�[��+#�t�3p7�@3{�Z�)�j�"�����v���{�Gq�Ow�<�@/��iO��u{ho�m^���$ҏ�:p�3�U<ɷy,�����ћ�?:�����]���㿕#�B�'�2|@DyZ������w&*�+�n�������7*"[8S�X���{���#��x\K����
��I�j�W���.f�o���i#��B Ƚ���O�nz�r,�T98�,��m����}��n��_�d��j6��U����2����;c�Ҷ��D��⿶�ob@�⿶obP׮N��9ơ[9akXt�G8E����?7�}����(v���L�)���� Y}^��7��6�P����|�l���{���&��x�� ��D�� H"�R�}d�0_��P_��ڴ�?�H�g춏�m!���ƍ��6�?�uZ�0<�����C�R�~�	ӕ�ue+Ɨ�	����q6y�����0zh8���'B/1Z�"Qy���K�Tm?A��k��Mg���>�]���-���3�3ҽ7Yp�5��Gl�������`=�F����:�
��P�߈�@70��x�"��c��?_6˝��72㴃�.�dƽ2(�u�!=�ݍZ�)���0�Vd�<� &�3�c�L�3�aޫg��6�Z�E��2�ӝ:�͸I��]��7��L�~�	j�W�𠞈�T��04��a�u��ܹ�@�K���!��]�N�kx$j7]*�z���|U�ӯzG�$�i�7#�Go+��Aw&yO���p�6���{Y�����n��%�zEKxE��(�`~�4�)�%;��N�i�\P>�ۚC�
��eG�y���y�c�j��ۀ���}�F~�5�_Q�W�Y��D��m�s�t�XK*��'n暋j�&\�z'f��̎ΐ��@-��D��32]��#p�w��}uG <�vtF.}�!�����F6Go�T��Qy��d�m{�=����\�"�Fxc�
oĂD��A��5�謑Z����-���jV�X��gЛ���?�f��/��#m	��{m��<�\ko��{Fx�����r�<S2mei�ܵ{��߷|�����}��g{�R�,}K�<ǽoYʕ��/`{��o���}K�����<�o@8��������o��%�?Z�$>��x�ry}�����>߷\�M���� '����-�����-)��}K�v2� 3`*� Pp����-�8Z�7 � ����-{�7(��xp�X�<��V~DȌ�"P��2���&6����̉S|�)�[�.a����F"���E�w�K���ǖ�q/	�"�3��	��L?=�0����r_�+�Y	Q��d�+⽖�G����Ox�,�GnE���)~#�����ŕ����Q�)Q��Bo$�N��%�h�m /�7�k�֦
j�E�N6O�6c>��o�' ���/�}Pk�~07�&'�z<~���.;nI�q[���^��&�,���oI��G�.�%��}��Q�;Av��0Qx�L�"^h�|���e���r㸕郋n����8F���{�z�߷cdc�~�°������	ށ�1�dAmz�Oy�n?��H�X�!��?�)���K�	����t��^����Vw�{�+Ғ�F" d�5��`��g�����+����(�@�=[��am�鶈���3N3�����I<���Mn�=6�Y,�:��77���2��^.�1���Ũ����;�^�1��n��-�П_46�y2�o�?�]�+���=����=¶�f���ݙ�u@J��b��ۑO�f��;k�v��+�X���kt�[0dtbB��Vv�N��:�1m��(����X�/��vχ��じ���c1�����W�pBoYo��E'�(4ć��`.c.���@�� ����������+B�^/��/?�#���μ�B�d�ǵ�|G'���#>��i4�@��K��!.�,l��@d�茬kz�,q===D#�[4�qo��My��B|�\��>��B���Ql3Elc�*Ʊ�PT���R�>O�v-�?Rq�%l-�b*Ƴ�T԰����u<�&�˓ٙT+�ͣb&;��Ylͬ��9���S��T���J��*�ءT,f�����GE7{q%�{���I*.`�^ɱ@_b[P�5܆ɾG����*��%��Jq~��H����Z*��?�ǩϔ�>*�Ci�n@��J��v��Ι�Y+;��s�t���R�xY��L?+�����j��N�P)�Qe�����*�Z�=�0Jq7+{�JY�~I�'h�����G��4�Tz���J;h����?��Jq�}�JqG4�R��f��Y��l�Cp��Ρ�X�N��8�N��x�fP��z*�w+Y	�&�t��B�p*��4�J(P)}���C(����I*MF�T���*�D�{�,㛼�[����-T�3&��T��٧�t:J���.�D�f�-v�4_?}$]C����!z
I����:NG��,�uR8�>r%�3��+��U7pK$ףNW��k���(}��wwv�$�G�y��8�X}$���t����N#���\������U�Ο9�}d���t4��ռN%�c�G��u�p:���:^'��I�Gn�uR9�L}d=�#�:�Yz�F>�7�	=w;=Vº���lam
U���I�C��PV�Ăh��)�j��Ԇ��97����>;���k�l�E���>�q_#۟Q�o�E�H���R�|�,�5K�g�R�Y���Z�`2��0�W�v4�&�-���~�xQ&t`��f�};�6g���V�L�v�X��lXJ���{�������z�h�Ay��A��YX�m�(	��v�},70r���y���=n^K7�]�^u�
+�0�@|J2�LrZ3�]V��:���f�~�?�C9�-��7��\����9���;.��N����峻q.�Tù�⹢b	�Z�{
���O�<�2�����}~ǐ�.O���euZc������'M�V��-�Q�m�pۢ�7wz������Z,���sn�������^��F���E�g��i������̐Y܏)�T�ytD�u{6N;v�G����?���t=�"Y	��M؛�^�Kg?�!"�����.���N�y��{�.���(�?f�� ����ǎ��	m� Ё��ư�Q��a��	e'!���t�2z>?% tjE���D�G,�l���L6=��5啻_#�[}�?s��\V�	�}���r~x�׺= �	�ݺVȶ�¼��{u��U�]��	?����:>�o�o�n�v����R��qhx��~�
w���<v��ԃN�`�����m���UE/|b/�ӎ�+ٓ��?޽���Eੲvtw��M��\�n|����^�P+������c�|�� �н~���cDt,b	����~��Xn)��VO�&�����*�V[jx����*f,��� -B�/v�����7�8ث�	������p�B{S��==襷��3��PP'�|��9��V�N{��4�����Q�|��;���2;�9��
�נ}Q�����v3[��߄p�@'t��:�w�D4j��V�ۛG���HD��䘧�)���:C�@���� P&f\�{l�	x����� d 0PXxP�88��¡��
`�6���
��	�� ��� ���{�(@� p/�A@��n�G�����!l�	 	`,�( ��pq�%��(��!̀�z���Z"�<����$��ǉ(���"*�������D"ГQ��Dd����x��~2�Ek�}����(���M����vT؝��+C&�z����dH��1��!�~��1����'�#��3�ZnS�p�),-)��V��3�Q�v�q�KK�6�u���2eť�ǤYx?��2Ɛc3��bg�k�_du8�n���'����\5~S�7e�������]�y��^���=בӍ¤�1O$����c����\�-V`�.��1��p�Gx��7�#.�3�"�$�1�x�~S�����{(�+)!n0��q�g%�ᇦ��o3�;x�NR	4ѝ��H>wH�4cB�4m��r�m��}?f���@��6y�= ����J����B��q���A����l�Mlu:K!]����38w�7ڄ�#|��M��������:� �@DD"��~�"Azzz$~J	1S�b�yj!QK$�����XH�|Aq|�T�+��ҟ�B,B�J�Z�I�p0fOi����@<��BRJc�NF�t�=p�vИӘ�P{b�� 2��9$�L���t�ÙZ WO���iBH��&)�Fo��M!*"!r���`/8�T�\���7bഌ�M}���F��(�j�BS2+�/�Tf��"�^��\d�\`C^N)i����X������+�����J����o^J���o)���4�\pG��xJ�j	�Q5ڜt9�1\ȝ����Bv�(�V����Y�ρx�����A˘���u��i�a.(��)4>��Ɣ�򈹧��������2��n4��4���3�]�����Eck�U>��m!��u'�\h)ř���hw�?��z��=$�S�N�.�N.�Ki�ay���{8$������B`��^F4��4Eg�x�X�8@�z�WQ���7�����7�T���Km���N��4��n9���+/��[�	�� � =ſ��,J�N*(�c�ũ0��ؓ)�^2�K�7;�1W�Kys��in�n�|�� �Bʙ-$�\�������𵜃�8�j���,�'�t��F���S��C��R�i=ZL�1�ػ䆞�Q�>��?���AL��f��'	I�_N�
�瀍 Ų�WR_�4�J��A�.ŴurSU���غ�~8'W����UD"��l{��բ�"v��@�A�w�h0�x�b�^"���T���6�u V����&��7/�{��F� bg�n"�	Ħ]DT�+A\� :A��o�5���i���v�_[���B*	?1�\��U�f���TҰ��a4��� �)ϡ�J���s����؜�M|�t�!��D�Di��P�s���B���~/�mC��w�)�_K~��-y���p�ex�v-v&���R��y
v��.��ȧ�� ���C�x酐�?"8D�2D�H��!�GC�xF@�j���Wq��vVqj)b�x��0�g��a�m��i-+g:�����R�f/+�8ܼ1����yK)���zA�b+#N$�J���N8�e�)
�L��	1�k��n#%V�u��ʁ1 RXꮄ�2��8��v�g�����{Iz�J��X�2vC�m�N[0�stvp,�:��;M���_�R��K2�=>Bx����=��Zh/��0x��!.t��y=v�Nw�ӂ��CI�,s��tP�|��G	���E�u��ޅ�NB]�zJN��g�����5���.�G���3�{Oנ�^��KZ���\�e�(*��{ɇ���ϥ�ϥ[D���E9�L!>_ڋ�^'�GT��߇{��.� ��У���(ߥE<���|ʢ^Q�|����[���LF2�c wF�@;�έ ��"@�턌����4@��mp��N��@�r�	�;�!�n..�O̧7�{# �@2�#���4?��Y��.(�s\v�==�B�݌G� �n��@u�Ӄ��n��e��5�)v��e��ӎۊڜ�6{�DL["_m��CD������,� * N�`LL� ̀,@& �P $�Q�D@@��b"@@ ��A"� ��N�����(�p�8h�4v �� u�Հ� P�( �����X	` f� ���Z ̀��*�2@`:� ��h> � S
�p�p�A\	X �Hd�L�=��>Ϊ�g���\�w�T�?B��P�1��~I6Sx1���������D蹔wӛ��7t, ��1}@/��t�t��:��씻�9���r�y�l�'+��Rd��l:��M�#���o�� _~<����S��w�߀��9Q��:m����gP�3h�,D/���]t�!���B��t�tc�����4,���t��EZ]I���f|�����QR	��c������!�S ivhBf�i�N,-�O����4S�s�e����Ҙ�uфLq{4���|�g{�b��X]T
� }��4��A�i�{t�n��
M��JidxT�S����z�v���+r��,��E5,^^�2�ݡ}��vМ�s����U��`���j��U������K�,���DRe��oӘ�H�6�q��8�jY�"����Ba�
�{���e�:���o��e+�oa��k��-�{��x7A���,��S
G��\������Ȑl������$RG
���P&r!�$�+���/���Ӭ�/��.��������_�/����?�����v��/�z�i�:������_��_�����/~��P�_d>�]տ4��pwסW�����W�,Y����}�W<���G����b����??�t��u�7<��s�Ͽ��ƿ���M�_~e˫�m������7�jhܱs�ۻ�4�}��}��A��}��ᖏ?���g��g��_|y����a�o;�����O}����9s��܏�/�t�O��#����00j��Ѣ����zmܰ���_Í�n�%aĭ�%�~��Qw�#���
�J�����))�::�Es�s�9K\���y�o����{�>c欂���`������o����?eljZzƸ����ʞ8�<y�%'7/괻�����E�_���L�#�[��W��<����r�B���r�]�
�����E�;M�����Pu.ht1�u�7>C�ſ�m�����󴅈_��{Q7uß�Ys�����҃i~&vS��N�vSw7�wS+B՟���[�-o�y��j�ۯt�O4���m�1ד��1�/�2pi،�z�X�yK�����i�7����7���~�&G�fa��5��?�ͼu�W���<��`����k���v|�� U���$�?߽Q��v9��ͫr�e�+ȿ���G�晿���	�Y"��/
m�*��:���	p4�/�l�w8��@w�`Fz1#_i�[��!�B>�b����	��Zys�ы_��f὘-��nW�B��G�v}�5^us����_���o�nB?�yY7�z�3|���,PO�&�}���&��M���������=����eA��7]�{���c����h�T
�k��X��#�'��-�w��\4��i� ��	��JȻ��x!����-���r���O��n?��# v��r��ٸ�pf񽘝�Qr�D1�bh<"b�>��~'��Ǻ�]�a+g��c=�[�n(_��������8�ڷ����1m�y�P��m?Ǝ�0
�st����m�0���F�����vC��=�g|���P���������Cx�]�o�zЮ�v��%�M�pn,��h �k@,h�ߦ^�>n.��}�PO�y�	�;��^o�/�W��6���t3�5�o�K��c/M��K�/��j���|����OL�4�k,�v���yC7��y�v���3w�XQL��x�q�w��H���/����-�ry~׷=�|(?[����p���}���Q.CDӘ���I0��7�8�9���U'�yی��`�������� OC�(�]4�pa����GD'���?]����w/w��/�����o�&������\����]�}�/m~�ӗ���k/���y��6��?rQ#�3!zA. �5�A��p~���r6��gD$�4�c�2��2��*�CY�\WpC!I�3�S�^AH��.���9�dRVzJn� �#�Xe`�s�I��b�T8/�:-�BN_�e���{迃k$�6��ԁ��qp��La���������k��%�i���� �v��z=��ɡ{Z��YJuKKJ�.[��eO!�R7�f�A��S�pAtt�Xo��<(�u������#�,v�o��ei���9s���^D� �xʥ�;���f#"�!����Nb"�6{j�ՓS��u2����������$��8D��FH~X��[V�4�z���՗����).���p��z����� �=�J1��4��Ebô�06N����w�B���a�n\��'/,N��M���5���Cc<u�u����'dXX�1�ؠ�a���-�����坻��PչOl7�h&�bR\̳�ƻ
=t	!e��|�j�g��{4�p凐��*�$�V�kz�B�5=Nw�;<�.$b�{:���'_���"&{�J��C�ɠ��(���(���(�ǧAcϼ
����}ec/�q e4U@FQ�-��'p9��9�dNDg�)d<R�1��ő<�:!��<�1�I1�S0W���I��( �R�aK�bm�c'(S�\�%Ed�Z�t��X=�����a�6�L!���2>g��0�0���;#�R�!PT�w�O�����߂�	Q������ȣ�̜�PG��@]:��X�[A�z-X q%��0�!�C}��=��S� � 3��l��@�� ��Nq�����1`�Nh��/7�m�u砾| �HH�}����A�Yh��	�9�g �E �����p̏c�0��$ =,����z��$�H$�'z�Ud }�A�jmFK����ZG�AЯ#��zr�<F�|�k�u����³e���Y�g�f�ٲY��e���g�YR�n����B�,�=eO��~;�s�f�d��7%ʝ���Y�䷦i�ݥ�n�X.�M闺�ߔ`����h��2�oJ�O�_G�#��2e�Xs�f��_!d���]��2�� �!�^�٩��CVvy��/Y�� {y2� ]�P�d�#���r��q��,��]���E�|9��N�I6���\\�,d���fd��	�,7���-y�p٥���]� ]����^���_�Nn^otRJ�l�m�� ���%'w1�<�Ջ�8�u�l�t��K��&�@u��p^Ww�� ��"�.��e
���s���8���fnw�a��Z5�c��J� _!�<쭴���_1,��^VxkO}}�<�|W���&���}�����2�o~۠����������>^ (���{[�,0>ρ�'�E�x޳?�֥��x/�����ݢ���zx�x0Կ��W��^�ʫͼ�)����y��x���~	!t�4��3���~��*��żx?o^͛��t�IE�i�)^���g��s��V���y�üy\..qF�gwkk��)~������>Q�g.�����x9��w;r�}�����[~�����?��˰p��d.�����x�g�ɉk����O�ҷ��UQ��7��d����/rb2/�����k`��uG�'_�c���7�Ek�l24<�?������d�'�������!�E�K\Ƕb��D��	�P� ���,, �ŀ逩�������� H � 	�8� ��@G��� �� ��M�5�����>�2PW* n@1� 0�	� � �~��C�}�]��-����5�U����0�H��+ ��8� p�#"j��l�� Ώ���r������R���=�y������.�>���g��B~Biv��.�d4���禑?���o:��2�o`��>����Y�}M�{	����O��e."9-�!�-}K���M�E����<\�_q��6�E�b�R��O�zJ��Qh>�ܫ}@�V�Yۨݯ�\{J���ݤ��Rt�uV��t�u����6�u_��y�b��p�!�0��������fr��:SB�⤇��MږDh�o� i�|+���������ʋ���ՊɊ|E������&�H9Ly�R�LSNU(����O+�Q��<�\��Q�_]��P���kR5�5��wjS�y�w��-��:�Φ{�s������W2�7l1�2�c��m�߸Ɉ�	!x�Tb�̕��<)�*�N"�.�����"{@���,V~��y�|�\"�&�O�g�y�|�|�|�|�|��A>@!R�*���+��� v�)�+>S�Wj���Le�Ҭ́MW>�ܨܤܢܦ�]5F�PTY�<�t�[��۪*�z�_���b�ݚ�4wh�Z��nm�v��U����V���ݨ����[����t/�u�����Iz�~�>�d�Ag�b�7���L�dB��$wJ�$S$J��Q��+H�3�1�B�CZ*���&= =.5��ʌr��#_,��p)�9ʻiZ8�e��J���!�c�5�����(��ܣlV~��T����2R5@5\u�j�j�*E���U߭�����UW��P���A��]��͚��/4)ڣZ���z}����M�C��L��&)�$�	�>�(�>�v�4K�'}^�I��t��K�)�Y�p�M2�l�,G6C断��%�3��.���H�Ê���+W(��Q�ʪ�Y���E}Q=SS�Y��H��c�1U�֚H!�4�b�:ٳ�d��,{M���M�~�Y�O�� f�����?� �u����u���gQ�Q���B�W����r�^PmV��ڥ
S_�NV[�T����J}R�#�a�&Sc�ܯ�i^ּ�٥9�!�~�h�P�F���&�A��ǵ���C ݕ�d��:��R�Z�J����'�@�~�ެ?�'�k#NC����[o���3f�W�_��F�~����OJ�B��,�V�T<�~W���U}V{B��ί����Ջ��������x�$�=z+�
�"�2����_�GFr��������@��n\e\cd�Ƌ��$6�jeқƛ,�i�R�#��7՚6=nZc�`zѴɴ��hz�t�t����s�7���MgM���nN�#iL�:ɐ��4>ɜ4+ɖ47�,�Ѥ?&mNz�w!���0I���$I��n(�;!���@���6�T�.�> ]-]/-�3�����W���������O*^��۬�P1O���I�s��T[U;U'T�UC�7�Gir4�5hӬ�4j��Z��a�Q�)� }�ަ_���Pi���!�x�q��ܸ��W��q�2�
�Ӧ���C��J�4��$��q�=[Z&���]P�>�~%&K�����M��d�do�N�����W�?�g)�A�}B�W�@.S(J��e�G�O(렎�%P���]��.Pߢ��٫�RsZs�vԌo������b��Ʒ�{�j�R�ʴ�4�suҟ��%���y�7I�a���$z�Wr�d�d�d���:I�t�Tq���h]>���]&�J-&�Qv�l�L++˖M��#�C�|Q��쟲���"E�����2B%TE�D*-�����2�r�J�*�j�U�긪b�CuA5[]�^�~X�J�Z�F�w�7�a�&A����@M����T�\�R�J�ZsAcՖh�����\�{N�Q��n'�{��h~�a�@m����k�~"=!1��eB��-�����m�햵Ȏ����+�V��@M�W�/�?S�Ƞ�^�yCs\s=��T�8m���Bv$���B���I3�S�ӥR��Xꔺ���Bj��/n#��E�E�Xy�<^.��A��%�ɋ�u���321��t�p� 0Fc����(��h0�A�΁�f3:��Qc2��Mi&�̕krJ�ⴢCqAA��P�}�2N�+����$��4����QJ���[�(+��Ư�|�\�R�J���:�e}g;�]٠ܥlR�V���ҶUyT�*O(�!�;��D%�S:V��W�U	�D�(��?��ɪ4h'�TfU�j*��*��X�h%[A��Gί&J���!� 3�rB>
�zU��YuHբj�|$TG����B�Qg���f�T�[]����U��^ݠnVRU��N]P4�4�%kҠ�6k���ާ9�iѴB���i��4�Y;U��.�n�n���m�u
�A��+�U��蚠�>-\�>N�ѧAmQ���:t�~�~��N�E߬?��8��0��*��-�C�Qc�j�0Vk�N����!c+ԭqP�&�4�n*0�ܦ
�Uk�$o3�2�B�)H&%$%&e&'�$-K�OjJb�H;7w)�$J2%�_#����K4��}�zI�����q�MЗq��tM�}��!}p٪?�g�'������hu�!� 2����!��he��!ِf�4d��S�j�n(0���J�U�R-3,7�4���1�6���ǶͰ��`�eh2�34C9h���
e�����J1
�B("(qP2�P6�ˌ����m�&�	h�.�I`����5ř�i�%B{$�x�A�9!�{U+M� ט�]�7m��i�h���wܯ|W�+ߕ��w��]��|W���PK
    +Q�H5ߨjE�   R    com/smaxe/uv/na/lib/jitsia64.dll   R     E�      �y|SU�8~�$4t��@e��Z�Jul`.M�F)�X��8�b�T��43�h��q�eF�}���������/�q��Ā�R��}��ܤi����}�����Cs�=�,�y�s��<�����Y�$��$5J�G���z�oИ�����8���q���w-s.�������qV�v��i������^�w�,�=��~�e��Y.����Lv�se�����ڧ.�kƔ�S�t�9�N���7�^��L��9u"�?1�K�mF�t�᮪�X߹`��I��?�J����>��%�ufgdIR;<</�r��c���d�gH��ޫ��$�H�=�d����gq��$��%i�x�T� ����`�j2�̀���AI���.��X����V 컥o�$-����۴�$�g��N�f���7��_&�IuWc�a(\/0���t�R���Xc�k��<�U߱�*I�1�8��5pF�)�
���s�Sc��p���/^#�F�l7��CNx�_�����c��^w��4��v�
�kS�<W���\в]�D���@4�rB�*3b��7pl+��0�/���S�K\v5��
�e?;�g=*���KRI����S�η�F�!�]sy�QԁG�*������J�@��.����̙{�Z{h=�ˬ��$�d�
��@40���xI���*�!X��LzEi�I�j�z���7��ōЫg\�T�)}εn�?���������j�7 CU#Mr�;&��@,�zd�Yo��S�nE��̈́=��O�wF!�T� ��L_σGH �*�f#����͇�@�ʇCb]�YK�p�m~~X��t����`�8>XXk�:�)ܩC��1��v����'vSV�U���EiY�ҳ�����ݔȘp@e>	{U��zEA����P�Y�������3
�H�f���\6o�|���g�y�XD�@6�
�h��H� x]?;�ݪ��_�T��H8�>�u.��:1? si�mQc�f�M+Pc9��X��}���_�z/=!(g�f~��}�
�1����]N~�)D�1�̠&�Be�PLP�]��l�������H�n�ߗb=�Či��N�:�ن�K|BL���&����:���J�S��u�GT�= ��v]e=%M��蛿6�Q��Q��j�ʎ�G?�����?q�$�� C��N��8o��n�!$l7��caqyY������V'��ϸ�'4�Z���WV¨@7�y-����le \	��KR�S��g{�� ��8��dL�O	�s`"�^���{'�ݍP��A�T����H�-�fR�w��]}s����9:S9���BZ�5)��f�`-"��dg*��H��4���alw��p؜0V���B�@6�t�>��p�} �Q�fnG��R���[�F3X���B@ߌ�� �����x�6�j�q�k̹b�ʐ��)�6C�sD�Om7��Mo��	2j��4>��Ms	��|�1]Gp+ܗ�
2X0/\�6�ȵ�lw�����:d�j*��[�? �'��Ќ�vN�*k�ip�u#	�l�K�.������u�6��S��n
�a*{$���DC�o�,��m�ax���4t�n��xb��Pd��N;���DF�^�����*�iD��G��ƫl�]���rTh������'��N!�����_w��w�M�!C�P
?��$�Q��*��cH���"dI�f ���c�OnE�t<L�2�dq�S.�I!j�����ȹ۵+l�1Q�6�A�u� �&սiY������1�`5����X I��8GM��T���P�LP{s��68�u�[#Td�`GS��#tf"�n#\d.ڦ�T����YS,��"�����������ԗsF}L�*�ߌ���x��B�o)�(J��`���o��ew?G���V,v ���̱��e��8��pNa��k��j��ޥ����>D�v�;G�LJ�U���렩�с|�m��uW#)1��IhZ�z��c��#�U�CU��k�)&�,U���#�5(���m����Q�ݛ����1Zs����Q����lH�?��
�9Qm�D�.F~Ij�H�t��jr`��<I2&��;�ɲQ���ng(���5
��+��V��NEr!	�1���r��O{��7���3ݎ��.G���r'b�x+�;`)��#�
��+���ֆu!��ŀ�X��d��ą0�A��˶�	"�a���$a� ҰnQA |��udb2�-�$�o�<�C��8���^2�dK|�i({����i��L|�p�-W��j��-*���6��mg֬�%�����W}��|�������������_}��}�����F�����i̚�J������t��#��{$����ɬ����J�`߇�H��5�@��g�ܒ����?W��6�&��G���{]�'�7����,����~4�	�X��#yfܦP���[�i)+�ޘ��2l���E��{��C�AWB:~��O,��5���_��0y}�ڷ>�Y�$s��Xm�ſ�0�=8WAR�W
Q�Z�#6*��T<��	0�D�۩�7�a�`�&��B�`��>�l0��[yKy�h0b#�+�6OBTS�	�Pz��P� ,�n�nO�5�`L���t�S%���M�K�����/V/�R��܃Ԛ���{��/�YL8y�o�'ڛ,ڻZ���=T��H�U��4�YZ��[�F3�X��^���p	���+�h�5�Ŧ@5�Z0m}:Eȯ�6�?{���c.���OU��)þ�
�~U��@��8PvG)�v�����Az���z�E
�Є���c�$0�?��|�%Ip/�1���`-��85Ƶ�p=���-T-�;(u`��P�ZK/y��)�H��g(��X�����#�H Eom�p��E���
�̔Ҳ��P&S�,�����t���W�¦���[�/�(�u*^n�epe�V ���7MNX_s��Jf઀���x��"d�j6DZ-�=��.�i<%j���4�F} ?���-�+T�R��gi\Ao� �l�=��ش|H�?�[�f���qh���U�H�*O�� ��.�H��U�ʭʼ�;��'��������+���F��iF�br�u��P�{
p�w��E�ŭFAө�A?���{&�;�&z��E��;}K�ؚS8���H��!$�_~�'TAc�f]��b>�<�;e1��"�/Hs"'�P���6k.v���S�C�o$M y�S
����A�D����P_�Q���O���jQ�>fZ���s �����&5:����B9\AA�(�$lf!������o ���&�N��s�0t��� ѵll��?��K�Z���( -,Z�t9`��x9(/��W�FS�@HuߙS́����V�����E&y��FҌ�$�Rxu�D	�u����R$T�T���<"��J(	ũ�B)�;j�@O�d�E0���w)v��6����`C�[`}5�*�=^<���3�vH�=TC�+NB26�	�>�w%��������KF���Oi��1?�|�h�qҬ��wF�R��������'���~!q�`!�`�e��c���SdIL8�+�+��y�2��g�0-R����Y��_~�iW������)���`!�L��)#�� 0���vR��lN��{+w�T5v���,���f���c|k�c���s��,F�'�
t�.Tk7#&����C)��5�"%���G�1�Iz�J���x*_8J�9�X��
L�z/ZI�0�T6��O�:���S�&y�Rd��� �)�m<������m�O��N@ ٪��$bG��И�����N"��V���
C�J��5z5QE�z���)&|��wm�$�PyZB��J`P �A��s��'Tr�Q��@��r*��?��s$!sTt�Ŧ9�a(�ۡ�!8(�YAz6��1���ؽ��
Ѷ W�ڍ��hwk��O"d����8D/�gB��X'��SH��ȁ�#PS�V�C�d�c��7
���׈���, F��� ��k�՘u�k��9H���1��c�Ӄu�bЖ��<�U+��D���۩N'����R
g;�@"�W߃�¸� d[Ph5��<�1�'&4�49��ձ�R�}�U��#t
#w)�����#�E�	E**aL���ꀨ��I���bdi�o��+�M�*ყ� S�£I����ؿ�$�^��d��#���Q���	o��}�����LQM�>��i�+����(H�pj���`�)M?=�߇ܚo��_��.˦���+�q_:*���r��/������� ��n�p9��+@y� 7'p�l5�uv��?����j&Mj&�95��G�䴰����Ħ�K?�
@�m�+���C����ȳX��;���2@a7��v��G�3;�k�,0��9�YҭF�����׬���?zJ�h����I��e�%�A87�*$�i-���YD!Iz�o�IB��$桄�m|0��f��x��6�p��25\�h�#v��@��<�WV���b��?�=lG�Ύ�����h�g4�g@������"�� m袔�p�@�����1�Jt,��}��-����ߐG����#k�W�
Xu���KE�o����\�Qd��2+���ɑ'�国��)pG)��&�ќ݆n����!eH�����w���� ._Ȭ(�:�JK�����wIM��-MV��WRբo����g�뎃/R����x��T'�4��598���y Q��z�w8�	���j^'R�-�)�; �:4s�hв:S�o'_s���0���tjOj�z��B{Jر�{�����$�%�@�����6���(�-sC��[��=�B)M{�Be�����]�#��xd~����5�_�_K��9?z�W�:|$�M�>��%d_�������6�ө�Cw�%M (X�Z^ %r�ׄN
��	�T���t{fm?YAS��t'�%�{��t� �K������"���&��^���@��I���鳊GZ?��u"���r���rV��o���\�JNŴ��Y/��:����+Z�%���$�ȒnZ��]_���M��U�LbU(���gC�2V����͍e�-���*Z�
���-�+*>ZP�����/�l�����.��YO�X�5�m]E�*�S��=�YW� 1�F��[`,)���iY�#�M>���:s�5�z3�A�@��[
��nP&?�z�Ȧ)F��v5&f���F�och�ޢ@���\;Bo�v6��w}*�,')�hK�^]������$<u?5����o��
����K�^�=�6��o�����χfPY����C�T����P�z�Z���>Z`ff��7����Rw��B���Ңɲ��}��Ԙ���O�Ѫ�%��jp>h���B� ��A�j�lcqANR����?���VM|�P�v��56�@N;����&cV�!��y�N.�ƝCP]��I����ޒ�e�F�=LR n"n��W�}yT�/���{�v>rլ�K� ��hC��D�h#u��[S̚�W�S|d��w�/i�{?��)�?-��������̲�b/�����i���v�M�+�֎���N�H/FJ�SM[���ѕ:�n�u(�Oz�n�`{�!
�؂U������=0n����:�o��L�<�֭�e-G~E1�v����@�V?�R��`	2���ã�KZJr��}z� ���/w�@�57�m��PƷ-js�=n�r}�� F��ȏ�Ƅ1V=��ۺ�3�t7���5�,��^oR����M^� !�3��3��-Z�H�P�ts��)n�Z�
�Uzi�����3��A ����mP�P�[L~�|p� ����0�w��0�fg��iF��@t&�Յ�=�$vAbO��ؘ����������[�r#Zvr�%K.�fy��fd� �!�6�9=���^@n3A��T �~;�`��
,��t��0�S�0�'�G-���=x��dWM�K�o8M���?�5����H�;�cD���i�Di�� %��w��q�g��L1@RZ����f�`���f�;���E3
5y��hx����K�ӥ�����XԤ����	�!~{�]��1��1� �ub�n��F�o��	21@8�y�j|6���|	��CI��������k��$E��ب/~B��)T�d7�L�D}2D�w��?
����=FJ��Oc¨��5�A2o�0#҉�w�8��!ɭ�Q)N�a+]s����� 4�x� 	!�G�%6�N�c�}��z�X���T�#�3m$��&�L�0��`��m��z�����̂����C�+T�?{�	��!)ݰ e��'������Z�`�h�?d0|���T���s$/;��:�cΛj���!�CWͷ�ͷs��뮲��ïmu��"��D~!v����e�sfP\��^��[s�?V��Ve�ݛ�l�Yo�W�Շ�'K���҆&��ch]N�_��]�j�<�PDۂj�B
]��J�-��?��|MaZl7�g����^��+�����8��+���S�fZv�.�.u&�Q�PV�Əy�4�;E�'��ѩ^�H�A�R s$!�kX{Uz�@�� 3�sW[VY�նU���$�Y���� %ܡ',^v�-P?�B.n<��TbR��7��=I��4o*x7�`΂�P��sz��~���-ޗzYn ,3�CvFɖCA���am�t��;XF���b�=��Ʌ��� 4��/d�g�L��*[���е	6�"�(\��$H�浅 �HcmV�K���b��U��1/B`\Q�ZL0��ښ%f����NhX���)gj�A��VY���N��$04Ճ��^�.��IZQ�n�A��Rb�`,},^r��рL���z	63۵�܆Jx��g�|т��b�j!�_5�R@[ 0}���?�ʪ��X5���+�}�C��Ǧ �ɯQ��A�K@�-q�J�B=w�J:�*�l~��#^e泔�V���L���u_����˲z��$��"{7)Q)6ŤD3�M�ps�{_�_Y�6T�(��!K�f�-�����KT�N�i��6�h��k�:'�вA<�O�� qt���!�qŴ�1o�S�*2P-���}���7譣�%M��:�1�1�d���f�5-��7�U�Oh����@���bA�j˟���a��������٥"��=�H�u�)ID`G֓I�k'����b�^.�˗���� ���EY��L�#�O�C}U�B+>����u-�_�x����#XK��M�ࠋ� �n4�h�H%9�q�k��҃$[��S�����'��s#0K�s6[���b����g�1���F�e�����R�ѡ�XYу����R��4�A\���J�$��B2+/�kzP<-/Hd��8�;���nG��:y$��j� E:BYBɿE��mAI������hy��8�m|<4�N����M@_F�Po?H���[�S��D�]o�ߕHRC�%�KGM�=��	&I�8�@�'0��cM�u�%m1X&����[���fr�[�8޳���
�(Q§L��d�)�6m��
ͻ#|�á��%C����KE�� XQ�g�������Z�%��g�Ϛ �������"��$�\#��bȉ@Z` 0��� K��d���3��d��D�I#����Fc�d���O���2�S �1@_4 ��	����'Im�M���0F�%2���G{/�ݵ�M4tO+�ȑg��]�nt]�8�sZ�V�F{���5��G����cԻ�V�����I&)g��p��=��V��=�tuh<�2kq�1��f�����w@�n��F�G���'/4�S�t�.�W@5�����&$~r%2t��(�paq�zM��	z�$��eV~�Iz���f6�ӄo�@ۈ��ud��|���#ܩ�X����Ǘ��u�����(���s�y��#�T����oC���FȜ�{s,�<��j��1�U�L�^����eb�x�?|\ײ���f��Җ�^R�ބ����ԜB]l�)]��41_�؏J���b$ށު�y�}�9���ɀ$�I��\>W��G�w1����/���f����@��W'�7�] MǦ��E��+�Hk����G�������%�K��A�<`�Rgk�U ΋��n_~���~(U�5���~ ��.Cm���k�9�4�+o�.�����%6�����E[8�p!��C�s%m�8�cSR�8b
͝ď��J�ʟ?�VFE�`�`D�S���՗#��:
r�eP��^#���@���^٧��P�c
�����0�e��,`�O5���ճ�޲f��P`�J���3"�a|���ߩ;v����rx��S�1Z�5�;��M�G�y�Ŭ(i�_�JjG�x��"��+p�?~F�_3���3�~�@��M!���!�6^~=�y���P�+��t�>�1[�΄"�7��N��[������H���C����s���<�j����=�s'�C3���p�C�����I�k���������| �ol�I.P�"pB{�L���>��MO����K���6L{�)���6=1�������q3 ��ߕv�)mi���2�Ϻ����n�e����B4�$�=O��$�r7�
�D�LE߃��� 훶�q?�-���10�9f"i���	S�*�r�+ً�UPF�`�e�Q7QC���E����	s��T�� a�����C[@	�l���[��̦�-�6�B�-W+ł5n4짻��DHHyV�� l�5�~.����K��M.��m���7�/�^�Y-���>��XG��]Y#��[L�1�@GQ���è������c�qouu����a� �c��|�9ҡʾc0��;��w���W@�F#e]��A'z&˕ t	�d��A_Rf������c��&���NF^��凥nU֚��A.��J��C?��8���*��J���a�]<��<���ߨ�����I&�W�2{����&[��U=��_��?n��dE��Y׭MS����}�_nܟ���mV]wh����=M����$������{�~{Z�uL�X��]DҼ�V�\��%rL���@�e���;0��>����h$��ѝ�����?i���e�/����VtI�Xc��&�5�BsU�H�F�h3�1�yC/����\T��./�=�#/ߦ2h�`�l
��ߘDo��Ww��6.�䏴hm	Y�SC	��������@��2�g�[ �A�daR+�ޡ0�X��	�ֵd�4��.�L��B��?[%�r0/arJ���zc� ��Lma�XWXD=N�T��L�S��=ԕ��:c���K�d<A�,ά4�_�����Z���m�jHh��ڬK�����u	8�}�q�Tw��8*h�A>�Я�E�	��ϑm����W ���.⋓��4��T֮;>=���	������?�F0�I�F#h��>LB�6!k��jx\�֜��5s��>�gM"�Ε��(]���d�r����#��wo�����_t2�����ɏ�D���/�,����@l�<e�jޭ�wW�a�����v3�56ש�߮��;�[0�j�nVc#{�ƨ��`TDw�'�ރ�s�X��A/?����k�V��j�g���i���v���;�Fs�`J�㴏'�����1C��&��p�I"��l<�y�6��Ye��Ӯ���=����� e�p$����|���w�c��We��ͪ���"o�ͽ�:lePL�����)̛eI�i�~��ɳ/XF|	���U��`4�n�YL`�@�f��V~��~��*0�7�����Q�1<3Ã�1�
�����^i���D�7�xK
�+ļ�=��=��oc����,�����5d]�����m�	e��X��_;�Y����v=*,�٥6e$�M[-���w��\�[k��
4�P�߸!��8�Ɣ.�H4^�س���kM$j�HH��#LI�����D��c�8����;:׀*��˯Q-����_שI%�/_�L�JX�}_��n��ʚtM�.�/1���9��k��`�Kw|�&50����I��m1�����LC#��"
���k��/:a�I�U�U�4X<U�'�xZ,������≋���]zb5Bw���������_���/B��8`@?2�F�5�F�٥�2�n��B�|l�B���Q�,�'GQ+B��A[��(��Z���{�A�k��@�qBM��I'a��$`{} )~�r��B6,�9Q���D��z�7nɘƸ|c�׎!�k!H��ix��(V�9,j����U)���N?l��O멆�uη��J�Oш`\����ݗ����u J�)����|�x�:�����"*����Y+)P�+��F������d_Be�n�5��y����FH�� �uս��H�&�U�-|x�k���\��>�����R��YTs�}�3>Q�U>K�R�[�]�����%�[���n��f���܆x���2�|�f�δi*��	�M����E��:��L��"��$�����I��&ƩD��7����֖g�uxmiղ{��xOx=�/�}�>>S)eU6/�q��L���B���ks�W��}t�E�G���1t��bh"�.��	A�:ú.�AI�����)���U��V~n����b���m��,�D�(��IK�4Y$m$�)-M��g��i�bn!�	����v�)(��X|�Y��;���T=J#�Tt&A;�z���<�$F{ٟ�x��hq(�V�M4K��Wqųpa���t�8�D1t^�T������4p�졉\���� �4��'�-�Q�W���c�+�G�U��3KQAb�B}ob ?��\J((��9��EZ94Pu�E����g9U�����on:S�H_���m�l�g���1��D�M���U+x��4S�lj�Z��cK�-��o��.Ɏ^�S����5���Ix��|�j��|Lcb	Bv�F�Й�i��K����b�^ݖ0+/��6����C:�>����oQדN�b��_�a/�;z���yx��%.<|�RC�D�\�8id��e��J�W`(�8�kY05xluq��Y�� �[8���$��uX3�޳���P��2K���]]d����F��x4s�P�zZ�DH!�E\��A���!F��x��x#g���=�	�2�E�ïS����	C�'�(���t���(l�Eaى�@�z��M-`s-l���(R�\9�wf��6��E��0up	�S;���4����P�ʉ�B�`�9o��X�)̮/��}J�3K@�=�)^w��6BW�V�h�8�	��)EP�YL��P3cc[�	u.��X`����.g�� ���yV�W��
P���xˇ����b"M���,el���hT��uw��^�t�Ȇ�6�����.��6�Zd��r%
�	�����a4������i���pcT��#���M�fu�6J|&%��H�GkKS��ln!���~ �U�69��J�H�\��$6I%~Yvk���F�${(�L�J�`�Z[)���{Us�H��a
��d�0K����߽�rzE�������ڱI`(b��?��k�,ݝ#:��7�b��W���]L�"՚ζZ������@/=�řP�Y�Hd��V�T�5|�)��j����|%{�e�
4��>bd7a๱Y6"٧�S7��!<�io�(Y*�����f�)r�(bd�/�!岯��W*H24��Q��i��@�A\(� E<�!.?���!�kŁ)�cqXz_Q��n�����O�G8'�v��X��C���P�X��2� ,w �t�N;�O�i\�?B�jN�[����~6�]�n��C~NUbam��dG@��)vD��]�?��`(*�Z7$~5��r`z�����1Y��v2i?W�N&m�r��tR?�-t��������B�{?@6#GV�x~$��Y�ܞ읎 S����P�em>����K���4�Kw�U!���W�V�b�}�s�!�k3 �뾳G~�����qY��Gժ�>^iq��3_��b��s�Qx�r߹+��\���VR��.�q��3�v{�<���Sx��1uDDzG+��蜤��bI�� �R�XNrAİ��T!��	�לJa]m��4T=��b��I�ڴ��c�7h?���Olq3HuqB��;d�&t���� �<x�C��U_#i?�s���`]���83�gξN>��V�Q!�dΥ�
��l����»��u�O�+��e����&I�ע|�#�@���9��x�j!��ɹ\�A9'G�),lu�$GP6��P$�&�u��6�$&D^��g��z$�@��Џ����b���3SЄ.EHB&���b�E(� �B{AL��e �!�E"g=&�.��Gj��{�#G~+�6�þ�K\�f�t�?ub�_�6RkR��EZ�м#��s��y$���Xgh��oQí�>�%��Ṹ[ Ձ]�s<�*6꯵8��L��:�?�o�M�?�tG�x�W_�_��h��qcr���HӅ�r�l���I�q9�`�[��|����͋�:��E�Sp��؜]�r8�v5,�+e��K~���4�w��a־�E�%.p��3��?�c�V�C#
���Dv�����JKe9�hp[�c���J�`���@�������b)�Ùo���c�ۣ�m�����T��Ě5���w���7���T[���/Ʃ_`���pv�֛����4|݆�������h�P�	Ĩ��[����q�$�s�*��	6x.Z���FjhM��*�����U�N0p�ɇ�x�["L�i�3���t}M�:��Ǩ�B����t�XN�N�U�{=���p/�kV��¨�q�yõ��(��[��V��}R�@�j@�!YJ�. '���v���ƹQ�4���`����;�V�:�^����\�'�����C�q�k������U��"��ʆ���U��֍$�{��!{��9���>��~��,[��q[k�!�Wgy떻�����-�/��p6���n�ġ"���S��]!�q<�a
t�{�ENCYm�ɳ��?��Xϟ��g"�Ή��`�JO]���4��Vb;�������bH �/c��6%ɏ�D����%���f��亿�k���=�s�����V</��&i�y�?��X���FꮯU~���:qr�C.慱�#��+N��m�D=<Wߗ���'J
bIf}��3��V�,Ht���F{ӗ�*��Z��x(���=?n��]��.s����骕'���L��`i��h�}Db2�A����~������*��Z�R$1p�ym9��'��E���O�}�D��H?�;�I;��)���on�e�>�����pX�'}�0N��j,w?�q�Z�A��ڡ;6A2�n�3յ��������T�id�P�7�Câ���A�c �ު�[�ؓW��xnm��@Z��Ur8X���Ss��-��Ujl��)з��Lf��9�&<��=lYA�3�	��m�HGh [Җ�0{Y��W/���-j�' �>d�����֖]�����.Ү���'�°[
��k�+bSM/�4ٽ�٠�M�w'A�~�p�괧W�^��J��.֟��� 5�z��'!���%#R]�s�9������O}7d���J�s���F�8�W�rX�!�7�ٜ����?�����[��+�����IF@��t�	�<�˫V��a������~�hI:����Czr���k��D�}�Ƭ��@�'�J��1������z��F�K��/�dt{v��Ԝ����)4f���ϛ�_*�^���rK��m�ؔ��R���_+���Z�4r���6����(�/h�ql�k`�����N�YvS>B��,?բ;����R�.z@��-�@���+�@���>�{]0Mv�u0�k�A?�%?���� %��^9�BҜ�� H��:���b�o�W����ot�5�iF]��Q��7���c��o�C�g$\?��}2-�u�wzKbd�d�G9�ד�O��z��T�> bx �����%{��DU�q�R��� >�7	j���й�pm���_%u ��c�u�cKǢ�9��2�x�nwU�k�(mV��^���H6���$	L���D}*}����CPO�I^����^�WoK<�4C��-�
\��E�,<ѣ�Om�����$�^h?����UD���H�"7d�n��E>��W^�%'�m_�E=�%��Ć�+�E)ڢ�[�]��5�MV����X��� ˏ�6of��s�ǈ�޾��2�Ԅ��o%�&�J>����A�Q�6�ԑG������2�����pYa�p.T�X\~}�ĬPv�PEoS�A���7����c�I�ީ�?�Z�`y/k�5���k���n�����������~��uǯ��r903.l��Ԣ.�
��VymNbq�F�&'?:�ǿE��]�N���2��[�U�WxspH^��������$�oQt =�;�=l9w���{������s����Ѝ=�3�Z�9s%1��������}{��f]�D��O�����nuk���ټ���N1�y<Z`��$��M%{��xA_6 ����Bv	�80>ߛ��U;��S���[,w�� ̳P���ؼE���K�)f�����ƄMwX� E�Ca'E��(���f:7p��6|v^��54�o�d 
�w�a�\��J�����8**�`�*P}�����D���O��
#Sr �ȅF�!����b��ct�4�d�h�J�#�p�n�0M��Gb��6�� ��U��A��0d�prԏ ��f?��0�)���TPx~�V�C\��Ρ���G,t�X���ג��n�}`_��OY��� )�����ә�+��@�-��I�zn�(I���-���</}= ^�A�=1�W�Z�?J��鐡z"-M����T��͈{��x���P� �~:������%�'�L�\���o�x����v��#��_S�����&5=z���j�i���֯R=�3�w����g���*z^I�k��;.�yP�t�ʻ�p2J �9x�A����`�X�&\���7?�.$���Y ��9;q����6S���u�z��X��nē�b9�jT�?���� i�m��	�ʎ�%bM���1V�ժ�^�a�f<z���b��tGU����&��3Rˋ�"��߷��q����3�O(t#}�az*��`
���%#Ϯ�'g,R�:�_����5U�ݝ"T$G�f��o� �I����0n1v�(�~x2 u�d'T3Xԗn؎[�W��0n(�,E�����|Ho�i�rCfX$�m*�h�R1
�q�E�9z�����޲݉\t�))1�W�skr�ێ�.��$�g��}�>�گ�&���jx�R(��|56<���}~��jZ���J�ݘ&l?_�l��w\)��/�Ww�5�9'�0��)1e�Ѝ��|W�����*TT� �\U�?<�*ڀAx����֨�$b�@��;�h9����h�+ZnK�|�d[����(x/��g�N/��3bɓ!�ň��d$���x@7�G�N)���]���ʿ���ڪ�+]W�$A�U���`�[��+V��Ǎ��٣C@{k�m����^����}�녠=�l��EH �}���mx�X���S�\	���]q�F���j��)Oc�Ȕ��ʫM�>c��i�r��Cv)dUt)1^�ζ"We�6Uϐ_iN�P�/��t�e�9���65D��
�=F�E�{���U�g�}��_�k�ȁ�_�#��1�J�A��,����+dS^�j��dMP|��mhf4���[�%��e0t�ҋ�v|��\G�>�z�9  ��϶ē���C��d�盓Ve��x?.0�)X�`�����x^��2�K������u�.��>�} t	ZN	�dtZ��_������qO��>�6hu�����������h���?���i���6.P��=��v%|pn$��T4�u,��$%�l��	Y ���C�Px4>���m��f�=V���f,�=��F+�J�\=��0���aT�����û�B���vy�ǫ�������O��X����k�9L�>��>����(��X�|0�����o��y8��#9aV�V�j���vx�T�Bx�|�-T��x���L\&�����[��o��w��GƵj ]#y�24�]~��r���x�Q�+���)��v����ɸ+n��uC�f��$�S)����a����T%������%��[)��r�U�6\��Mhx�g��?��W"�*ڴ�'ޅK����<����]p��R݃� o<��g�A_UX�<�_�6c��n�N�c�I֬��Qۉ��IgT�[R��'�z}��ӄ
�7�Z��~@�П��#^*+k����$�� ���8��B� HJ����Pط>P����A�&~
1���|�׸l�s�}ុ亯	�����}r�:�Y�U�{��u��XzBr�VJ^!G�@E�"H3��E޲<�|� iѥmS�K8���6�"Ko���i�`QB�o������!��s����'pj+x��;��B�L��x��7�^W01K�`3�y}ىĵ~6Q��A���V��G���Ԭ�����hf��pTI
�l�Km�j`�#\D���$���	k9��­G��oN�I��1��������cS{z3�#M��G;�s6�?�%�5�X�̓6�BB�J���>�	�<��p�d���R��J[[����"��A���6�&?LϣG�)6�8�S�ʬ�[�ͪ�-��b����Z�ZT���E0��?��],�'g�6�P����	T�)5'�M2��ʀL�՟EW�x%�&.�U�x3���[��,T.v41@y�Y�� ��n�� ��'ժn<�Zw��Oku5^\g
�������b<��N}��N�~���@Wh(Tشu��TÜ
�'`�����_���q_����
8�KۈR޲ٮyrd*�8dW� ٖe"�]
�ҽŤ��p�_7H�Aj�FY�	��$z�fӑ#ޢۡҢ/ KNh0����=�|��/��E ���� �6{��Ӄ�a�M+�_K����Q�U�%Me�R��"��;T��W~u��Yy���+�8��]�����m��؜�#{5�qYl��2�稘)z�e:1�.
HB<�ؓ������E~<���c�aՆ��݌�L ��"�q�wl+.�c��J*{�����Y�$��{���	䭷t	�`C��$�<�:�
��I���ݻ�ͨ8���@~�j�]���-~��~Cl7�k���@�cN�X�=�(�:�x��LbEʯYm�24��J���'�P��T��r|
��.�]�W��
\�b����r�p���W6�H����v�<��B���t�9]�l���P�8���5=�c���7���JAg/�[$��Ә�t�i���r�D�덭Tw�)>v<�:Yn�"8 jV�J���Ex��hgB�Ff����c^u7f�O����`�Ԝ,������-�#.Q�->¨*>Xܘ��P��OQRF�����
���?��G��/�BD�<�MkJK
XQO,�����Mg
�鸽qF�Ƥ;n�Y�6��c?j��!R��q��1T	�ϢYc��U�A�#�;�ܻ����j������)���V���r)�u��4�[_]��EX �	F������^�����/I 85��+M"�q1-]��U��$N�Ŗ����9P��&�~B=�t�}z4�߰�������������f�ߊ:��w�2E�U�k~xyM���� �<�明���l�}+��(����<9�j%��.][����mJ�O2i7��������J"k�Z���-@��ӷe��?3T�Õ���fq(�OR��\��z�Mw4T
�.����m~}�?���>����>��T6��=�o�[���rZ˪	�m5q�����zݶڣ��@���p���ȧ��]w\t#B�U�'D,��� `v˯4��K�ឌP&V�Id�{�!+�ۀ��v�s�Q��	c��D.eW�,n�P�T*�f�����Z���~w ��q�8M��d�[������.N�՝Ǩ�F��ox��h\�y��%F�b����f�uG%uLʶ���Tβ�����ǆN��36��ܻ�vN���"~P-6�8��KLs�I��	��}���+d���Ҽ�J�*�O���H,y�~��XĹ� �tGp.����i�1<(��
:��pi�cxX�u�c�hP#���\/��ۡdb��"6�75'�D�$=��C*��/����n���8T��9�"����	�еL������A��_P�?��cv�|�e��|���7*V�6�HM
�2�mڹl������ͅ�>~Ȝ��k}mv�8h;[w#������v!lq�:,�<ja ��w�y�R1���)��V:��/.~_I�H\.����^�X�אh�l�7汹��"��o����r8ܓ�| ��[j��xL&���A�<��E]�0o�E������4��1��0P5�d'1�?�����׍����8e?ߗ��%�'Z�7��P8�����U�a�p�E�f��98�ޣI��~�3��v:.����F�B�t.t���٤���#��hI�?TXB��R܇B����m�s�\���a�8�����{Qʻyq�u�����{�Y� F��I� qRq�5� �C7m���W��� \����(v�L��7W��)��Bo�;T��s�%zl������7����I�sIz���[`={:��wIZ��r��p$;��b��m�ކu�'�W^���$k��;&߀O����#����$�՝h��������b�\i�N0��L�&�磣g^�	Y��������d�3��i�"�|�@���(ئ;��Is���xk硸������wl��g���q\����:����5���N%��?����e����@���� pX}���ʩ�H���ˆ���qD:��d�������I��Dc{�V �J�=�u�Xv�]L�~�:��H��|�UtW�fx�,M��&�ō�6�Ԡ�pI:[��1P��X���Ԙ�ܬC�Ud�{��{�DZ_����/��cٻ^v�Ƅ_ c����m�d���t�6�Ϸ�<���l�Wʑ�h�=��c m0�G���x�Jo����cMЍP���{����N�}�z)��P��H|�	T&��|'�ė�L}ԬQ͏�7�<��W�s��m�ps�� �V��ŵ8զK�0$��!Y�*��x^$=�I�ARA�;��qЧ�ڬ��)��ןa��.�r������oTQ�[o��)~;�G�A����������"��{�K �i���E>�!�\ �`��>��n�_��-��I�0��2ر̘������[���rnUe��>�'W��57�m���=�;C��
���CK�sy�c|=ƫu'��ʄ+]f��K��}����.!�#7<)����X��I	]����\zEt��|3}i��d�]�_,����H>&_zflD+rQ����Q���"�V��@�5<�@l&�����q�j�7~%�i;f(�/#Vz&>0ƒng�zzo&��u�5����{z�"�U��\|�z��H?t+�yCq��E��B)�N�2�pŭ���D����a��H�o������D�4�6|G�q��Ŕ0琁0��MV��l�޶��D��7��e-�ǿ�VF1U���\%P6}�������&j�H�|-�*��J#��QP�ч�c iN%g҆�ǫ	��Q�I� 
	�o@��K`^�5��J�� :��;P�����t�FI~n$�"�j��ٛ�C̘�t�"H�8`�p` '��C*,�;<�{�*lI�מ���F�XYx|����g�eÓ���?d�����70�WpF�)���8	8|ʵ�W��3�֘�B_Ħ����������˺������VY�&ao��5�I��&�2��dH*_�M|�,�C��B���WH�LG�W�jU͝PQ�U�t�?����1;����A|�C����a��v���oQ4�� d��ߨ��0�-.��Ƴ�e��,��D�fF%|ZM��V��j#{��@4���5����a�+c��|���D����\��5��LUo�_)�7;�o�/jH���S׭�����洓���~�y�Nӥ:�K�Mrn~�q;5k�{`Ȋ��G(�҂ .l��De�)� ���fӛk��n�u[C�h���TS:�a��lD]������yz�?�5s�� �HG(��͈t�l�ڴ��r@����|3������ n��aA���l�g�-�F8�[�7�p�v$#{<Ұ+VP]�s@�1-7-:F��x���6A�%y��<������;��_n�y�3�f�~���I�[h�	1+�����C6��@a��'~���OK�Q�G��S�0:l�e3�X�ս�Z���#߈�/�,]����o�z':騣�I6�0�M��p�:d�"y�4���/<���iȯ?M~y�4#;y˜x~K܍u��a@p�Zԉ�bu�	`��e��&� ���0��"S�Г�8��}#Nr�g�j��X��5+���.F��	�\?4������ߩ��<�U��D6=�359��v��/&=f^ڹ8���� �o���Yӿ�V��\���\��}0 A���t�w$U���plXO��ZV���أ;��u�WJ>�ۗY�?����܀ZS�:��g��RXC���ߦ�<'�W�$��^@���<,ѿ�%���&G�Q�*����T�h �G�=�ͮ����1Ijb�a,Hn�5,½��^&�k1�1J~�sD2��x���ɴ4�&Ֆ���Ŵj�OK�#c�k�~����.�-{9�7-�iCk�^�4ֶ������=�BR�U��Q�I"��HQ����?O�/ڟ%Z�7T��C��=�l-�oЧ�#l���R2���	���ҧQ's�i9���x.ٳx�+����K"�Lwl/GwQ����{��r��*M&<Y��>�LɁ�7�!e\��Xb4p��0'G] ����;׳����~����="X�D��v���B>�
Z��wF!��zt>\t�� �3���w5%lF���̢~|��	��[�1����uc�`�k��8w�`3}�T��^�B6y�nRY��$T
s���u�},��X��S*�諥�������޷�EY�����ps�N�I��J�a5ؠ����i� �4�(���h�llk�n���-��fv�Ki����.�Ke��х�2�9����3T�����3��s����wZ���Y�#��:ÐZ�\m�R���]�G��5t�T�EC�RH�����M���B ��xM��I~r_�ݵ]�.J��X"���U�I5ῗT�ehj,��������Ӭձ���G���c	ʿ��W
s�7����/:��&�����[�����c�n���c��Gp�T���GN�Ԑ_C�M�&�ec�����~3����y�a�*�h;I�)�`���� ,Զ�ז���',� ^�r�0�bP�s�-�ϊ�G��������P�m�#��5�gh}t��:��4U�,����>���^Q���Ri�F�lwLv�Q�Xsm5�c��.�Q�0��m_w���$�-k�r��U�/���U'�>z�O����D��0�]��֦�x���F�v�7`}�햬�����񋛠6G\'&�x����Zz�ox����W�mZݼ�f��g5<W��AW�*���R溕���iai���f�.�ʮ]R�YZгT�F}�.dm��K�����n,y�:��B&�׎�R��z��E���m��V%B��BȨ{Յ?Z�)�z��'��nge�J4Ill���5 =�S�ڿX�1|��mF��yN�E��s5����{��OՖ�n�Z�b�i���ʟ��E��u}0:�ŗE��~~@qJH�<�X���&����iF�u�{N��˴�7s�#��^t��`��{`_K��M��ȥ�?Qi��m���Q=���O�L�=ꅴ��Gxu�~]F�{}!r��� �����Y}^X-�Ф�{�0�p踚���>�p:Fי�eZXS7���F����nr{��=���S�&�jJ7�aw�X�1`�m�rߒ����N������|��F%T����7҆ӎ2q`��|��}b*�P���8��j��t���F��z�\���Vr#��f2�+n�Z�eHOޮ�*������E��^N��LsӴvT�/�F�H����9��?��g�8��a*�i+�y��w䞋�L�7�9����r>	Ύ�o�u�Ѫ�q�C�M!O	K�H+Iݩ����S����]�����*Y��O:l⌦���[��x�p��&��3�;��ϧ=MNLK�i���?�mϮ�B�V{��h^,�ϑ��4���{=��TQ����Ң����B(�3fu��"%�,J��{UH��Qt*ͨ�m=��~a���:F��k���)��fM�W��G������#B���g�:��J18���}���j�6+x�sOY}jk0��s�
qr��v�</:BP���,���AԮ-��+��)Q��ڎ����z�ң�{��Ts�5��C�{��l���50`���yK��c#��|7��ЙQ�q��v���R�i��v��v�iRۖ%�����.8-�x�VC�9�Sۖ~H;�R���\�ڜෳF}�|
����|Se��q��� �'юH�a���DОA{J�)
Z����t�޴��dO��<Ք5�8�z��b�Zt��G�R��^���L&u#�ｂ6��U��Z��g�$�Wi�Ce�>,T����{�Թ+�~K����1������[-��B~Y�[�߉rz mgɂOjS��ci���}��̿&���[�C�FW(e����@SP��E�O��7�����ӡ�i��~��m����0]W�R��):����DTm�wO�nv]�M-����]o.|I�x�4}qZ���"�Ďwݯ���)k��˺����k�h�gp�wh�a��J��������$P�I��y�w����򵖂��5H� y�k���x:F�^�7�P!�m����<��;j�#t"�4����Z^:Gɧ��
��]W��I�r�=A�/�U�?��'��p�p�4&��)|�}s�r�g��My�3���_��'N�*���d��oX��5�ƠVW�&�2n��D�/P0'j��ZPh�d>0�u���L�7�Iz̴x�݆����.L�DoJ��f�F���{<?�>3d���6
=9{��{�S���芝݉��/��%ģ���F5�uѓ�h�E����9�vg��H��Oj�:tn���ʰ/����V��\�!�B�뫳�(%��m��� W�8��a�y�8�G�E��K�|��~�7��Kٔ��fN8�E�\�GtVci�kߌ��#������Ĩ�"�z[1�F9�֐r�t�����Ѣ��̉�q������S\��b=÷�wʆJ�V١۩C��]ig]k���w-��Is}�Y�����Q4�G ־���5�:&OsH&��,��p56�v�/�HY�q�\�<�[s��t�f�ԅ����J�b&��|Juz�`p
s?�������ܙ��ns�'~�8#�6�����<v���V��#(��C�F�9�2�kLT�Q��A���M{W�@4���5��E�xYF��V����b�c���ƤF��X��4B��|�IO���c/�$��=��պ�M��-^�J�_䕵�{��b��:�5j�'�:)F)���y���T�K=��*�j~�x��)��O'�R�(�0��"�!�ŏ%Oʇ��8�EZ�w�A��u�:��6s#S��z��Ɂ�Y�ze�c��r��-��|��k��*�����A��þ��3�R�Y�����̽��륏.�b����O�~&���W�]7�6is&��>�pC�����c�l��t '�Xe����Μ����Ѵ�IՉ��Y7�]��~kK<�77�F��(⦔�}����o(^v{B)n��1�f�$��q��ʻ��"�H�a@o,��s_�z���'h!�~��D�
�+*����2�-otLz�ǐ����9(�����K��Mo�ρ�ǥF^��\x�\�NS&~�����=|R�9���i��&eܛ>3\=������~�.�@�Y��O�I�;���Z1!�9��f�+����.�?A���1�Y��|�ɘ%�Yz�Gs�q覹����'�s����iI���-���@��)İF�7{F��&]9/1����fu_�{�^��=�`.�<��V� ��o���C%J�էw�ъ����Sޝ��{joўޭ׭��@����Ysmp�4�;� =W�'�A���� �X�p��𥣯2{C���H�{������`�kh
�=�^�u��L��Ӈ{Ԧk�~�*!��<�����]��z�������_}��c(�e�T9O?DG��*��=}�'�p�i����_ᷢ�Ҽ���^�a><�F����%����2�;���n������w^�@�ٻ��~��!��e�y���ڔDo�^����
��C���o��O�=���w���6:/fB�uL� ��=Y���Y���J����tN
hTSEf�lu��ϋ�@��8��#���>^��{�T��ӎ~����h�1�FKs^W[be��g����	j��3������)�.��HI������C��7e%�{k@{Oo�ׄ��~�2rB�&��y[�S����D��b��L�[�h�?�.3E��E\w��$���������{˱�6�㏞�_�-7������>��x��)� ��Uxݚ�g�}&�W��*��zw�v{����=K��h��e�<e�}(�Ѯw�8²G�6���S���]�Wg�>�($}���1��L=Mh���?�Q#_+?��/�y�z0j�$⯽�ߵzz
x���{}��i���Otl����1fzV��	# N�?n�^��f�rx�x�:��=� O랠~,r�����n��Ss��J���q�Y�d������N���.��Z<���f���˥ޝ'��D>�����L�O	Ԥ����//S?�?���h�YJ��X�|���5��L�K�wz�e8��>J���]_�/K����f~���,ٴ���ِ�	U11���-޿�8F�]ߴ/}�T�AE	�	y�s��c��?9���V9���AU�e���� ��O|�{��)q�]Ǽk=#AF��·�^�T���I�eg���1�~���X��[(�鈥+���2�7������/��&&��������}Gi3iǅ����*0��N������ʥ��̧���ߜ��6��&�G�/0J�%Mb�)�@*�w]���x��I�7&Ѓ��	��G\��/�E�/���>v�r}��� ݠ��*9G��x�<g�~S#�8�^Ln�+�~�X�mB�K��)�w���b����]�~ݷB�������s�Z�V�������r]�6�}���cC+\� �{O�����dѫ�t)m��Y��3"�.'XـJ� *?���g�{����&���&�ч�I�$��,��f��u?�����NZ���_��.�)NҜ莶NDn=B��;t���GV^l.|�߈q��耖y��L�;:Lǔ�?�+�i�|����s����7g��w|��p��ՎP�ˀԿ9�����e�Z]�S����71�˨�<����w]2���6zm�G�����}�6�C���Nך��#���SJ�F~g��!����3��b�1z���8B�tk~�W����&
���k2ݚ�5R�C� >��|�\z�6����R�e��W&׿G�o���Wp���������̈́�=^�{��T�B��6��;:��7���4ߑ��M{��w,�F�/�F��c���z���аN�V<�\�W�����+S�ݿ�9D�q�vt:c�I��=�Q|�����v${����䶼6����y���M�A�O��m�#�H����g�͔t'g�s�ẗ́��u��;�{��:yƂ�n� �	;���
����������w��\b�
�WQy^r�%3kc:e�:��{�O��d�Z���ʗO����w�~G�64�;��t�YFGN�ҿ�N#ƒ�����fhqmB��_T��y�ˋ��x1ۍQϞ,���3�Mx*�8�6$6��Ѣ[�'q�#1{ԑt��!��j�i��"�����Ir1z�hO��rzϖ��,���ٴ:SnG=�B�锓���ޭ{\o��?��܌.ϑ3fρ�������]�=���5՘݃���ǡm]_��v}����� ��ܡ��^h��$�Uf���o��Ęү/a���>���*�ݩd?)�i.(m͊�!�a(�|~�wn�~0���0z�%��TfBe�>"���M����E�#N3��[�V��Vr�;aP�¨����,�$�&ND*�B��XaV�
"W�.�|%Se� J�	�HQ.�M9OU���+%J�t1��M����k8M0(��x��*t�M����}��Ee��[�n4E�� h�6T� h~u��i�SY!h�
Y�	�_D^$h~�}��iZ]�4�)�$h��"YдECI4m�P�tm���t�t
?��+NS�P>��w3���+�&帠iAY9 h��ByZ�t���"���
��荂�H�zA�]-�m|mL�-D���2_���|���4��!�6�S�@�%�>A�Q��D�	Z!Z+�N���M�3ѝ���t夠�^r儠�D���VA��G�H�6A��n�A�]/h�z��4ݤ�T	���+e��'�"h��S�M7�(fA���2I�UD'	���Ⴎ!� �z����h&��?_+҂hE�-D�-hZ�Q��z��Q�X�U��ͩя������M�P�MBe�P�Ce�P�M��C�u��*�*����r�O�b �|�8Q5Be�P)T�b*�B%	*W	�`���d���Q�@�b��7�b��Q�*%P#T�*6�*ۅJT
�߯�V@P������DPdBq�o����b���x7��R��h2�v��l�]I�š�P�ysm�ֽ�2����4�}�v6[�֪�3���i��L))��=��h�:�\/y��=��{��5+��'2��*��t���7鶄|�G
@��� �i��!w�+�Hy�x��	zE^@|������uk[W]/��Y_~av�	�ϘV�=Zo^�C[��4�9u��`l��;�9�$�vڔc�)���}�M�(S|�t�~�qH^O<5�w|�<�!����?P,,e�����Σ����+��CR��_��o�v���"�e�=�ܝc�|Hӎ���nBd�йg��4���̹��X�Z�X�8���v�2}V�e����0{#����;���[H��qN�~�uy7����z�F�ڷ徾�ޑ�6AIrLrg����hJOo�X�w��p��~��rV	����Nsݴ���Mg���jx�nF��@���h�)kl�OdN72���ΪW�<�͇�h֑�ar�ܴL��<���gq2����iH;�L�����D���Q��+���>"ï7�o�ܔ�΍Evn�i�,�u�V���-,c&*cIe��ejcng	��}*�ݙ��z�ig������xg�Q�QP���TF�e�3�{��٩���Q.�{�Ÿ޲���f�$J����c�˛=t>كW cM�{?��ܪ��A��Rˌ���_昢�X�;ǒA��W��P�2��_���9��}}��$�-�t7�#�J���C�U����6�{�Ș�q�^�`T2��Η)���}�s��5 ���ſD�qqZ.z��� �i0e�b��8>"���ɹ������ O�~u��_�ԳVb�	���}C\����%�S�i��±#���
��p~�b��^�S�����N�z���\�����Hc�A�yȚc��gvy4�pӚ]T|��_9��6Y4��W'=�~�>�|H5��u�=�DӠ�����oĪW�B?�$M����)��Uh-V��?��,�z)�Ʒ�'��������/+�=�G+]Qz�J�=�m�3(�='VѮλ�JG0H��I�+���Q�g���)Pr�c��F�z�l
_i�n��O���)Z�#J��򥜾��g��Q�=�{�ORB���ePnxV����L�\H]�� �t�f�^��
~�����o$Ғn�Tw���^<��?����+�_��"$�y��S���c���}*�9���uB?Jιj�кwP+=�^� �娀̩ฎ?k���uf���w^	�@��9���m����,W�0��n�� u��cZ �p��+�Q1f���ETN��^�G�v"�����[���..�b�s.�iuL5��.�s�3�..�x��]�����Ǧ������<��K�f=�9˿UKc̮NOv�Ѭ	{���u��2��r��c�ӎ̻?Ѓz��u�#�洳���؊��q?����??F����+A�z;���O<�'y�3khs�4^�xGe��n��p<�l��/������%�|
e�{�������~`~V��C�靃&B�����}E�JP�M�Z�}�|Rm�p����^*�1*cJ�Io�2�'�Y��z9 2iMՑ��swN>�ͩ:��f��Z�0�Afw�p����_��Zn�=��c_�T���k�3�����S3i�����)|k}���-��H�^���_x�_,���Qx�{϶{O
��D���OH����gލ|A��ǩ�k�湼���.��u�&q��{-.��qm�����j�!ʬ2�g۔��d�k�	M��[�9��fw�g�ո���e�ϸ��D{����������I�ʥ=��*�=�(rx�꽻MX]ӣ��&�Թ����:�W��
��V��R�O�%���ړ/"��� ����ր����(6�h�Kk�ǡ�Qe譾��oU/��nWK����-��9�S�̈́@�Iܟik����a��]U�g:W��������g�Іͦ,$��5'�'NMt������Z|폳�b��]UI�9L9i����"k���3��>@�F��;3�[�Q8[��D�:����Ȩ��G�|yj���m��[���nQ��oQ9|��%|�4���{Y���LY[M�O駶���م�	��_�B7o�u>�A�y���d�X�,�OE��0��gn����*��).���Ȁ�=j�{fSO��_�����P�Zuv���f�O�ঞ�������oz�u瘔淺4�u��E�^�ҕ�K]8�������}�w�^.�2Z��K�&
\$q��z��J�)�����ĳ#.h�8F�Ib�D�D��z���G�k?�xFb�O?�C%^,�$1W�"�K%�+q���.�D6J�#�B���J�H,��B�:���x\���J���2F����%q��r��$n�x�ĝ�I<.�D��
����_(�5N"K�7�۷�F����Z�v�{Y���{�W?S�����������
u�Pi~�?�cZ�~��`�u���Z��ZD���u�2_Ze-�Ra_R�`S!_VZ�(�XK�8�=����q�deM��[co(XZ0���6��b�gyia���>�t��ll��b����`lQ��Z�,�X66c�t����JǤ�����
cYE�b5���e֢�΋����Cg�ڐ����ʸ_{�z�Zo<�ʌ;v?�����绵W��/�Y���^�5@�M���Ć��Ӭx�j�˘��8�f�`S���]c��a,�!?R�HÖ��&��i�5��(à�O/�����|ߕ+h���1��ԓ�������I>|ә���7�YY9+�;�7��%�+��l~�1��B�!��o �+����%�:{�#L2��3��=��%|6�M>|S��R�2��pY�f��:n�j6}h�����E|�z������Wr�������~����G�~y�+1�/e�lڮkOHsm����]~cyŲr����js�V����������XPVV��ʙ���S�"�z�=h{?z̵'�i����D�M�Z�����b���G��8LD�%�"n_b����.����,8���C233C�4��rƔ��>ZvyR���>p�ț��Ă�U��ғ�}�V��&I���v��W�3�J���Bke%C��d����b+�s{���e9Jk)��F^j����f�F�c�lJ�,?U��,��kz�e,�sX��g&��i~�2<i��"T�8 w�������]�E�*�j���%��!�U���ܖE�|���e��-����܆.�H����\)�Y�U@=���_�k�R�,�nᚓ�O�F�[�]%=�5U��1����.�j%�獰W���E��s����5����������O�y�(.Ky�]�D6�e��"{�
�~�ςc����rP!O;����d�S̖�p��xoz�Ä��r[�V#\��l�L_a{P�VM)���'F}�{�~ uOw�O��Þ<�>v����
{T�~��oI�p�~R㯧��Y��'O�E2V�/6(.ȟ�v��]�/��2��/w=�wٿ��ڢѽK���x���K�o�)'�������.U����/�ZY��X����RNM����&~ozW�5���(�R�jť<WZ��%_�����l,�>,��;����]��-��`)/�vn{�����WwT������R����P��w�S��
�Oy}[��&#�5[�rI��5�'�~��C�QJ�%\��ѿI>����/����Pm��!EU����b�F����y)���[7W�s��a��[I��T���~Pg���q:��rդI��R�����Hy�����$)��򶏅� �)W;�z)(�	� �>)�������R>Lu�Cȍ�{R~���N�~�R�\uO�oV�'��J�V��)BE�^��_B�J�9��Sk�t6
?#RڿG�j!ڥ/"|�m�16	iM�/�KdC�@���s�2����t%�[�������v�7�ԏ�_#}�C ��.@N��i}��� ���&@~G���r�f�W�X��ƌ��[!hNژ^A�qƢ��cv�V)���e��Fs��^`/,Yn̰V�Km*�qrA�U2���˥A_�.#��Q�ʍy�m�@��Yh�Xf�t`�Xht�ح -v؋�eIAy�bk�q)<+l���awr�R|�e�E�-]D��!�.���hyy�x��a�x�Xd�rCt٧�ќViAY��V?����?���rƓ���,����g++(�.��SP)�\��XXVQ�[�=��~�ЯXR^jDҖU�.������e��J��Ŏ�EeV?��Y��7�Yf���ܡ%�,��E���p��K�ᠥ[l��{:�>|=F�_�|o>+�;�AQieW�-)���o{�?��?������HĔ�E�|����Y��-���ż@�*�����wx��DE�O�QI�ʔWՋ���dlą�&]ɮ��J6�X��� .&��Hf VA$^��%@�-�$�8b,��.f0�4	���\��
��[����`��+E;;	]�+�7��O�:�Q;,.��$�S����k�m�e�@k��R���)*��_\P��RX��QRZ�+�t���
H�y�E��2 �W�:u�Z���.��$n�X#�Jb�D��|�f�)/��$1Q�p�F��%$�I�K���$~���3?��)�C��ē�%�-����$�x@�>�����K�[$6K�&q����H�(q��z��%�H\#�Jb�D��\�)%��x9#�'�Eb�D�D��D�Lb��2�7J��X-�Jb�D��d��Ϝ�� �Eb�D��$�z��2=$�K�H4}���\+��s[$��=B��̠���%������UY.�����c�
�j��I�/��Rż���t�J���>CΡ����69?�˙�GbN>�A�T>�]�g�'3/���v�D��)��E|��.�)�3ت���տ�?U��Q�!�[������XOr��"iB���K�fֈ�2�o.��6_�<p����1p�,�O_y�pWuO�_�O�G5�|e�bɒ+*���%�|F"���3��h����K$2�dX�uXd�f��K��3��t���P5Ҝ�����Tg�o���'|��^Ji�C=}5���h��6���K�.�E���d'�Gv��r���!�d��*@W����3�^*)�K��^�!��E�V�<���T�s�YN���̓�#�g�_Xu�mի�QA�V}ۭ�q�����k׮�@.)�:��C�đ)�s�YZ4�ͥ]y���j�b�KII�Vۧ�f[f�u[/�ƪ���--/�X6�!��>��j���r����]��`�:J�Zs+lN�W]�	�XlF�|rE�099'�X��ҕ���_�g��K����u����{kz��s���i~�����>���S�������랦%��������/h�~A?�ו�����~q���|�~t�e���?6�]�T��x��շ�֬��W5�����~}{�o���;������{�x�}�6o����ض���yǟly��G}l�㻞x򩧟y����{��{���^|�僇^9�v��㯾���7�|����o����������~��'����Ͽ8�噯������z�&(8$4��6<"2*��N�/6.�� C��A��f<�����pd�E��d���I��OH����S&^�:�ʫ�6,���xqI�7�-)���d�t8�.�Z~�u�\��һ�-+V���;��m����O����9�s��i�9�g�^;sV��9s���B����+�?=�������SG�dG�����VM�kd)wߔ5o�_��9�'�ɓǍ����g��o~�l_�l(����/kJ��{+;.;9c�+1��b�#��
���5i�c|[����_6P�������3=@���>.@�?!@��+g篞��-�N�//x�� ��<�����L*kx1���DަY�%_=��Y�Gb�b�|�����*�6�x�+1-W��׮�h�u]���o���osG�i��/�Wwk���s8�=�U/,��b����Im1�֓��9񯟸������17�L�����MV��=�����~W�tkO�&��>�4���JxM]r_>�?pվ]z�n��raw
x�}{����W�n �N��u��#��{�wJ�[6���w�?���>z?䗍��sb/����^/v���.ս�K�}����Q�P���`��J;�΀��{ҁ£�w�'�{Ώ��ә��6Mê`_��w�)��}�[@���Ξ�C��wP��p���$����	�տ�c����%;��/?�|��2Qf�_�=�R�w����GdWO���=v��i���N� ��,y�4�Ql��zv��6�x?�/�i��x��HM�[�h��D�N��:���"-�ׇLc��o%7Z��k&7�CXtQ��S��n���lS�ճ����c��H-�	w�g�K��X�������,4O맧���L��IrAcB䓹� 
���%�� _5MXd�a��g'��?dl��k��v_��ժ����nf�6��M5�nj�4�a,�(��b	�J�D ��g���"�aܯI�w"?N�G��#��p"�����q-��3���iՎ��y !"�E��}�j䓓�fa,�(����;�l��7�I�5�k;}�mh#������B�)'}��	�	Q!,j���'7,�ܨ!����A3��[�j����w��&�i�p�b�PW�m��_Jwc!̐�"f�񰵜|���!�G3�.��h7��(��E��[��z/B�/��O>B�F���X���kt!L��жठ\�3E���8���fw���� ����q���8 �v�u�3�G
�����DY��G���z�=5��<������16�"��@����5m��f�O�ӓ:�����ȯI����~�����M� �83��t�������Rn�q3�H����~��j��݃�|Ҋ�`�tW7Z��:Z�M�3�?b���!��}����eڃ�^�k��#�1��X߇�����̵Js-0� ��塒_%	�o����{�$����j�s�O�[�tϟ�qBo�8a~���I޿������:	����K��)Rn���R�C�?3�������pWꯓ���W�;��7	��>��S��Ӳ~y����~�m��EZ4qa,���"p�ަ	Ѱ��]���/���~=��`62W38�F�L�d��:��ǵ�k���J���E�̐���2�x��c��(��9�=Ҧ���Q,./��`qvi�=(7���%��Q�cl�D�Q��nn$��`�5�������<DmzC(�%!�%8�P#Y�L����J�P�ݜ�س3��8H�:ĭRC�ar�iS��8���Ty������m�8�M��<��0��ʗ�&��|y:�9դ�ш:$)F�ʗ9���g$_x��ţN�G�$�?S��xGd�m�z�y6�E�0 �)����|���4u#Ĥc]y�燨 ������^���v5���L�s�y��y]y.���(\65���F�	�D�:�N�cbCX,�?v��kf��ޟ�e�K�c�v�I8_�Ο9�sp��65UT�s~��Gێ	
wƆ�l8��ѓ��g�~��1��<@ F~�+�O��ۂX-��gTgD��-���j�~X���M���|����*��=��ŵi!��������z��E�l@^?6 Y���Ӧk��EY4�^r<Kxeë��?"��H�Fh�������mq��l1}�Z��<F�<F1�=��ǁ}��f��3cr_f���nh��g�u���,a��%�&��	�'�>a�e䟛�Gh����}ۣ�"Z��Y�d��8������1���H[�E��'��F�11a,�3ޟ��K!�^�y��5�q<�v��tWkS���%z9cIw4�0�w�az���G�jX��Pԛ��PF(#�N�%$E�a�El����0�{*#�9ȃ������DA�	G��I�ˆh�e���f�Q�F<�&��������P8��fv�U�f��հ��P䳘����?F:�w�լ�7h��`�i6at$Tt-���%�`�4S�0!�G��zm��8�%n&�Ԑ(6���C�>�C�'�h�ou��#�[�/�C�ɓ��>^�hyݣ���h���������0u3c�B��y al8�x�-z�M~�մ0��W�3��>޺���'��B\��1L�<�gz�O�N}=^����cg�{�Ԇ툟�.�xZ��XnoB�C�&P�aዀ�"ؠ}:6��Ah����#.W��I�Wv=l�*;^����%ϧ}q�+���$y�Z�jg�Ì�����l��@�`�= q9`|�M��fhh<�����-����_$ӯ�vz���>��NS��:k ��f�v��T�O=�ز�Ў��5e��~��r��/�Qߦo�;>")att�0G?�o�gc���ѩmki���c`^�tG#я��t�]�P��<�N�k4��5����L�p�����{]v�!Ʈ;�U�1��(�^&�����s@Ԇ�n�A��9Lu�@g?Z�wgK�/*�;_{|ʥ=�I���D�mP/���L���qYw>}�@È��%iD�n�[��I�>��e&%Q�R�E]�6jF�m�q�ݿ��cp���=-2|?����\����+����5���QP^hE���]@K�J�W��>QE�u��1EeelFvf��<)a��,(������Bf:�r�*���Y�ւ"��#�슊��)��Bb�,wЮ��3�|Yiy��'��՞n�Ӆe�������lk�Rk7��i�_E�5���̱�a�W����2�v���z<d�b�"�/k���ۭ�<~�'���fJY�,�cNA����s��%K
ʋ�K˭i��!�n�`���Y�KJ����^�UU|7dvy	l(�y�	�Cd����^����*3����[�vk%,eR���3DġF"����i��W �U�
�5jH摌��\�|�bɡs�VJ9f�[ZdM/)��U�8����;��A�Hy%2D:ڶ�}�9�y��>ge	�1�Y\l�#V:��rS@"��Ͳ���W8��HO:v��+��fG���H);�Q$���Anҹ-v��-@$�hs�\�2��j��� �#2����Sl(���N�VnF��4��L�� �,!��xN��|vO2�H�sh.{��򆺑�2��D�r����4�k(�2˗��+����,~�r.{�Bؓ�|��j_�k�s��L�HB�����+-�Q����������J�uI^)|Q��{[���	U�l.����F�����Ctr+r[iQ:���V6A�'�?��`oNʫP�sP꒛j�eH�'u����i�4-8�� �q��������o���&R�d���)F���\6���UT��f�2gN��V�3�fN����1bmm�f��� LPo�E��Qg<D�X�i�kP���6�;�!����a����@����ɂ��h 5�N����M�66A��۵���oC��a��81*Iê B�av� �װr�=�'h��B�Kְb�� ��jX�.���4��(��r���5��1�
B�,���0�����ɢX4C�]�֏Ţ��g�� ���@6�F �������=�`i��r�c!]����Զ��ꬅtu�B�ꬅ]ff̒�]�uii�u!���3�[�C+ϥ��b��F�0Υ}��6[��a-^=w���Y�ϙe�V5��B=�v���#,�xL�y��\�[�΅��f�9�vf%�O:�vNI�x���I��9�'�s�O`g�9��'�K���\ۉb4���N8�>�=���N�z��L�I��=�vΞw��h�O�Ci/�s��scg�8���H�7�}��=�����"�vҬ����}���O9��9�
��;0M��"��W>�=�?�w��`�"��s���1Kr���E�7����Y��Y�y2Y�#����9e�KZi�������%��=�ѕȸ�`��o��0��C�G��{<Ջ5~����ԏ����y��_�+�������_��5���ɞ�@�����s��?5�S��?5���+�3I�ȯ��Ց��#7hIWm/�%ҹZפ�����0&�a�ǳ�6��p�R/�G��4K�����;�O
uO0�_*�iR�.���L�>K�\i�<�v�T_ad���Aөv��0�_-��Z�R�%��H{~����^)�$��U���T\������7�q��Y`�� �ֈ��
�Um�$�H�H̗�+�$1I�p��q��$j%�Hd�e�H�\b��%*�%�I�'�i�o��R�,q�č�%VK�I,�X$1_�Ib���37R�(� Q/Q��~��G��#��[$n�X#�&�D�Eb��\�f�&�)�$&J4J4H�Kd���J�I<p���]R�M�F��m�%�$&K�D�Ab�w�=���z�:˿_��M����2�g���2je��(����~w������^���ү���B�����]�����<����9r�!(�oڊ���州'�����M���v~e�iU5�m�߽��-�^�_}V�I�c?�?M�N��|r�@��fe�u�ۿj��E��7����yÛ��;�����J�<��.�h����B��s%j��)�<io��_C���5T�Y9�X#�jX�sm����Z<��|:���M�~V�+������u�sބwǢ�
��#h���W�@��9�C��,7�a��	��4��`�@�~�g�N��}����v���&�� �{�O���v`6�m�!\�o����	3!��	�A�A���&�"4�f�dо�}�_��4hB:����|7a.����F4�6h�?o���)���?�U#���+����I����=�M�|��	� �&�BD��s�WǸ��]?��t�pqn��`х�?^�wޘp�H�4�+͠	߂X���&b<���-᧤�_Ñ�����=�K��4ᴋiϕ��k�@��p���%�8���,�q�D�K�a׍F;�δ.@�g0 o;F��3���!��G3�4��"���x>����xa��g�^-��z�SD>�=�Iؒ�Y��K1�M{��/�D'C��@���[�z	����t9 <�r��av8p��'�\�+����6`x��i��e)�'x�Tw �H���<t�a�D�n.�hmn��0�&��J�f�[oC�m�W1�!���\%�i~!�3�ث�[q���N��M�lMHG�E��4��Ak�� �@����� ���da�A�YI�$���"�`n��/B�?А)�	C� o�&��C�y�[�������v%�'��Y�k�K�~xQ��7ӧ��0;�����~<�t'02�t0+G�-�#G��,�.ԫ��3�ޠ	7@�����M�x-���ɵ��~=e��cg	�Θ%xr�o�m�I`d��1 g���������$�.���/�ڀ�����92����B<��us��z`t����y���|�/������n.@W��X�ԭ|������=�?_��A� ��~L{XT@{15G,bl��Et�<���p]��M�@�-~�.�ye����Z��-��� R@7 ���} ���ghv��:�ȥ��:8}����\��R6Ct�&�P%�%8~9��8IV-qE��!KԳ�.�5���'�%m�0�gp�
a��ېW��xs-�5�+��Ԋ|x�����t��������oDx�a����h[/x�%M��z��9u"��oI�m`��]�{;�z�z`��>.��
�s�n~�-�?��q����ہw�~^|�a�Q��w�<'�<���w
����'���ɒ� :~/�0�?��w�.=	�t7�4a���?��&��Q��z����- .��J�n�8 ��	� ��Cm��~q��[bx6�t�
�f����6#n��@�E�Kعqu�F�#�P�7'�/��!~@?
��u5�����m@}��[��Bԃ����P����G�m��?����� ����Cg?(�*�ڂv�����8N}n���>$���>�z=pȣ(����9�J;��w���&L�)�	x���?�K�/<.�k�ݻD�����P7 WAl �|�)���ϟA=C�$p��2�='��c�>�k�'�"����;�A� {^�5�/�(�k�'��/��|�%�;"΁�_F_t.���蟬��e�n0����x�#��F�����%�� ޡ�
tF^%`h̃���d�&��)A��D;h�s��VQ�]�#�>ݑ�D����{?�.����n
�7"v�a�?��?J��qI�4�I�]DN�4�\I.�4a���΃m�&|V�t����&���&�N�_�yh��:��4��&���D^$i�Iәc��	�$M�$i�}����?���]�(C��6Wo޸�as����6��ܾY�ܹ��f��[�[�[[�[�V�_s���o���m�����~����M�M�Ͱ͸-�9��A�Y�l:�I�tf�v�as�������K�R\ڶy\:W�l�nik<��ި4v6�idM�&}���ؔؔԔ�dj27�6�7Y�J�lMUM�M5M�M���5�4�jjm:���t���Ii�l:�Ě���fC��9�9�9���ln�m�o�4�4ۚ����k��7674okni����|����Ds{����|�������0�0�Hܑ�#e�i�yG���%;l;�vT��Q�c㎆�v��ص�uǁ���yi��!�!��ְ�����A�)i�e�mS����@�����o�޲}������m?��}���s���Qۨo44�SM������FKcI����������qccC�Ɩ�]���E��4q�qr�ـ��	/��e~��&�E�E�ŰŸ%qKҖ�-�-�-�[,[J�ضTm��R��~��-[�mٵ�uˁ-m[Nliߢl��r�J������~�~���?PK
    +Q�H���$  �  0  com/smaxe/uv/na/webcam/IWebcam$FrameFormat.class  �      $      }R�o�P=W�(�Ӂ̩t:������3>���df1&]|��+t�2)l�C|���MM�>��G�[J�-�I����{o۟�>���:4�:��8� ��Up|̠Y��x��w\���e�Zm��\m�����``�+���Lb{[zU�l���~S�I����r�"��y0�}�a��E(V�슆OŋP��¯������tkuҦ�Ď�����斬�4�Gz�i�^�^�mTe�:��BG�u��:`/���1��a�a�Z۟�\xƐ�
k�s�L�9�����a�u0��~30�RpS�)�8���c�+8��\&��Wp!A`%0��	dGPP`+(*X`�����?��p<O�W����<��џARm����U��'b��)���r�Ԉ��Kv��E��d����.��Cw��b�Θ�!.�iL��$1S�؟���)�	��@���;h�^�;�7A�����o�BM��Ҹ���W�U����7���_�}:��ԑ��������D�
�S�9��3>������b��"��E� 6��M�PK
    +Q�H�>eޣ   �   .  com/smaxe/uv/na/webcam/IWebcam$IListener.class  �       �       }M�
�P������8	�tpv���V��� ��[��os��(Ѻ���@Br\o �&ii��(���gMR1��J��/L�m�j�Z�Gi���%GMk¨�q�i��Ĩ����%��۟]�Y.����ZĄ��`ٗ�qN�G���=Z���!ڬ���PK
    +Q�H �#�x    $  com/smaxe/uv/na/webcam/IWebcam.class        x      ���J�@��јX[km������:;�B!XPP��4JJs!3�n}->�%������@��?9��9�����{�n�Ҭ7��ȅ�T2�0�E�
���H%��X�{�DěW��?'�72�F�EB3��$7�Piˌa�+��o��!��P}�3�c�C�Je�P�;��"���a S&�|D[�ho+1�eE��k*��B�\j���9�Nґr`;pL;�uPf8p����"�	�L�˰#��1p���1y�@������q����[�{k^��?��������y��y������[j�ē�PJ*���
�h��b��l]�6A��-�2E*X3_�1iX�x�ڈV�rM�.�Ur[�}����c^PK
    +Q�H����   �  ;  com/smaxe/uv/na/webcam/ScreenWebcam$ScreenFrameFormat.class  �      �       �PMK1���6�����j���^��ޤ�Ba�
z�k��ݪ�gy(� ��R顈b 3�`2�����;��	�a�����Pn�����c%��4���za��rZ=��T[�ܮ��mLsm�4˭��~1_��1n9��k�=l�ӂ�@(PU����2J54��[�DD&ٽ!4�bd��'�(LA�~4��5�=PB�XE����"�]�NB0���ݠ�X.ю���k�>c��$��/���� PK
    +Q�H͂���  �  +  com/smaxe/uv/na/webcam/ScreenWebcam$a.class  �      �      �S�OA���v�H���F�Ti�ꂢ(E,�1$BhB�L�Xhw�vA��A=q�B�q�@"�xл	����f�!D�d���7ߛy3o���o��#/�5�� 'SS�K%'�Q��|*/蔠�a۱�	�8��F��%��r+f��6���n:�|Ë����ǹS�����j�2[gf�9��Ć�W}�u$�?��d����i`���-_B�i�՚�b���;���r&4��qV��S]��sv��ZW=��g}f��y̢��QJ�����������=:��QѢ⼊VQT��hW��n�2�Ɇ�)�B�1�ha����K8����L���9o��;�
���Ѭ�":4$ut�I�k�u\p��.��lJ�R�K/-roG�w��぀�<�X���Ѓ���p}z1@�x�-Q���po�̪U^E�� �2r�>�^ND��T�2ͫ0��%"{�H`���qC>@ƈ����$�~�$J�$uRRY��� T!����6�_��qh|�pOv�T�D6����T�fv��ۡ�|���r��]$�ߊ��
I��ek�ږ��M*G����0Y_j��w�9�n
�o��\���-�a`:}���f����]���Z\lR��%������S`�y���l���!�PK
    +Q�H<S��'  ~  )  com/smaxe/uv/na/webcam/ScreenWebcam.class  ~      '      �V�WW���#�R+X�0�������`Q�ې0�$4�j�Ͷ�]��]l+-$*m���=�E����;Ʉ��9��;��������� ��	��zM�/��j�2�Lty��_��W�%0�E;��n<$@h�AnET�4�d�Wǌ�&��?������hP������U�?�ܽz@{"j���f�T��6�W�n�A�PnlPo��#A�ຉ�קG-�E�-c��hZ�ʾ=���$c!���U�\5�n�o���Q���"�I8�Z�4���֌��x(%�M5(��W���﵊�ڐ:>j��CC��xD5�pH�D�DF
PHo h����V�dD�.���Z���D���(�����V'wGD���%Y��ڴ	�O	�S�T	�.
Ãa�V��AuXs'���<�V/n�"�%��PG5kc�~���ۧ��Xb��E��ô�сB�J%�C��l�)�RU��A��):j�S�<nI���f�F�ǈ�!B�pRT~a�Ƒ�G�a�D��(Q!�R�J�DT�PD4�h�Y�nw��*�n��y��{F�lZ�8���r�o�IW��F��N_&�$*�-�8�ynt5�n~��j]���m�vݬ
i�5�e�Z�#��iC~�m��<m�9n-���'�jP�Zη*=F:U�\rv�IwYz��s}�>�E7���XkF���31ߓg��k�׀o�qnn���wK=��)�*lqe�8��Z��|[n̗��q�6˸� ����A&1و.&k�-�=2d�Q��d�@��R�QA�}LM�,+dR�Dd�!�����e�Ǔ�����x��T�0(c�<Ȩ�&�����2ng��8Њ ���e�,��(��8�	&�L�𰛇�<3s��e�I؅�%�;��&�2y��q��_�Ё��"a7^��ū����	{���%��.</a/ޔ�(�H؏瘼]�6�g�5�AJ=O�X�d<0��6�7D�uT�F52,��{B�)u(g��1)g�LNoa��0��P49�jr���.��$k*:E��l7��ة��B��'<3X�\�Ƿ�ξ�9|B�S��(�.��fS��!�Xb>r�B�X13�6�;�8~Q*��<N(�<�29���q�ɴ�4�3���5���<�)��5��i�)�>�В�-#./Tb��J\�C=�K]������j1�To��7������.��h�-�C{n���q|�cEo�=g'?y)�ގ�TQ��E!�쳼�SJ�|ŕ�SQ�����ѧ�͉8��r�1ï�Eف�d�j�� :	D�%+��Zý�[��
�r�Rw�1���P¬.���I��͍��&+0�T�˛���������Pje��8)��D�"D�ϭ�9S�������0[��%��/��e/
i?@'�<�kL��Ι�ǥ~�j2���|����~�a�:�b��g{���櫘/���j$���9�ǢF���9��Dח-����{���,&��e;��+r��-u)���V���O$�I�De�EZ�����L��t���
�6�W���l�]��e8�PK
    +Q�Hy�{  �    module/_004_.class  �      {      }�_KA�ϔ뿶2��ffZi/+�SE/҃ �`=ɨ���l�}���(����;�,��<ܹs�����/ E��D4�X�U�c	[�l��.��ʔ�sͰ���|%�-���{un�����0�U�V{�F�P8o\2-y#'wZG8�6C<��t��=.;FͱM�!eȒ%KJ�rt�f��o��Y��8C[��CB�>�Jt�#���_S���&쑰�ؔ��Ð�ؚ�Qmvɧ���/x�����qe�3��;�t��,BUvڣ�m�8��G�O*���S�R<�������1��]A��0�#�:eig���'�H?SGQ�'Sa �R��)����^f �6<��{������+�������?��=~��S��f���_PK
    +Q�H��Y��   ^  X  net/java/sip/communicator/impl/neomedia/directshow/DSCaptureDevice$GrabberDelegate.class  ^      �       �M�N�0}�ICCJ�' 1�1�H�,HEbw������v�w1!1�|���ʝt���{w�?�_ ��d��.����:��Fn�/Nhڐ$5Rǰ܉Q�^�-lw$Ý���W�V�QR��C�YM��S.��}��S-��w�Ш$1l���މ�%�PO[�@^`Z��0+q����]|���e��Ɛ�{�=��I��,�c��tv����{�g�f!ҋXˈ%f8�f�PK
    +Q�H�MA��  �  H  net/java/sip/communicator/impl/neomedia/directshow/DSCaptureDevice.class  �      �      �TkO�P~����6@E�6�އ0.b�1�x�L�Nf�zI[0�"�z��D������)-DE?l�M�����}�������_L��Щe3$���n�\.eKɹZӴ�`�rsѢ��ڣ�g/V�7�7����Uk:� ~CK��3��\u<�Z?4,"Ѫ�㺎���k��o���4솾��-j�/�j��v�a���}��k�e��f�O7-���±D�4��鑆��y��T�7��Ċ�5k��F�"S<ckKx+�)F@���Dcw�+l��x=���U����`)�UpBA��~��+m/0��l�w�)��/��S��Z�ZX�_��)/��s��e�5�(mOb�$�mc��F
��b��:����э�]`Itp�0�q���Hc�#��S\Pq�d�RA6�Q\N�cN��Wd�*�.�5���,;u:N}�\^�m�-7�>&�=B����h5(% ��(�p����I7����zn�f�A^��,�d���\�#f�q+�$�J�Sz0QF#
�(��p�m����a?	�M�#Y�}��J)������2�"�$Q�L&�*�oP�c���������NX�u�A�����"�0Dj�4WB�9A�B]M�nlQ:�r�_p�f�}-Ⱥ�c4����PK
    +Q�HC�L  �  A  net/java/sip/communicator/impl/neomedia/directshow/DSFormat.class  �            m�MS�P�OH
*�|�����!iT����
�b�H#C[�"�g�ld��U]���pt�?J=����������=���ܤ��|� ���aʺ��u+f����q� ���#rT�Ò����	d�)4,4.A��4�d�j��n�͎��FA]	S�4���L���3����ENҍ<i��{!,C��b5����b��ޓ�q�����+g{:����Z�xQX�aޛ		�8�u��$O����0��J�ȄV.�˅�r�Q��,�t2Ea�EA��ʥ��ѡ�����l2_�t�������!�����S��X����U�������$|�I~W�[�K[ݶӛ�³-g�P�ɪ"�swԍL*��v7�lfWuS;�j�ɤ��k�	w�%3����g���-��9����*���U0,A���B�����쮛���>�F�#i�f���#9O�F�N�A�I"��3>� �^�)�i��Y�$Lr�d�$B2O�P���qX�G��n�G���/���� ���d�1ۙ�Vf�`=�� 3$���gA��8�+ n�'�Ae��C�"���#ae�������"�*l5٘�d+�k��bT��z���C�:ނ2x�=�/�8 �2�R�F�a-�AA'�8���U���H	�	|��B��e�K�r�s�\qR^���;'�[�\Cͩ�z�EL�E<B9��<r�/�<J��'������~������`�0X����[)���~�!��"�3ȼ��a^c^g��3����e05�μżͼB�PK
    +Q�H����y    B  net/java/sip/communicator/impl/neomedia/directshow/DSManager.class        y      ���seǿo�6M� P�ł���%iU4��WZ[�6R݆K����n&��ܽ{�\z�.Lw�Xf�����_ϳi��p*Nf>�7�������� H�'F"������i��@o�s��<75�8�[,\Ѯ���ӹ1O��c��t���R1E^=�k+GEV��F���Rm)��jt��۲���f�p�d:M�1�T�k̟����j��a2N�M�N˘鄰#�����F�qu������r c�훬�ݾ��'y��s��Xx�H3w#�aZ����C5����u��.߬e���W̎�T�v�q�2˺k�T�Ѭ��a7�����E�m�Guf�kE�}%����W��n�U�E/��2[�-ٹg���(�3Q����&�ߡ3�R���<��K��;%�K��O�L$Fޮ		�$D�/!ΐ�013�0>f��S	}P%e|��ރ�p�1�x�1�8���1�8�8��E��0�8�H�`���s���/_12�lI�2.2�_3&�q��ǡ`1N�S�i�#ǘe�1�a�3�{���Xb,�#��+5�����yx:�y�@i������%PZi�O ����� �G�Ê��������>nyX�Q�p�G�C��m������M��Km��s�Q����n#�o�����7�Enx����-ɻɧd@-eQE�����ܻdo7�N��H';e�5�����A�c�GX�R��.�n�S-/�*OR�^\@��e0([x��):�I��[�.��X�c��&ނEjϻD��#�?ǬL���F^y��������'J�8����	�چ�)C�n��/��@\��U.G��:q~��p��|��W�9�>r��x��y�Fx(���KPK
    +Q�H�J ��  �  $  org/bridj/AbstractBridJRuntime.class  �      �      �V[WW݇L.L
5�(U����F�E��X�bo�0�`���	jo�b[{o��j]���]]����]�k���������L"	B�9����g�3���,�m�B`��'G\kt2�=��\����ߑ9۳��0���I}ZO�u{<yld�4�0�K��5��bX[%�@h�e[^�@ �2C�*��7ae�����)��l�����
4$�J�\s,M������eH�r%����@x��}��D����gM�{;[*�G�ޓֳd�P�\���a�����J�9�J'OrȆ�V����"�S����[v��m÷�w�c�=��P���C��H,��^��2-5�L#�Z�Ń3�Y���J��@Θ8jz�h��&��$48�:���4���|�S�	���FZw�r��3�P���*hcN����v�X[��D
#)PC*ݶ�x��eQ/��P�M��Hi�U<���i=�3�J�a'RQl�.�Z�S��ڞ8��U���$:������R5��2'�a�UT�)&e���ZƳ��O��.��YYb�z�O���G�s@�QB������9�챱�����-C^���4��ce�M�.cg�ָ�{9�nK%*��x��2�<#��c�e\��<�8;�Fc��/�ѣ8��+�v�b��sVz�d.WqBv�M=~��e}5%���-o��������LƴG��^@��yѷC8%�zN�1ѻ��<Þ�9�C�-�P��/�E)��@|1:~S�Ulƈ@�����W�v�\�`@����.
nX��(��n��\]S2mڔ��hq1��L3f�V1��,��G�3�� ��}Հapܴ��k��	:�o�f��U�kA�nA�6���)R��鋧�@�F�\6���W��*�Z�=a���7d�_"�%K���5P����N*�$���vg�r�Fr�)�a�ox����>���H��}����tג��r��}�m��F�h
;�狑p�@�{B��2^����?��:��\�<d�M�a�C��E!��(���%9���[�~�E>�+lr���QQx�c-V�w��()�.l�j%�8� �q��CE�#��Fm�����i�c�m4�<�W;�W�&�/��"��P�"�n����#nU��jyz���w(�2�
R�x(��vM���;�Z�~k;~�֎�����"?`7��5����吸�_!���<�H��$�]L�jJcS�����j���	�h�<v���y���MURj\�W_�-W�;�ZT�Ŵ�m��j������ѫĈ�\Vy�_7�v%ܳ?a��p��-ԟ��tc����-wh��8�;l�.���<~����?�A��#Ga2��؈1L L�u��$�Sziƻ����*�k԰���7��jp��?G�(ޡ�ԍ�
v����6_W%��G�CV�.�Q�R#�߸��4G�g.���(��G���{x�ҊS��5�*�����V����qU�8O���y��4��:�{��W~`��9�F'_�.��A<��8�^j�7��}�����8ٜ�-�~�^9I�;J��3��`�6��]��O�4�"����O������t�����O��v��6�6}�`�f �ĕ��hh�+�m�q����x�KytYa"��ܜ+��_�x�>R$�&S��w��*�{0@[/s�����F��`G��1�x�y2A�����,��Y��db���6��R�Q(�o��o�����.�|�ˇ�PK
    +Q�H���R�  N     org/bridj/AbstractIntegral.class  N      �      �TYs�d=�n�I[7ii��-xi��4dh��:��`�R�h�m�VF��-��KY��B� /e��CgX^x�G��z"��������s�O���/ .�)a���������ջvGm�e��ZՈB�pxS�Q�j��+���։"(a��{A�I�FO� -K�-�KK�VJ��a>H�\�Mݾ&!�^��$әZ	��a4��qp�v[�J8U�w~��Q��֪���U����j�v��81��Vϴ�-ma��mۺeF���U����=�h�R'd��(y�D]J����ۚ�֝OW����!��5��Y(�yVE^����p|��T�*S�1LJ�W,�E���֒��s(�.����1��wӲ��u��T춦覭t��p����pc�ѦpQ�+�|����v�.>D[o���dN'�8��2'���Ss��C�������"+mZ���l���QO5�>"��M�a�f���]��I�4�h�]�W�cd�%,�XD9�"��&ڒ��B���m�&YE��_���&!�Eܛx[��V�ښ�C��Q�V��aU��6�u��zW��6�I#�{<21|@��evm�|ڪ��#U��QS;�ʖ�	�D����Y���4�E��B
G�`L�Aj��pϱ�!SO I�!-����=ʞ�	G~p�T�c<�)��Z�A�Su��̕#�����>x؟!�p)�C����f�<�Opb�	N���T�L/��r��<�y�<E���_?s��G>b%����:��C,夼D�4)��\&��$�*�O����#�qe��t�^�uYX�S^�5/>�ŇE�7���P�<�u�p�������[_td(�L9�E���F�P"z��m+���������X���G��/�s�!���CDC_#�7��l#
x��Rw��)�ܭ5���7�m��:��>k��WA�m~��w��O�q���*�&OX'��q���>� �t�ݞ�}�C�ʆ��PK
    +Q�H�R&��      org/bridj/BridJ$1.class        �      �R]OA=Ӗn��|�PQD[�,�JC�ULŇ�oL�M�u�%�a�B ���_0Q��̴&�6���w��{ϙ;����� ��i"��&RXɣ��*Z3a���uw�5�w�]�t�r(��G`����~����)4���e����=7��|�	람"��b#�v+t;}��;LR<�j�%,-�+��|+�$v=���k&	��M�K��;(0P�T�Q��]�
l�V��Ԝ���e�|���2NB�o���{���E�����V�iǄ�΁�Б}���(
�$a�yꪱ�:kS��U=��^1��������<L��X�@��=ܷ0�'=vO5,]��T#�|��ύ��ƴ�$�	���8a�����A}i�<%x��lzA?�q�A
mV�_q��$`��5f��#�}�R�ΐnT? s����M�:Mk�o$����ciP5옣�"�ɲ0d ���jE�f�uiL�)�'�$y��:������E;���8h)%�W.�PK
    +Q�H��|�J  b  !  org/bridj/BridJ$CastingType.class  b      J      �Rao�P=
�ҍ	����TT`����	da�����$!��U,)ŔB�r,qF��g�����{J�M���=���^��_���� $�d�%#.㡂El�V��q�N Q���xޕ�A*wl�!TԻ�i7O?�'�۶�-��5�륎���y�ҞQ|�c��#X�]�o��[Få�)__nϱ�C�d����°�z� _�z��f*=�+;g�.��Q��s��->O���eȦJ-��k�n7���Ps.=G6R�4t��;&WIJ��6x�?9�7m�=`�O�v��R��Τ3+f���^Hɛ�@�a�����#���ϴy@s�J��4��&7��6�Pq�/G\��e<fH̐R�����"���(1D'1��ءX*=�v���P��1��7"�,7�L��vhii��
�P��r��U~F�@7��B�)�G�}��
ޏ�V)�E�'�X���_�����$��L��)�C6pS��(r�,��rfk����2�#�#8Ip����:�B�Ed�%
�H�P},���h�j� �J�7�B����y��}2��G���	m&`���PK
    +Q�H9���
  D    org/bridj/BridJ$Switch.class  D      �
      �W	\\�����#l�M�W�)�x��FX$�@X�k�����=��[�Y�Z���Z��Z�֦��U�x�ޭ��}��������{�&��ߏ���������'�{�q '�E5�ދ;��&��c؊�����ǰ���Ǉ��G$�G9��ON���~9���@�p�尟� �A��8�x���G�i����9l��q<���m��<�E�Oq|��3�,�6��q|��I	|���x��_���9\��p|��k�:����or|K��(q|��ߓ��9&9~��C�I���9~��4�O%�3�?���/%�+�)�_s�����N��s���������_%�7�K8���ǳ�ǥ���ǿ%�(��P�i���"�햗�`�z�y�I؆�.òT�ou�얶7���`X��������&C��V�3ڻ��{��MCY;d:S�?ZpiStvV��d��02��1��5��,�Fm���x°mZ��g8���2^�e�Y�j���gf<3K�:MW-�)�NˡR���vLvIj`�:�v��th��1�i�%�vhE�P4o����Hm1&�6�ȏ��YV~�uȤ�\�5݌c=��'|�P{jS2Ͱ��vedR�BZ���"l�D!K�SV��-�FMg�PN���}c'6�׮�O�Bư�ǒ���ʐ�:+oyg1����=����t��	�l�K{Ff�FQ�����(�i
������d)b���J��Y�%�M�pP^��؁��F����1�/�ֽ��"?�҅��1�,鿘Zn��5�IV�k4<�CQ�0,]���p=���0fخe!��Y5yEc&7��g�.��ҋ��^v��+p��7�JW��j\�p��fv�,;k:$�i����P�Mg������� ��N�Y?����c5$���b5�e���p����5뗏ڎ���#�ɎM�ǫ���([�F+W�-��'��	}R]v˛j�z�]��CC�Y�������ԑ��Pr`�k ��ب����N��r�n�^J�ޘ5�t�%Hr�RĒJŹU)����w09@w�c�12�́3"(�\}����+�Y�\3Wp�t�u�*��mR��:��p��G��d{Z֌�~��{zVU?}f�^����g���YԽ	S���Ly�r\ofۋ��H]��NV�g�+H��CG_����K{*������g�͞�ﯛ��oՆ���=A*m���J7�$�.�G!�.UD2#���L�'�NVDr�zLtzΤ2�Kһ�Vf���Mb"�9���0Y����	|ў������ԑ"�6��)&������t�P�g���TQ.Q�.��O9Y�<J�ҷ%�d��N$�*VM��KU��س�^��G����M���$=��T:�IS��n��f����Xp|h�)�fx(6P�P�T�)vHyK}y��=��|���6%G�z��NR����'�L�ͥ̓�t�1uY���4�b7�����e��Lo��u5LI5�}5�sz`w�@�`21��d�<��V�N�������7��F&cʞ�I7�)uv�c���~	$��/7J�"#��vW]^4#K:S�z��rt�(�'H������=��r�k}21�'U��W0J�uY�K�8i�M�ł���;��(Ć�'V��h],�i�����Q=�"�������J�o�"0�
�8u~�׵�^�n�$�R�w)	�����GtQ�� /:�ZȾ�!�i�t�d��U��A��-�S-����/I>��I�@^�$�!�F��c�|f.,A�P.UW��޴#_Cze3v!o��n!ы^�;�pZe7�����#�:i�B��0*���[@z�R��t��l��>#涒!KCC�|[����йԡ��(�<]���tv�4��1�6�-�Ͱ�%5f�ʽ�?_��~�l����6  Z趀:u���ɀn莀Ntg@/�%�TR,����W��(E�
�ՒƏ�]}W������]G_���2�~T=��>�bx��Ʈ%�]xk�*�Ԏ�7D�K����w�\��6�C��h�X;B���y���4T�Ac���ߏ�[�DĖ��V}D�{MCۋ�E�,S\,�a�3���P=���iě�����yyd�~�R�"[��E�݇Z�kXl���Ȱ���CʂS�S�%nP^�3�א�Iφ�L���^��4A�����(���? ���Cı�RA�z����a��Mʥ�"ߌ[���&��˻�Q����A,ޏ������h^�\,ۋj�\����Ǌ��2�ڏ�����G+���DںU[��s��qR�=RS�[q��{��dR�����!��W��qp�X���b�xUH4*�Ia��b�81$Z֪���X#N
��v��N���īC�5
[���rq�8#$�)�L����׉�!Ѯ�&�Q�)�aѥ�n��Gl�s�R���+�B�_�8����M
R�y�Zq���
�@���k�B�Q�E
4�ubTd�"�@S�c�Eb\L����-�����2=.�)=\]Fkz8R�)��hk�ü�3��q�:��M����26�>D����he\D���Ȣ2�� ���w N�밄�B#ۍu�z���e7b�	��͸���v�b��iv�ew�O�����a�Qy�nܮ�{�W%�~��.��/{PK
    +Q�H�\��>  ��    org/bridj/BridJ.class  ��      �>      �=	xT���.3���%�� ���AT��HA�I@�"�6$CIf�L�}�}��V�um5�@CWp�{�K��֥.ui]������͛�$b�_���zιg�w����)�*/�Px�"M^�.2�"S��@���Kdkb�tz�x�K��0�=DC]`�#5��İ�'��pM��}���Q���En�$ƤAX���8M���/�^]L��$'�J�^#
�F�ya�(N%���5q�.�P�Cuq�.��T/�И��4x=�k��G ������^1K��đ��z�Ӏ�����i����{�B�D-��+�՚��B����K�"z,��c�,$&ӣ�K�Kͱ��\F]��b�Km+uq������iN����I��M�L��X��zM4xE@�I�բ�:���A*���u�h���D�=��Ң�S5�Bb�.Q>Z�D�XO�^�Q��b�Q��i�q&=���ٺ8���s��<]�O�tq�..��E4�b]\B@\J�y���4q������պ��.~��k��Z]��@�N�{�fq��z��7��&M����[i��<��wT�==n����ǝ��.]�M�x�C�K��h��5��ؒ�*�V*uR�6Ml��?ꢋ����bg�+���إ�u��ح�=�x�h���(��}>�&��ӊӽ�1��jb�z�>����S�i]<��g��9]�����5��!VQ/Q�˺xE�������.����u����Mz�E�Y⯺x����;���.�A�w��.����u�}}���t�/]|��Ot�)�}���\��6A@~I����������+����;/d���s������~z�H��(A�L���Фԥ�,ݸ��t�}�:��C]��Lӥ��t]f�2S��z �&�葭�A46G��u9D�C��G�a�s�.G�r�.G�r�.su9F�c�y�.�{Y��@�'��]N�b�&�uY������
EA]�r K�QJ���q���)�<�އQ���Tz�J�Gx�tYF��9S��t9[�G�r�.�u9W���G��4~>*Yy��\���
e^.�ϣ�T��N�P���豘��c	=�t�T��h�V�r��-�+h�c5y�������x]�@'��$�>�~/r�.W{e�l@��te@�k�l��j����k����A�_^B���:z4�T
Q)L�*�J�=H��Vz�Q)��鳝J�Q�t*�A�3Q��Y�<[��h�\�������P(�h�G���&�c�V᏶C�K�[4WG��` :�]�b�Y}�����5�TZ�o���Sl�[�"8�6�u����5�Fk�����P���h�l
4B�3�Ñ��Ց`�)������@�Z�}�l�|���`�Q�o�u�{����?ì	�Ki��*ӁU28"�,�1������*C��V����^�cm�;�����k����Wd�Y0۹�\|.�F�ճ���p��\g��S��8���g�I�!4G�GԷE"�M�8{0�k��H��P��7����-3�Ե����L�g���b`$���"��<�D��fi�]\���5q�Av�Y��#��-��]+�{���MO+��*�&�k�K�2��O˒�]S��͔ V~���!����;�Z�k���� �H��X�p[�A��%���?J�I������(���J�Sۂ��)�X�oj®6�#!Ҷ����@SV��D­P��&܀�B��M�y�������y�6l�!�����8\����pc5B޴��Ԇ��*�t�nc B�'&���SR���a�?Ԡf��Ӫ�?ŐrV-���%�sV#�c��IU)�QJ��ЀZ$�7Yse�j�������D�+?H}�<}Fl�����G�D�ít�5��@K ��+5��5#"|�yP�K��2ԋ�J�#S4#�#�!��=p��s�a�F�[g3y���
�T���P���yu ����2JS-G�@�V�l]�Ւ���O,Z�`x^_����fP�sh_}�3�i�$�����P�R�Yq�T7M����p�Q���%��}50�����%@2�Y�t)1�̥e}*�<쒯�e�����"����@�H��'�E߾���4B	�I��;��A��V��-$=$�Q"�҈�W�*�mc1�Q)?#�7wk�_�a��`B�m���+��k��C�k�*#�4�0�Z׆I������)�_G����M���v^`�,"6�A%1�f�8����&��@0*i����I=��3�I��)���P�ieM/@IZ/�?�-9|(��mZ��c-WЄΉC|.W�r�%�8C��KZxx4к�2;��+����?�r�-�K���f.ꇳb4���s����;�j=��p�IC-��`�S���$�W�Ⱥf�7��� g��^ɘ�r7�{0��"A�Zb�d�@�zg�1�_,P�Dm��,�~�O�@�Qĺ��@�,��&�\�U5�	�&M�h�d�I� �/��	�����I}��v�:K��� �k��ԥ�`l���]�M�J��F�%��E�%�⏝~asJZ����B?��?p?{sL��dSE)oԖ顨),��n�Ⱥ0���S$n�I��ERZ�%jW�1❹����ISY���f�!���Zˣ�1>�?*�CZ�s�$M�o4�7 )RQ�7�&�A3�Ǥ}R�U�6�Ԡ�p��P���b��C���[��xXW��ג��}�\T��փR��o��k��2����[��E1����of���Cv�Ai�J��б�v�����)��B_�%)cUP�] ���w�?�,�.ހ��^���l\�){i�BM^�ɋ5y�&&`��~IM<L%W$UTJm��m2������]nkj�9��=1�a�����/ ���M�a��7��)H�#1�@A����D"a�F�� ΀Z��������f�ЭH��޹"4k����ρ�KL�1��j�^��ަȑ03Q��]�Ĵ�&��`��U�����ؼ*"k��Ž�(�M�"{3����+C�Q�B��(����y���ă�6!6~�RM���v�_AV��:���fX6�)9�� kT�7#1ū�}J^b%uךbf��
~Ջ3*#C�^�=�ɵ*˓n��"@c�'�I�IR�3�	�b�u�H+�ǪI���U�g@R%sL,����t�����5X�S�_D:�{��AJ��P`#bŃ�v�B�j%E&��S�0�L^�}hډ����h:��I��+U�~ǰ�e✔'C��ͷlBxP�&wK������Z=#.g���n���$X�D�Фd�y��k5~��J��Mİ[��ːvk��b~Jd��و�BE�|� =�c̜�9�N�hb'���]k���%y�ݘa���5���6T���ˑ�9�<���D���sDn&A��Wf۸>9ʩG���Ô���7(���%+�ڦ���W-r�����*�'*_�w��9t`r�����ZU�&�.	F��N��RT˼�}E؋Sb޷�a��g�4������@z�7 "��E/�0Ir�A����o/�Y?��:����u�ͫ�Ms����m֐õ�9�!Ќ�4U�L��f_���FM:�!q%�i��;���Wr��ǐgُ���|�4:\�剬�򧏲�;�+�;��;u�Tb�쟫�iL��v�`p���J���Kӈ>V/�s��>F��ce�U��
��PC�B#��v��sEI�r��
�@u�j�����)B-z����&.�!l,Ǿ��@�>\�Ţ~�R�KQ�'��pf���l�Q���À��&�D�	�Iϒ �����/�F\&����b]�+�� :(�D����^��Ilii#5�e��Abdi�/}�jr�&1v�g�7�C,M^�Vn��L��U�QBsl{R��0���<ߐ�b�i�C^+��ً�y��ސ��v�,�t
�P��niBMJ,��S�
gT�df�n~S�������~��I��ֆ#�/#^c�0�q��zV�����m���������I�)o0؟�o0Ĉ�C�Uj���}t��SZZǶ�8��,��˔��m�և�q��tJ�^�K��k���y�
�f�1~�!o���zv�!o�����y��Ð�N��Aᦦ@�������e!��<�<�P�܅�K*� @��]���Mc���m��ǐ��{y{2a��5y�Ę���pn[4���)W���!YnYn���Zn,'���F�+/�(�EEe48^��|~�Mn1�Vy3>�6�[�fCv�m��.�h���$tg���������,I*�&��6��q��٭ɝ�|@�2��7�|А��1��'��G�6��<Ӑ�����n��w�Q|�|�!���vv���Sn�5�Tl+֠�̵�=r>��2����8t�a�����̳Y�����$��]�m�[�	ﴔ�|�V_�4�hr�3�|-2FN�dm���ȼ4�k�iC>#�5�h���~�,�K���bX�(�C-��b�?��q���vA?�'�|L���Э��@�!_�/�e��&/4�+�UC��>^3�_��|C�iȷ�_5y�!�f���ŀd�E�hyO2��hoޑ���=��j��%+�w�
%�y��+k�U�VTU�)9W��\ۃ�p�|����I=≖g�X�?���X��D3�C�����O��&/1�����r+�Kp�;Ӑ^��7Ɏ-�b�����
�������f57��vyՒE�5��KOZ^�������\�>� 7?��k���1/ZC~,?1�6��`��;v=�Ⱥ���%M~j��3���o���~���=��'�c?���A~�3P�I�۬2i(�<d�F�W���v9qÐ>��_������ꝑhM�_ .E��R~�����kC~#�e0|i���G9@�Ԑ�sQ��'��a�M"����q�I�?C���+5�w�IC~��K��/�4��`� 0g�b�3��{�=`���d��D6R�2�s���؆�~��>��h�sy$�o�ViVB��y1�=iq����f8oeR�+�KIV��J(4��4&'�*Y�&4"�7��J����T=<jʵ*�#VC����}�t()�bdj�(.F|�a�8t���T'�Nå*��Jk�X6\�XV+Fvj�X�^W)�P�Kۢ���ʈ,���f�0��n�Y�&9�}{���ǣ�1M^n�4�����������J7\$vF^^ّǗ�P�_�o�2]�@R4���q��L�ws��Hq�oRn0������@梄2��w$`;�MI��Dhhנ��@���"ax�`�&��n�����\ɯ"w5^G�N���S��$�OyX���^�|�܃([�A4g�kp��d����`�b+`b@8F�K�d�Ԙ��$�}D�����ߋp�W`0{��q$��ghȵR?XZcu�N�=t�J�ڱ���K�c����C�Y�wciyKKS�^���@d}�>-YkN�ŃpD,���=9r�Oz��0�(�p�8Q���#�z�6�:��t8s�(Ws�4\�\���k�ry��CZ�>z��6�X�{��a!����e;�w����d���g5��5�5�p��g\W>"Uߧ�8�I��dѶz�Gݽ�vӋ�ߗ�K��P��ܼ5�Z5S>�y4gu��>ɜvR/$��]�5�]î���9�U�*2��{�6{�>����U�%���?e�����?���K|����fvp���I��uc+m幆k2jo�!&T�!EItM�g���--�}8ԅ
�i�'>�J��C��k��:�5�p��f�rmj�-���2I����Q�qb|��.:|.�2�j>X�k6��ґT��Js�K9=�ң�y�YI�[�s>��R�(*uRiǸ�s��<ҋǯN�b������_ ��vKB�h������:�u�	���ǫ�>l��}$�l��P��؟��Ţ���-v�{�	T��1��ZZ0Z8�F��f4�J8JE}�t�p>�
zc�5Օ�>�51j��(e�A3K�p�5}F��9��F�`Oq��
�(-GcӨ4��R�<寮�ʤl�Ͼ@!�����B__��/��Xt1(��\����;o�ÅtxB�
�z��x�P�|!�ϕ:-��JHl��>E���t��{�I��(������Hr3Q˾4U����H����*/a���9�����ԍ���4�E�	�uv�TFQ�������B�6+��ǸTx�2Pe� 1>[�ȘD�jn1�!�'%$���8#!~3C��K�g����ty��6\��
�~R�[�����$9	��~�DA�DYM��_���х���1�n��� J�(AHq�����%�B��M���c��씿�J6T��pG%o��ѱv��%V��8[�	7���b��)O)sI	ە��T�ꍉ9H�e7֧�i�5o�Q��-���hq�N(��Аt�Sut�(Zo�s�T,�"�������/�����AIl4o��A����[���Gk���C�U�E���kv:�5�����aP�ЄY�-���T��Ll�D�-�5�L�&��ʨb͍���L�C�n��� d�:b��=h�ꕙF�`h
�ƺ�Vҷ�N}�MV��_��r�l9�F~ʻ6�(Ɲ��1 )�Cg���������8���7���&�s"Wn"YPx�:����3��ɬ���
�zb��-~�E�%�I}L��5��Eu�"���Pp���z�\u�H"��6�t�i6%G��B��u�&�����#�)��5�\�C��Z�.pj[ �a��o�H�a��6F�m-��U)}9]���"�My��J��1L'S���~\ʔ���p![���/�T(�ō��Ig�q���ݿ
�*�6�p@^�.��K����� +�K��9sfE�N�	��w$DʍBѦ�J�?0���%��:�d0,��+ZVH�c�~�W�J)�Չ���1�������(��sv��X�Xm-�")����H�
�L���#ܤ���ӄI3�� �$����F?����%�O5�b
�����)<��u�%�Ƶ�u~*�S�����"��z�
U�=�`̅^Lrՠ�֢�����<���,M!�*C4��Y �9�$�.��&��z$]QHb��{ �^)� ݢ@EA�G�?�Θ��3�yI?����g��~Fm�\�X?���FMg�0K��tZy��ҸrE����Kj�j��1p=� ��P:�Ʈ��O�]�߿p|_�߿t|�
�����P:������ߛA��V���0��S��q�[�o���9�>:fŲ��V�}����z�m����Z��������{���j�;�{�~�_�D�^��G7��d�߻������w�������H��0:lP�<�@g��X�º}�I|>�_���_ W�`[Uק��V���|f�,{��'��9��8�=V�����f�v���,~�q�:A���,�*z��U�4*��NŌ�qhV���������� �������=L}�\���F��e��#v�(;a4���r�5�.�r�]��e��	�D|u�������+��j��S�D=
Y�
ára=L�P�h��p̄ӡ΀8����8�p4ù8�yX{>�l����.�[�"��Pdl����^$��n�{	��Er��U���Ꝺ�4�Z���M�_6Ԁ|��:n�e�� [��鄂��P��(��`��a��un��06;���`o����bu@c����n���p�w�w"��V�	�������]Pb���^����}��,��C�n�GAk��`��~�V��6,����� �PP�*L�P�3��~���c�p��Ђ����#,��������޳�bNKC�:���T����b�n���:$%��S���޷��[$���G �wA���]�A:qe����D�Y](�fu��n8������'�#�
M�-�s�l�E��8��(V ^|�4xA{)�{<
���ۋ=G�}��>vW���ǖ��!��P7}�����!�c������"1��>�a��>��"Ƿ�>���@�~ξ�� *���eeUtü���*�Ph�Ǚӫz�����`�,�%GK��W�?	�Im�ō��X[r�=����}g�=C̓f���CU,섣oMv��&�b.���0�=�d?��l�R�?����w�1���O�Ow�,�:���E�``'ԌB��Zd�L뫨��jKK������k,��{G+��Fs@&�2bg�~�Z�J3��9�s���ȇ#84S���-I��萅4kA/].2qb����;�&Wm1bq�
d�
�L�$���|.T^u�ܝ�t3���2Kk�t��>w���d�
���L:e�X���V��$2e��]߃��jX��C�vk)�ݦ�DQGo��N�h�]0����i(:J��Y,ei����2�K@GQ��5�#�c�P:g�=/Dj�!�ݰ�)9��:�<]����0U��3��^h��@K�سe�f�]s[sd+����?�� zP]j���`���P��4>�@
�t�)�m��pk�Q��H>�b�s�^o��U�ŴQE;�8[�.Gb�m%��h��d#��sy�KW�25�sf��^c�������Zd1����Vu��qu�X��2�i�1ApȀǤ���x���z�����ɧ���"oYv��N@�?���IՅ�`:U ϟ��+�M���,�����P���a�mF�����t6��0���$6	�XŊl���!O���+��3ynsl��B����W����h^CvS\5�¸)P�6���w�����@<����0��f5�{!]2j:��UQS�	�ǳ�����T�L6F�(��~�8eшsx)��� �
���c`��C,h �Fi|
"c�C��b[Ųp�L�;a���G�ioXj�y�^6������"s�:a�fȏmX0�aY��.��y�֊
CuV��O�A@ݰ
�'�Г��a��Qh@6��!l!��P�ja
[ǲ%p<��	37�� p�����MbلQ���j{�r��a���ḭ=$j���u�Td��m�~J��	2�X9Q^WS�{��*s��� �(GN!mO��&�:z>� /9�M
�nrn=z�B r����R��l��`.��4D�v��\�3��5{�j��!�كn���\����ǧ�2�'-����5sؚ�]�kA�NE�"�ݩ�]b�!%v�l��ݴ�����&��݋��	��5��B��õ��0�(T�V-5�,^\Dl[d�m1��%hIK�p=��Ld۳�m�A��\(`�C	�d���l��Ą�+A��LP�f�9��EZ�t1�PxN��rDsn�=c���n�-(��m�Q�G�[9����k;DwB+��Tn3�js_��a�N��0,�Ƞ���`3��pCҝNN�]p����N8�c����5�?��QO�ǹ���b:�<T>I�|U�M�qALo\�B��蹲.ꂋi�Kbk__�2s��/w�}E�����U���VXCj��~��+�����.1՝���ȧ�'s�S�s����.�����9��F��\lM��+a��������C5�$���<l��ܳ�=g������"Fܯ�u(7������eo�S蘾��{�}�ށ� ��{̃^Y6�ݖ���	��>e��3V��͎�`�X��b�q��e�a7����N�D��W��Z��y1Ix�.� m<�W"�Fa�꧱c����G��_���,��/�C\��G�;,{Ea�Qm�����X�w9d���ti�V�YdJx������x?bpf�A�~pk�GE�&O��a�%����Q^=��/����V�HG]��mpM<,V�� e��|_��+���K�'���ko�!��� ���knuDN=���#�9�n��yt;ܚ6X�c'\�2��G�����uX�Y�����y�������l�ʚk���� 7$�s|�*7?����ѳb�c'�����&O0<�s4' ��~"]�e�ۀTY�d`@t��6@ϛ�F0r��c�e�����q��R�wc2xS�w���W�?~��Ԁܔ<OIJ@N>x@����~o`M�h9�Ь߬(��P�}���[E��h|9����� ��Dk؃�Z<�ܥz�`-:��~hL�ޖ�&��l��G:h2��|��F�ֲ�'c�ʠ "��F�Zǘ��[���-Ih��$���2?!��*'#����Yj������x��m�!s]>�(��	w�������YS��G��.���pw��{��n���$�����1@_	���]��n�R����a�����>�Ͻ�����vB'�2ͧYֶ�J���Q�8��md�t25�M�{B��n�O2�ϳ����{Tw�(J�u�\�xt�3�B�rx�*��"�FES�Qc�0�/�I|1z5����{����mW!��J؄Z�R�-��;��'���!�~���Kd��Z��Rƭ��&X�[��to�S�$0,�3�(�t8<ɣ���Ep?oŒ7���׫�ﱶ>W0�>�_�#w�#w�/GlQ	�� òyC�Ѷ�ގ����� ,{���lQ9�}�O�"���(g.y�t;�z���Q!K�d�t®�� �Z18����A��wб��T?��c�����
�x�䩐ƣP�[a2o��a=����1`jG�}�-tE B�|?����{t����L�+�9�.����h��ݚ$�g!���Lr��%��?V*+��,���{ӊ��^qWl�sE$H����ኗ8W���:�I��C;��Ϸq,��Wf'<�+>�bɶ�I)s~��_���ڡ�2�&���~_d)��q:Ң� �6�(	�ŽV<k>��[P�O��Dut��A�v-n诡�_��١��!��?V�G��L�R�]��T���d� З���$���9@�����	��������l��[)�ɨ����Nx�-�=7�W�nyd�)�n%h��J7�)9�GY����.��wC6�|�>���|j��<&�xLV�3d�q�r~E�x`$���Gؘ�ѯ�LLĹH	�<�Nxb��A�?�L�I3��23��R�s�⟺�yz�`�_��/u���~�z���]��ʬ?�&�׎�J�.���x��0��77��n{+��ټnx{3�Y� W�;k�}3���@��zN_)�ޭ[)�ޫ� C����)�-�=U���W���9�)en�ɺ�}��V�M+�&~H��`#k��W�&�_78��+~��k���mP��l�Ik�5��)ڲ�/~/~j�ݯ.��~Qa��װ��a����>S����o�)z^ġq�|�D��ѩ�#�][쀉�e���wA95�Cp�+���G �E�������$������ix�?o����K�/��;�?�j��,���.�a��:���������-�7��ξ������������G��X����-�C�J�_�rԠ���~��$����P�+�#.�k�>���kQ�1���:R�1ٲڮ��z%��[Ќ ��F�sJZzh��QV�4�cƄk���Y�Cn̒�a����b������q�J����c�Q�/�*�o�ǰl��o�r��7�3�m���:ዘwy/�]S�%�+k̥�)��p�Q��ͥ2���B��B����Si0U�;4�4�i�&KS�Q{�5�Y����=�	�GWg ��o�Zp������d��I��0Q�Ǚ�^D>�B�PE[Nߊc5����X��a��(#�R��Z,/c�C�2�NnS��`�x.�C�"���s��A M< o�~K:�~�j�|#�LsO0��OuFU�t�r���02�Pv�����EC����r|�.;z����E1�(t��� Q�D�S��hi2�`��"�ϡw�5�ʮ܅%����[���A#e�gi��2�ù�FBS�=��b�zm�t��܅h잪���O�~��i9�)e�b�Q,K�u��h�}i&~�>�^Hj���i>o�{�1]n��������mQv��F;�� 1��Ca�8r��0]L�r1������/�  f@���Hhs`��������݇�袙�I��H���^������<*mQ�N���?�����=�R0�6�!ʄ�o'�Q�,W��T���� Mq Ww�oAC�p�'م�դx3NG�wy��@'������l<R�N~c9�lfD<!�1|bO�<b�a�
Y���Mt3W �m�-|�xO�=����aj����nZ�� D��~�ˏ~4�����	,�Qoss�"c��)j�-��!��'��h�7gԈc�qn�*X#��Fq\*N��E�Iϡ&�*	��Pa���Ԁ���l�9��y�g�\v�H�U�e5W�=�`�����@kf����Y�����5��~.z���"$�Vud(:���N�\��7�K�ibMȤ�M>��G���Ň�\��*��P�����qʫ�0�<�$��6��H.ώ��&J,��u���[Jg��WU&e;D�ҩ�F"p�hu@[nA;ƚNi܁>�H�,�`�;�'����6"p��i�?8�~�o���W��Ĺ��ѵ����{iٛ�n�ތ|�ʹ.�S6�y��ҋ���41E����L��
P`,s���(��b��0��tr��B�ݔa�y�,ӤA��� U3�:b���b3���x��JVb��sw�,R�{a�O���^��ӻX�fȢ��-e��tÍ+��`�!�Slp�ؐ�����ge{l8訄 ��<& l�,@�>/�������i�覢�3�ذ�Y_�^���ͩ�}��Z@%k�5,͗�v�H�+y�/Y�\�B���Ȱ�4�^�����eXs�L%k�L�/ݗ��F����+�̙�� �P�#	�LE�QT�}���F��U�o-H���"9��҉��Q�ϥn�d�\b�٘��.�,��E��f�v���AwO���i9i9�۠���I�R��(a�·̍�`���xe)	}���ރ���UٖMih\��f����t�y�}Ώ��^+�P�9��@�>�Iz�gKǏ��b�+Q��Y�VB�~`(,��LYW|w�O��,�t��檀4]����|+6A�� f�a���Ka��V�_�]���/a�����w�u�������o�72�����!�wl���Dkw�M�.v���m���Ľ�	q{R��=#���E'{Glc�۹䙢��;��͗��2�?A<�O{����O�x�G�3|�x�_-���K���&^��W���u���3�R�ƿ��a{���p��E�xG*�s�{�B�/�������0�y]��`:dgc����GP��e�
�(��jU]&{ڔK���Zc�Y;|��~il|�f1X�yU
����3Q]:�26�
��@
��wq�H�jl ��GWGk���oT�0ٷe��M�Hd���� �����|/��I��˱$c״�yw�z6������2]R�c�L3QJ��4���ɂK;J)TNo2��?�@mtb׃K�j�t��>��Og{�{Х�$u��X�94Ͼ�A�3�%ݍ2��s�Xe�������}�

� ���V�`�S��
�OH��~��Us��7,R'���@&�{M �:2��$�β�XW0k:Y�>��d���C6�'Ȧ�=�d��`�(v�ö�Rug��'W���Z�M����������o`����P���G�a��>şN>#f����4��H8#}F�^�Q��2s�X���{̦9�R���p��G��V��!��
��)��r(�>��0J�qĵ�x/��(��c�J�(�M��Ny<���X�<cp)tX��#���ݬ�B�9�l:C3�|��ѿ(P�@�/
��1b�f:��X�o��{<;�,t�xx���%���l6۶�G���d�Qi�]���Xg�{�9w�1��V�����(�S�G��B��=��$8��@�e��*���l�n��0@b$+a�,�\Y�e	̔�p��
��48Y��2x_΂O�l6H���r��b�<r]�����{��yw���� M�@q�Ji/{0n�1����a&����U-�juD�ރ���7Q�e��R:�i7`��8�q^�/Y�q�u�C�w��LΓ�P�&]�G�KV;��Ahp��L~
_oy�e\0��Xiz�/�W���[��3�Y�}ǐU&�[��$�%<�U��5�f�.�?r�)����E�#���Q]l>�wًރ����6��t�\	c�q�'WA�<&��Py������_Ww}3����e^�����u�T���M�C�_�lcG%+�zT
	��1l塿0Ϛ`�uqBv��l�Q#���;�����;�yA5�����`'��P[TL7�e�O��-�I�=�;n�*jnlxe3d���0��-0I�� <̜[]�����F?�ALFY��`��]K�t��`-�J�����l{�y1���R��X���;�A�{��El'��oH�����]�s
n�Y��C+��ir=��(�a�l�RyZ,iKkX8`���ӭc��w��
/�Vs�u]|�^.d�
/�}Ȝ�=u�S�0V�w v�K�}+ǒn��W90�z	��"��n�K�LՊ�v�hݬc(��0�S��<�1�`�$$���3�g!	�u���Hy.���A����0K^�E�kL@lrT��vE�*��E�y69f[� ��G�_�6�a�0&�q�%0�w�͚Y�X̳Hd��t��S���ˍ��#˴��l!��bI���e�_3��;�����y5�,�{"�o��Q��2���1
���5(�:�2z�eXk�W�����X�&\�柹��E�~��H�:�TNzWoR�)������fr�_Tba	Yz/���N����2~b,��.�Cj������~7�c��n�b_s���k�M�Iު���2�_��u�\�4�|���V�{�aXX#f�*GR�݂��"o6[��u�T�I��S�g<H:���]K��b�U[d�*�uс[��cc~��;��2�Rv��+�İ,�
*�ia�04�(.=����Ӳى���ʼ>��KN���k��ءҩ9���Fu1G���^�/�P�X="��3�7�5� �w�@��k�u�5��5nE�mC��tG�g������H�W���wn*���|��n�
{��y����|�8,By����'��l����YxE>����u�'��|���#�|&_�/���|��y���@�6X�Άɿ���6J���ʷ�D���+��a��=���(��[����V���Nee�p6��~dCT��G��U~ �+��F��C�}t*���g1]0�1ӝ��p�`���o营P;]A��F�~��OU#�応	i=8�K�S�C���0Y� M�i�T����u�Q��զ	�J�z��Qp'�����(cO�bժ~��c��ݳ�_j)gr�.�v��wإ��Ү]�,�C7î[c�
v�&,5ola)�j���R���t�S1\�K;Y�
,��ZU��������dm��n���6�k�=�,��n ���������d��^�v���tSb�3:ٙ�ph';K��d�¹��<U8_y���&:�7�U��l�}��1����v�lvA7��_�U=q��<�g A��S����4���S 3�M��/`1Ǳ����F���oQ1|��a3�n�@z��d�Et����{�3��s�/p�K��/e#��ȍ�C�wl��`�b,����u��j1���?@�\Mh�]����.�)��]׳��e���2|7)3�CNb�s{�*�����[|��PK
    +Q�H�'��Q  �  %  org/bridj/BridJRuntime$TypeInfo.class  �      Q      �T�NA>C���T+Т�Zu���!$J$)!`h�^mw��4ۙ:;E�y��P�3۲]�.1��s�s���?}� ;����]�-�۳����Ő+֧��h@�# ��7�S♭�=o����O{��my6�Z��Y�i�h���X��o�A w]��c����)�`\Q�_K*�@�q���o����D�}��q)��Jth|�{&��p���(9�ڊ^P5���}es+��7��q<�����F�suZБs&Ts8�����C�	n�=Y���f�.c��Ӧ	$�x���6]7�<�={�2�?���$��lI�˿A ����;Rf����m�1OW�H�Fq놹N�k*�x�*���E\�{,E�:C��Q4\K�u]I}�@�ɺ��@�j�i�Z3k�����s�h[��e�q�B�k̞���5���8�����z|)�=R�b(z�<ln��9�G��������_�
��!��<,����?���@�4�/o!�%���Q�<��Ѳ���Ke���=-�`=�/o�f�{8��<�N�����i��]HM��o^�[ =����PK
    +Q�HX`+Vx  �    org/bridj/BridJRuntime.class  �      x      �R�N�@�H���|�p�4�ѥm�Ĥ���ƅ����S�����𣌷���G��;=��s����� ��J��z����c_9���m(��$ J}:��C��\w��
$H(O�"����/��=W�,��WF@�YeNj�I�����zkBﱞ�gJT�b'����G�ZK���ȡ�@#ҡ5����4��l���P�W;�Y�Ԏ�`����uЇt�~���VR�~@�����i�n\.p"5y�Ym�mn�r=h�i����m�LSՑ�9�v����X�C�_[����m7�,v��[(B0/0�d z�:2 ��<�+�
6��J�+��-�˰��ac|��k'�-�.F�H���OPK
    +Q�Hj�s�  L    org/bridj/CLong.class  L      �      �R[oA=C�\���B�U�w��ҋ�Rk�ZC%�%�/f�S��v7.K���3|��k} ��������+��l2;9�3�;�����'�E<`��j�l��l�2�~0��6�)��W��鈪�?�B�t��qo1����5a��(	��[���[��������0���'��(i�0�'p���x��N��wč�`�_;�����P<��0D�����!��U��*:�nVeY"/ݧnVSM4�ag���T��k�YkWh�AD�1�/^ֹA6��v�| *N:���.��K�W�U#�V�l�R�)�dC�5�%/A��wڇ�f1'�3�}��!�y�H�u�IӰ�4|��Պ�&N�%rԎ���=�>��z�����%5��\�f-��p�!�LD�eU�9�5u�T.4Hy���ò�]$T��vElꆠY�%�:%ߍv� �{
a��4����!���d������>���'a�j7�T�iRgK�Q'q������=�䇖���\�u�%�ۤw
�]�2UH��x��40��K �t
��9H�@ʽܗl�\7��s��gZ�;�续�'����Va%g��f�FxW��:4�-�����L����`��@d��>7/}���7��dG�x��I�)�c�&��u$'*�$}� PK
    +Q�H��뚞  �    org/bridj/CRuntime$1.class  �      �      �TmsW~�faK"nLҤ/b�u�*���61j0Qc�}]��t�e.Kl����t,ft���L�����sa-!A�0\.�����<����GO �A0�e=[����ͭ��@��9�!�io�Y���٫�M�:Ff��k��.S���v�K�0��B9��3�{�uD&����~��r��Vl���V��
~U�^͟/�I^s�R��[�ϧ�{H��a�]��{,:���83[��j�^����0� <,2D�Bz#��Ǡ� È����2�49�b�*�p�A��(�b���`��?^����CҰ�+�z�Fح8"�G8�0�W�H�՗�­��>1�R�fV$�dH:���f+ŧ���lr��p�*��"-_O�ZH��]7{��?7?S7�Q�+�*/|/H���3I#E��vBCY����rC�w��	l��0�/��7{����/�����������K�_㔁�p�47��j�ۙ�a�9�8K�#y�%��]���5�F_
{K�!�⥣X�̬��t�Dsط�-���ÛJ>�U#$jB�N)�E� �)���kW��MC��	퐒������x�{W�����k]���~�
�y�2L��g�+�-L������b!�Hՙ2UD?�W)S��S�o�R(�e�м��W۷+\�'S�n����XI�=;hK���_EA��Q����+����9��"�zoC<�y\�\���-���$�A�DB=-�k�51A�?��$F���`2�����ش�ɇ,��,�V�;�N�?i}��B��"(�k���]�}��͇8l������'��Nn�s�\���+�t����]�`m��q�."�20�����.��^����������Iu�#��Y�	�/�jϰ�=�%���K�i��M�n���Q��b���
�ucQBǾ�ؿPK
    +Q�H��T�  #  "  org/bridj/CRuntime$CTypeInfo.class  #      �      �X|S�u��eYB6`�1l�� K���	L�
��`�$��,]%��r%A�5}��u}��u��_c]ӕ�X�Җ�/��k�=�&ۺv�֮]�e]�n��?�^]]IWI~��������?���_~�s �U�V���ȴ�N�12v��-����������~(���S�&*T��B��v`�-Y�1qG�Tb$��Ύ�K.��|�-3-��>55�cTaI�I?Z����
�e���Bg�~�"
�ތ�)�U�Z
|U�q�eh3�"��X&��+,u��K��]++ܖ/�d!~@a��H��Ua���قf�r���2iz���"�D�`ck-�L�7U+�������ta��Hċ�����ЋU4�O�9"߫�!,����
�b!�9�Gޏ���Zc,�PL�eCX�H�`(���1�*ח���E���l����c�X��kB�� 6���a�Ⱦ�����I�5u'�p�H�
i=ˣ[pC�GoTX��~lU�MәT�b�mخ��&l�����4cZ�S1u[7cW ;�[��J5��DAK���L�F���4�0��jn	�
�{~<���[�r�y����!�	���I��IK��̤nɈg-uB�ľ �`���ؗ����nQM3�x~���h'���y><���p:n�#3��iٔ���,.U�QŘJ�1���XA�6��Q���C��K��P��#s��i-\8�͇Ok��]_��d&ah�p"��3�dx�P^Ȉ�4`�b�2Ւ6K�r/�h�$RA��^��Hq?f�|��!�R!1��$��+$f34��^�Fcc�0���œ9)�,$
U��)���)�����wkf����Rΐ�9��N���K��]�_i�|��VU�-���R�����$�����U��d�;�]�lqN�nyIR���
�S�C��z!\0���>.;��j�a�N�&�{���� G�K�܍�I��*�ܪ���+��{�ꣂ1�&�9�7�>���m?�J��f��(��v�#���Ki��6���5x��ԙED�O�s9�ϳ�k�Y.»�1�{�CZ�d$�x�H�ߏ��T2<�(f�5n����S���[Uj���4�J��x5��V{�=g��nȩ������iY�t�j|5诈���'�k��z��*�]�`�-����T5��0ɤ�ϻ�X��mϞғ&é�A�\.���h�Z?D�jL��evt�[ѵ���Z��Y|.����e�1=k�\�!�s{����:D������l�OI�ǗX��쿦)���l��&iė�
�0��[�?�3_��I��O��\���F1A�5v��ӹR(�I"k�ڨ�i���l���8�*�\1�!|�%��̓�4�Ȱ+(l|&�K�?�'��_1)*��duI��)�t���E��=�s�ۚ��]��w�����0,�ǰ>�[��=�
���Z�:i���e�c����B�a4�rY��8��
E�dN��jh2�>?��3Ѹ�7��S��n���c���.�|Z,�J�ۚ+���i��$�M��O���7����e�ɭ��ϭ���2�����L�R)�1+��>3_r��Z^j��Wd�������/����Y�`T�3�ʹ˥��}Z3��F���sy�e<�Gլ|T\���*�O&�)�m�y���rˌgǊ�����E2��T����X"��N$J3���W�l�`�|61�N��I3Q�Z�<9VN�c�d-s����u�.v2��!Ĳ�V�9���Ȯ��ɯ��
��Ss���MܫKb�^&�Z�H�ҭ4�I��9ݘ7��k��ґaR�R������o�GX!�FȚ/��+��d��\N7x�;�ӌ���x�~�ԁ=��\F��5l�|��;��mj}P]#�g�k#Λ��h�,#��eH��·���x�����H�I���`��Z�fR/.��R�:k�MV�tʪ�f�E<pg\)R"O׷*������m
k]S�z�y�=���9��)ߴ��M�ϪQ0tFQ�pz6�`��)aLO�s���9�0�R����]�H����4U���{%am�_��8�tkO��Y�bAǺ��/2d�61�Z���Q���Qu�&�W�[�}�<�w��m����3㬄��!�0y�9��g*<��$;�1�fY��HZk�"}��Њe�[ ��J��	]�^���:/��z��_�[�D�׌���o5�pg��D3� ������u��F�/!���h���~�6�u�O~.�%��I��Ũ�}�CدpC��ź�8t�"w)�8Y�:_�G	ӗ0sLXo��;0)%�� �4�[��&d���`���Mj��!*`��u+�7b�9p:��͝u<9�"��)D��y)�����y��U� �R��[��1�q�%j��%|�Kx���:>�Ư�0�j[u�e���ø�^!_A�e�{����W�����Ehe���?����_	�|��X;�هߦՕ�v?�,+U������|C����f�}�����7��;q�
�<�{��R��F�����ЯR����>*�~*�!*�a*w��}�V.�s�G�p��/��#���5��_] |�OV^v�φ��Ƚ�6������"��]E��P��<�����j��UuBV��t���D=Ĭ�l�d/��"D>"��̐�F�%|z�����x�������3%|qrCK	_��/_	,[�⣬v�l$Q�_���5<Jy,D������� ��,We�Z�_7�ElG[TF*��KW��e}�|��S_dq���gj�#�Dq/.ٚM۟�/ls.���J;�?:L��z�������r������|'Z��5l�"~p�4����KU�̨m"�U�'SխNLo���U�6+|��e��s��|�ϯ��|�R%�oت���I�*�\9?"�LD	�Ǳ�nM~R�@�Q`Ux̕�>ƃ�v���P��"ɂ�w�n��c|~A|r�k�.�+~dþ�|vW��s�Q¿�6�.�~]8���w���b�w���� &	�g� �/�� |� ~@ ?t�O<ax��}��V5���J;*)�`�J_����)�}J1����A��x�T��.���O8<i�;@�ͪ�Ɨ��c�[�H���J��Ro,K�8�z����驳�ψ���/l^l���u���9e��y)��ں�[W�zk���Y������کt�j��G���g����3��%���V�C{4�d�?�ڲҀ+��a�[� xEml�p�v��j'��pY-�܂
�U��[�2BT-�fՉQՅ�Z�����Z��ǝ�{y��b����
>�g"Xa5��p�o��iM.��l�8���5�>�P�X�����������p��.���q�s@���w�j/_�S�l�fCU���Cx�ܵmQ�ͪl����~7֭l�-!s�U��I��+�A��:.�k�w��E5t�b����>[TT�Lp[԰�@q�Q�5� �� �ⲙ9Ǩ!��N'�.5�^�R����l��z���n�?eK���J[��fi���jLҪ7n(��c��u��K�$���v���Y\T7K�he�Ŝ^!�.%�Mf���R��AЌa�Z�W7ʙ�J��N�)�TM�C�i�k8�C�@c�H3��~;O߄��f؉����!}��g���2���Nf'�
X9��`m���48��ŋo~�mj��j����Y1��Q�v��4Ȇ+w�vt��PK
    +Q�H<l��  �  .  org/bridj/CRuntime$MethodCallInfoBuilder.class  �      �      �P]KA=7_�lcM5~�Z��X��/~<i
��B�dG�0�	�ݢ��}
(��Q❍��V���{��9g�=7��� 6�F���4�D*����Ī/�}��B�Csb��Cy B�'~�@s|��d7��%L= ?�1a�oN��?�	�eT�G����%����%!��!a���"�	y1��V�5��j�1h���<L���J˶��61��yWbe��ׄŧ�f�๗���|T0ϋ��.��4�]h�P��-��XDJt���a���l'����;��Tv��l��+�&�ҡ12jh1�!֑a�ݗ9�9V�/�L��#�~��e��qSx������7��(�-�E�+�x����#,�|$��	\��%O��c���3|�m��c��Ӗ��(�PK
    +Q�H�ۃ�A"  �M    org/bridj/CRuntime.class  �M      A"      �{	xT������̝��@H0,2,JVĀa�$ 	 ��ę	�u[�j+���*.qPBAk[P���֥V[��v�m�~mm��;�޹3�� ������yȜ{����v�/���D4U���$_;�-��R��+�w1�q���m�d<L.��{OSQ��������\X���X�>�4F�c�����T�w�it(���;�K#��~d�g�T�t���L�'�Ab��F�L��-���)]�pdJS�sbC4߬Q)X���Q�S�2�Ӡ���F��d�HL��0�i�@�4ɤ�\ɐG �R�n4�3�ؒ��c�`e��h,�R��O�
���H8�v�Bsh�'�l�h�E4�ui��Mdr���F�7/���I�ZaD�@Bn��4$g]�
p9��ip�XN`�I�'0�4��#9��"{f��BS�F{�&�ȳ��b���P��@p���ƎΈ�aȫ�j2 c�`W<��)�d�#�2_��0ځL4h X���?{i�Z���qH�htE�������Ő72�_�b���k�WP���gcI�-�8��>u`rpr�7�B��X2�S}$�HHF���j�µt����XN�"F؞%����s�
�+V��2�/4:�F0�4B�t�Ms��S��>75��t�NS�D	Z��ϟH��-����[�Ӳ}�E�FK������� �\�����8}��x<���Aj �J
;*?;�L�˳2�Sn���/-���<c�>�ڊ�fU���i��bZ��L��4�fr$ׅ!��Ks}�1z��P��&�W�Bf �[�+r���\:O��|�	� M#����|�FA��,�w�DSd����p�A�^
�Z��������a/��z��`��37�GC-��I幄��Y:E�C�#�I:!�c�#����7�i,�<`-��Ec4�@�a,قJx�YO6[�԰������ȋh�d$b�0��Lv"��-�s39l��Y�֊�˳�R����^�i��R���
/]FW"�w��5"�٭���C�koÁ��H� �cb]�+Z�Gۛc��F$�h�³v����)��#�r��WM)�'�!*}��K^��t��B�i^�6�qMg7VLzA0�<M?8�+U��#og2_�#�ynb$Q\�:�c��I����N�w�Qs��Ws���p[<ߜ���=3�m^�د1y��)�t�6]�7��:Z����`wY�!��v��������|K�K�{[��cIG�QO�Bæ��iƝ��?�vo�����s�QzL���*�HY�NO�}^j��l�vAށPH��M�w{I�1Y�h��b	�Yl��4��a'�����<5d��?,�%�~7�q��ӈ"?�)��R*r�R���y�����%3����sX�u�6}G�����ZƆ�%/I?�̹,��w�ɲW�G ��X(�6�	��u�>�&y�dX�R�~H�z�l��uzC*史�n+WHeH���:��[��\��M�㥷��2��pF��F��2�zh#>%�Q���ⱎ�������$�@.�ؒ�p4��G����,{T����F\'���_���O���k�k@	˧d,�E��њ����
�7����u��E^H4��:�����)�r��������_�����f��&�����P�*�|fN�����h�	�L|�js�3`z21����{i2f��9��uF6�,�Cb�#s�<�u;�i�
rU�Ѱ�n/�أ��t��S������s���F�q1\ă�U�଒Xe�2��x��K�ޕ���F0��+d�a0nLy��y��\�\�a���x��}���ᄉ�ΣL�Gg��^�ܸ ���c����X2 �9e�=�؟ky�e3�aTť��=�<n$�����\*��F��L�u^����D>���hNv}�qy!W�n�|8��љ�.UA繂�����|�3�#:&��'"�I�if����:OG�'��L'䋚y+�'�3�RVbB55��ϡ��۱d����5��gI�����nF�<8[lD5�f��yb�x>��.�����!N���y��L�q�Q;�x\���<�.c��Q�ޝƍR�K�ܒEr:ia˾E(r�g2�OI����͟�V�x�������u�y7�d��37�����+޲|P1/��$9;*!��H��KUG�pށx�F�'bSĈbS�	�N-|�/\D4�2�ŀ��R��Z�����ؔ-[��(�C��_u�n�E�d{Q4��q��_3�(ǋ��^ �=i��u��9W�I�Lr32�B�l_�����9���S�Q.�o����04; ��zo�q�"���-]�F<h/�����|����T�,�i���\��^��±)��2<ȕ*5[���\ "��%.)��}��טݓ��:8ؤ���t��Z�>������P~�Kqb<gs,�H�*<����l�r�gD�d�,n��oBq�_�W�?�A��f2*��g�J���:ْD�؊D)��q��	�BF[��6U"2J�2@���f��4e����:$�K��5f�u*CU��F��{���{�i��Z/�>wrs�w��}|��W��j�"�6
u:��f?(@Η�����x��ih��%U.��QF=>��z3�M��OB4	_����ո���I�N�����U�<�ӯvt�MI����(������h��	���gp]�, �A�P~4 �gy�D� �#��j����)�o����7Z�$���vk3&�cv��P�C�d��/"���SB��?q��_N��J�Ƣk5~E:��iƦT����
������*������?D��]k^*��N:F��^t��񸟦#~`��K��r�Tc�w�ڞS��7���u�c���=���xc�?g��f�Q��e.�ew�?��?�5�Ҵ�e��S�q�f��B���O�H̖ C�7�_�����L:���6v ��g�C2{�V��(��F�F�PUq�7^f��|E��Z6C�:4����]�!�%7�+M�PAU~˿��o����Of�_+��?Bx��x�h��`^�5��'���?�0�l�nD�!�F�r�#U�wZ8�|�G:������o:M��<pS���L<ز�]����A5�ԸlVŒ��d�y��+�9�o�N]������BF�5&g�B���f��pzp��վ�٨	�����օ.WxD�ο��9!�pk�|�
"��☽�e�\�qF�ܕ���]v�JU�5G���$�C2�0)�sa�u �&�KbF�i͢ 9�u��EXz�T��\1��T'#����+�Sotdy���b�l�xl���&�}$��8�?�/�nI��r����@y�8u����������p4\�8��͑�?�Z�����S_�
�,�D��+�dW<*�t1Y+V��7�GRi��)*�T��i��s������ԁ'�S^��cYN�k�;�vHqy*>�T��rr��^��k�6�����Ꮀjw�y��(���Qr�F]��J" �
Nu�ݼP�k�/sL[:��ta%�/��\f�W��4!ߑv"��r��+�	T�q��Mɔr�S������>+4h%����+�� )e���q�|�M�U���%���],���yLs�������NJZ0�9Gq�2�a~�ʶ'Y��X�ҏ7�oS��B�A]���Ȑ
S)oF�1�&I��@&��Ĥ#������^6&&c>�4l�p��Xg���6"��BF4,�@��j[Wҿ��-b�>|X�|�D#.�70�6O�t��r��6�˥|Hq W:�<>>���DY����e�~YԂ��ˤ��k�7��r��ï�+<���"�����ZhW�&���i0I� �U'������'�}�'�2!@4�)�c�<���9�@�-_�&'���g��7S\����:/�	�xZ$�:�M��qۅ��Y�|3(n0n �o�ɂ+-��G(����t�9�3n�w|��D����"�("��G�47j⎣�xKt�Ut{ŝb���r�u��%�.��w��"�ЂӹGU��^$�2�����jj���H�uq�x �ă2���"� t��[cv}��|�1�W�?���F]<"�R�xn�̋Ac�!K@�+i�G�����7Ӳ�&���/��t������t1�t���Ld�/�H��A�����2L��zG��CX�j���4_����<��-��5�z�)�[ZԎ�o�l��V��3s�b�ݙ�r�����\N��O��[�s���.��k<��*����y>r�:�9�o�g#ַx����H��&�삜~h&�g%��#�$J����k������6�7����v�"?��)f�>
[�Q�EVA)�=��=^��]m0!sƛ�(>�귮
'�Y���,��A�cvk� ����[&�x<每fWY��9G��?�(U���$[2k���x�a�_�g���ӓyO��}��t��J%�qp����d���ࣼ��t�B1�F��W G����C�H��$�����+�L�%uGt�s˱���O��1�N�WޖXW<h�~<���h��|wB�H���\4B~&F,~�'A��X~�l?O��4:	cM��1������33ΝR<B��'��ES��	��H�3Qu��W����C�����k���qMA��-k%M-}Բ�V�3wJ��=��ͳ�������(���w1�����OI���E~Y~8�$_����R�45���S�ҪCT������:ൡI.qu/ź�]���e��a���Q4�:�B��&bT��1�
��@2��]A��'Zi������\��r�ĊD�x��"�h��9�<�E������D���ϓ�hr��6��]�r�J<I.8���*�����rt5]��;��%���H�mɺb�)|�!X|�D��������8���}�]SY��nL�~��bc꥛�_6����#<}��j��(�Ui�+������[�6u������ ��ik֍�֍?�ӝ�m�?Ϣ�]Y��Kw��G�۾םA��T�xi,5��6�U��2*����v���{�A��PM�P�M��W!=���?H�b���N�y-N�I��;�WAcK �EyG����'*{i�6���S�w��5u���s�^���������C�u.��\����}����4�g�i�>zO�K��o�!����}���>G/����u��C�W��7{�Q]��!g����^S��C���b��I���}���n� �<�j/�B�M�>��~����T��y��_�Ur��L���:�ϻ��!ǣ|9���z�{�������;˜}����^֫����^.^��K���R�u��p	�@maA�^��n��>o�>���W��#k���1�4�����
��>����|_�^��ȶ���_����Z᧰�Y�$��+��}��]=���
}�}<UqI�����Cn��˵@C�������>��Ч���9=4�NW��$RʧB��^^��R^(� g1�������=�7��	u�}ܴ�>�,K�>�^�\��>����%���������}�6�b�ߐHC�B�~n'<�Al������%���v-=�w���.=�Q1X��#����R�&N���Rq�zV�'�x)�n���E>^ɫa�ߤi|&���sh,�$ĵT�g�9T�~Z���y���Q����B.G%~&F:?J5|0�O����8�l3+���n���|#J[	��/�;�m^1��U/}���u�n��h^���~1���-�憈��bi�)����50�`%�(�1��xAy��*��N�-|!���6q�9I��s1c�gU
;��m��[�ѽ�h�#�W�	�"^O.�/E#�;c���5|!M��S���y#�Λ���6��˩���k�j���������,�����:��o��G�g~�>ㇹ��b��vr-��9�7���ʻ�<̅�p�Y���s7�޼�����m~�B�����!~�_��%��+b0_��b(O�̯��������).�ĥ��s�`n?������Z>�����)�˛�>�ZWA�V�������L�V�����t�6��z�<q�J}�R��*�/P;v���@� �\����&BK��LKh��R��h��2�i�#KsJG�9�#Y:B��:bGL�н�UZ�L߅Lߣ	�>U�w*@3�C�^Q�T�NoX��� �;���ҡ���	�M2tg�)7�ӟ�_`� 櫬��K��j�b��4�/�-�/V�������'9
�)�y�P���(3��-���,� !ò�C}.����i>�9v���:��O�buq)�*��t�}|�j9��Y�~��xU���ne���u.L�p�����9!��!D,�?(=�!�X��C�2�?�q��D��}O���Оm4L>� � ������[^P�̳A}�&�E�K*�|�zz���&^O��JRE0��,�v"Y)�
�`ݴn���.���o)�y��Mf��C�j$�Q�Fҭ:�H:S�I5uA%u��;���M��Fb�o��w��� �4��E��o���4W��D�..�n�Lx�j1�n@0���~1��#�}�_���(zIG������s��`k�-������D���I��4�!�#G�{�]s��ɘ\����=�;��2@��G��09.���}l5nH�V�1,^��'����/v�/-�'�O�RQNǉJ�j��O@Я�5˴�le��Jf���V�I���z��F���ۿ[�}�ş=�{��ZCE�yn1�TDb9͢�E��OU�J�F��4Ĭ�'OF�XK�bMu��_���u��I2��~��O4U�!�O�W��,���u�T��A�<>�q�LǱ��D�P�H�d�r�o��I�D���qF��`�q*�4V���eZ�,_�UV9�;��;L���~�<����sj��Q)@<�
F��c�Qd�Cd�ې鋱k��s���\#�΁ZgA���U��N�>G�k��{2=v���1����r�Ok�9��+�g讘(݇&��8�j�a^O+��]wu�.�N�e*	s�LZ%&�h<q��9 �ޜ0��*��$]6'n�La$]�|���t�(�YS~�`$Πb�-�_+�+�T��#�Y"΢fq6��s�&��*���KT����+K��^Q�\�?uO�sV˿(�|�>qR7� +�&g�c*���N�kT�O��Am���mr����b�4�v�2�9]����nw&�	03����^%f�8�F3�N:C���� >�t1#<u��(Nz�`�R�R��ü����o��o����~p@T(�i�XKbU��t��@D����p=x�	�K1�y��T(�=.�&� �9��P��%�� �X�+Z@��8I�T��>�h�D́ZGA���Y��N�kʜ��\��$]0g���dt����8�4�%�ƫԩ ��tˁa��-�*>R\�*NS\v��F�fm�jBK���an���{M_ K��Vdx�"c�U�Z��I�	&>W�XZ*�zŊnҫ}.��T�S��UÕ�K��*��T��TU�Tͳ��gY��@$�*sf��|0����
Pu%(�
�W�\q�6~
[�1��]VϮY��K�4�2Y�W���j���vE�YndU�93�1������[T¹T�Q-����,:�����7�q#|�M��U��_��a���q'�(��/�����\Y�G�kf�.�c��<_���!�M���y�Gi|΂�"$Tw���pP�3��je��DV�O������QU��ұ��c�ȡ�L�O��d��q���j��iZ���j� E3��)A9Ӡʴn����Rqa��Ṝ���M�J_��P�TX�׺}�u��ï�<i�mG"���D���_I�-�v|G���<��Q���3���N4�g���6�}^ds)(���_.���E��Y�σ5��)�SPĝɎ�1}Z��q���t��'��R陂��҂�s���"�V�i4t�Vx����n�q��m4Z|�.xһir?sBlG�y=���D!�|��G�S�8�U<�B�`M�d����)�*��b7�������^K[[!�Z�q蔹�r���m���]��I/��	�6:�*�\�����URQ��bnZ�&�`�R���k�������r��x�]a������ԑ��Y�~��Z${t����;����HۦG�m�2���is&e�ꍂ�dq��!��Kw~KW�ka�&w��9��X���A�-��N?�����E�F!fT�	��P�� �5����`�� ��*n���,]�t���+��������3���n*�f�G��+zzd����GEk�{��}���8MW��o:�d�!�	������I�HUCmZ����T5�b�����Ř�a~��e���U�,��<ݴ�w��D>ӻG�m�����?_S�'^�є�@���x�vrղ��x6i�#�`�+Ə�����X�S@h�䵊����"qP�h5��dF��j��ڡ̷4���?`p��I��//�M�a��߃җ����ZՌ��y�J�n�tK��>���W}_���Jd�H��x��>��/p���i]�D��K�(đ7��^��6ˢ�c���Stw�x����n,hO�g'N��i!|�"��>�� �S�Dj�¢����P�!T�� �������^0�O������	 �#��ry�PK
    +Q�Hן�l�    ,  org/bridj/CallIO$GenericPointerHandler.class        �      ��]O�P������"o2ATD�)�.L2�nY���l;Βڒ���{x�˅^xE��(��x�2>g-����&OO��y~��9���� ��3��AݮNm�.p�-�������x�p��@c��ϸ�r�n�WvD5T�Cj7AEC���!c�P=�A]�[/w�x���c��rg�Aۍ���*wn���;��0L�ǁ��=fv�� u�bȀ]���������X�!��T�}<>�2��1�q�0d������`��o��_�'�w�Ș��t�6|DTq�N)����Z��A�sf)��$����c3*?$�R4���f4�ak����my�c+�4��#c&$ɖX��i��g9-�����9L�4ܫʋ�p��	������+�ؒ�a��x�a�i�)ڦS�x�h=�8ۼ�B��M�T�=GE�Ϊ��FC4�R�J�E��I�+��F�ӻ��� {����"w�o�r��r����gR�$��<pg��Jn�ֽd_�}C�[��P�#�w�C�MY_0y�K���Z�a�cl���{�nyߡ/ٸ�9R䮢�YF�Ĭ�Y�827��������jI�kI���?�|Z��c�R�Vʚ��k�=�ڜ�w��<�Z�*��-��^ PK
    +Q�H*�|H+  S  *  org/bridj/CallIO$NativeObjectHandler.class  S      +      �U[Sa~>AVpK<���%,(f�A�C�	�:����C��,��U��.��8S3iNM�������$f7/��~����~����u�2��z>����v$.
�5��l���Zf[�+��+(� ��ݖw�HA���)�Ah�}�ݖ=ů0�1�=-K�H��L�]����x��˜��a�_�<]�;�-$��D��Tb�M��P�!܌�B�z�F��<�{,�ͽ�a�ᮮ<)PP�{(N�٨
k�[/�����_�����[dJq�TM5����	k�%����D�0��E�E�ы>n]яn�28��*us"}����x�[���P�'��!kYB��`�fӴlZ\�e۱�l�r9]�s��V&"Ƀ B=y�h�gٻ�V��ILq�MV��e)*�x�ꬩ��	��+|�|�VO���-Nw�a�QF%'�"`���Ԋک��G�c��3�ڰ"C�=9�D��"�b�Cg�x1���P���:M�/�NW�uݒuU��M~P%�Aڅ��'�j�j�Y��i!�m39�5�~���i���(�����rYbR��ԣ�p�z��?8��O��e�)�o^�`����R��I���~H�����:��>�%i� c_	w`�NɊ�|W �7sq�OY:L��q I����SvV��/e�:�|E����R����*�Q<�N�n�}��GK�0r��/f�J-�XS%�_���Y\fޏt���
��s���Ǝpg��$Zx��~����۠����(Ws����,b阚��%��~�m�*㵹��C$��r�x\x�T�K�H���'��]�Wх3p�PK
    +Q�H�#��  H  %  org/bridj/CallIO$TypedPointerIO.class  H            �TkWU�7�2D��G��Dh��YmSP��A4�!���
3�ɤ��p-?��ɵ��B�����rߙi�{Ϝ{Ξ��9����o���@�v*��,�e�F���6��݁,�ۦ�JgeM���3��aU2k;{��j��t��=�}]����	�]:.曐٪Q��̜�-���_��/2��d[5ש�\ۡ��dG�VI2�m0~������,���.
&;No
\j:��J��5mK�E����f}��#���УaX����ˬKә����+,�Fq})��T櫸ʠ�t��"o&�:Y�Dxq$t�b<�^Q�^��LzP�\s_��yC`�y^pӪܩ�ղt4\ӑ� ;�l�UYN�v��HÕ�n�X@��@Ze����m\�`�r�
���F٫ƾTM��`�n(Ao
�]�I������vm?*�wTP�
��`���x�؇�NU��|_�n	���P���ϫ1~h���/�>jN-y��~V�����閤MՏ�j]��r�TH�|P�du��]���6\ò���A��l[�W�c��`���T�Ϧ��5U�����������(�YcaD���ǻق�˻ 9���Rr���g0̩�Q��\|�#^Batf+������s��ԣ9�h��X�[w؏p�.Kg����j6�B*�N���%W��;�	<�����K�$�g��
���䲩�c+�%S�0Na�q�zehC+������^\�݇~����;s���S'J��b$����b�/+c�)&c��sL�#Y<��@����1n��m.i�>�{3'���g�A=Vc �6������c��"><�gkx<E�页C{�mj3�-s��2�$�h*1��}OEa��x���Ǹ���.vşa��r#�d�U�*�3l��dV)�񥤐PC�8&<!�lن�,ְ���Ϊ��g��,��S<�h�У�Cџ���FB�B�x��6��F�"v���>o����n|�b��G:��R} �"O�4���'�p"��nh�q�!�x�-���Ϻ�PK
    +Q�H"BY"  �    org/bridj/CallIO$Utils$1.class  �      "      mRmoA~���/-�-��R�T��R�i���	�	�/~Z��Y�����&��� �q�8��|���gf��y�~���@�m��;���k\��E�2p����`�>��W�����:[cb�!9��t	Cn1���ٞ��hs9�35�3��IÚ�_-6g��)$�dX
	�#.�B����9��G9�s���)�b͂�,C���l&�C<�r�tgn�:{R�u�\قa��(6gu���	�w6q�f���K�k	����s�<�Bcn�w�i�)�&��R����]�'�Fc>֠�{"8��oh�ʄ�����̏�3�ː]�Y��v���6�m�9�#�[m֚������"$�r��-Ν0|�l�������eHՕ^���qL�= X&�����8}�z@��0�L��b����t3pH6E9�l�����yF�&v"����3�[����O����O�$��>�h��T:�;!����!�k԰>�b���#�ʧ�*�W����Q��~J���P����%̢�4��X�PK
    +Q�H��)6�  �    org/bridj/CallIO$Utils.class  �      �      �TmSW~nXv��!��J��,[��-D�b�h4!�-�[z�e����L�����_m;����wT��n�$����L�^�9�9�s^�ۿ_���]��/��=)�k�vݍ���P���0v`�b[���[[{�j�2����|z�kd�@����,j�.��w�ǥhn����k{�˥�a�ɾ&��F�ן��):##�3�33vp
�n���s����0��'�U���\��L�a�!�(��jI+D�)��8L�X����"�pu��I��?��SK�V�R�x����sL|�`�]1��u�j�&ذ�w�^���Rw�u�rӟ�D���.2�\�*��^�R�\^Y%��
U�O�(`�D��lŽ9�0D��@�����@&�q�@�3�H�y�򘘅e �/ToD��8�:4,1\$�;���ŷmir:O���O��/	���p]���ć�H����8�:�V��= n0��H�p��YkA �=5��/�k���-�S�u�k��TYJ�T0i`T�F��Z�'��!�JM7���!�s�U�D�Hq�x��nR��}�r���M�m�R(�u�!qU�������I!�FوzM�[���R����P�Hܴ��4Ć�sr+�M:�k���ߒM^������� �Qus�~��)Ul���������E+�u���?h��C���C�����k�t�=��%d�S��.|�@�yL' ��٧+P� 
`Fd �p��Z��rr�(��f��e���c,�o1��Z�����=#"Z��/���1�9���?Q:�D~����0|���K�ys�Q%�nG@�}� �S�X�e�3�GUzDLjA�D>�e50������n�y�����~G.�J�v,Q�A(�|O�
��F`:=��o�hh���9J�� PK
    +Q�H���  �    org/bridj/CallIO.class  �            mP�NA}%��"�8�\L1�ŉg�b���f�B�t��`�5~�e�c"C���^m_�� �qFh��4��$��=�u�$:SKje��p2��y(jk�U�$\n*;�l�&�h���A�X��P&�[S�N�Ɠrɒ�M�*T�-	�yN�����o�l�:��?Fh�T/.ѩ�}Bieʮ���&u�D,�����Mn�5ew�;���tOb#Φ�&cT���.�R��7r��Vi�i�A�+	�h�G�W��12���/�T�B��x��Uk�`O�!�<@�PK
    +Q�H�$l�  B    org/bridj/Callback.class  B      �      �R�NA����"����&J�
����e��u�,�$���4� ?�� (z�0]��]==�}{yp�]���5s�'�\�;�����R(��k�Z)_��*�\ˎ��Z���	�3��w�m�gX�,3dX�Cj ��-��KC�q�r_iy۽&��/���.�RI]dd��b��a�!��e�!����׈�h�ҕ�u2١�>M=�1�����K�����I3cX²�E�i��۠'�ʮ͝:�$�Q��}���e�Ĺk	��D�����=�W&=d`�Yu}����J�ͭ˶�1'J���wU;��)2���n��ܦ�J_'��0����#%�Q�}��E�p}�In�	���9����q�Xy�Ǹcl�v�"�g�v��C���F�PK
    +Q�H��;z}   �   !  org/bridj/CallbackInterface.class  �       }       ;�o�>CNF���t���̔,}�Ĝ����lϼ�Ԣ���TvFF��ĲD��ļt}�����vfFy�6�Ē̲T��VVF1�@�12p�%��e椲1201�002�1� #�db` PK
    +Q�H(�7�  q  +  org/bridj/CallbackNativeImplementer$1.class  q      �      �T]OA=�+u�� �,��ʂ(�c���� ���ۡ��6�mc���F���$>��Q�;�
4P���ܽ��3��3�?���U�� ,;�P����"w�o�H�ņ_�/T$Bk� c�OA��T$}am�h?(�����I�$B�S�x�3�tq��$�`YD�����d�hN�yYy�X;�J9�@ՉL�ڎ�X+������=O���Ө��w��[��k�Քy�F�i�
��鋏6p�a���5��HM���4��'�{�K^��'�ӗM�!�˪�Dw�Ѕ$:�T2z����*��wM�V?z0f�&��u���֑L���CB�0�͡�2��+���b�#ms�m�ϖ&�48y鉭 �5UZ���JS0��=����	�Nd�f��(wV����d���<�4{?�f��M�w��\�Z"��=+tkvy(y�;za(H%�j~Q�-O�i ��BW�v]�^P��6[��J�0��jUT1MZ&��I��� �$���7�Q0<$k��{i�,b<�=�D�w���G���0ޥ�1}���V�P�f�E��,an3�����x��v�3݌�x���8�Ha�Ş��z��L�/d��Kj��+1W��>��5N��/���Go`�� PK
    +Q�H���&  �&  )  org/bridj/CallbackNativeImplementer.class  �&      &      �YxT�~�d��9�$�� ��Nn��P�D���� ����$Lf���VDAD��U[[�z��-�2���vUZ��nw׽uo��nw�����n��?g2��LB��>�&�3����w�������/�u@�\�4�F�}�Z�P����4��]f��P�4�q3�*�����hh�XG��SK���&xǃ!{}��+���)Y/T\f���F'\�5Aj�����..#��]��&�=�A�E(�	�y����uf|[�O��C�����lj'�藜���T�����}�{�p`8�FJ��p�۶�jDfH�ܑ�#͵�nlS��7f��j�sVP�T�4ͮ����ښF����*l��j�*�椉뜴Fjg������lϑ�HC�`n�4 "��o$l�vQ~i��l׽>y�9��z#m�Һ#�5�#Mg����4��X<}S�f��6�)��4n�l{����#�P	��asO|�d{���.(l����F������ꍓ0�>d��#�A'�������L��KM�P��J� �)��7z0u�\13<;� ����6jX��\�J7�p�i�DFpa�b�Z�ZP6! �˯�I1�U��Zt�Q��<���J�#�-H$-�8Y��S:�l/����s1O	��N��~���P$w���y[87�F��I�3���thh�:A�oZ�ڢ���7*����q�
΂k���i����]Y11�zO����"�∙t�7�ngMb���`#6)�������mLC�2��$H'���q��la��\u���̡��vd���5'�^4`�^���* ����k�a����YesO�O!AlW,v\����R~ aA1��Ri�T�z0d�����*�.�I�ƈ��XjC�╡��G�9R�MNu��KC9v��TTN�04)r��N� ����=Y�<��p'�T�'W'�Q�1�bv�W�>ܧ��m���
��G���s���m�-#q�֖;򛚩�i��Ԙ	R��F�>Ơ�"����*��d����h
�9���W�Ƙ�W爛F��񄊤'���9�Z��ۖ\ζ
�L���m��[��'��f5��|--1|���1�!��*�
DM#nVǓ��������i�*�DwU��V��,�J����2���ف����5�döhd��2�(���g�9p\�d.J�jK6_-��5A՝�2Bt�԰'�PF�Uf�����d��3N��&oI�Ak�V����
)R/�he4j0��zZ��B�.�.�֬,�by&��ʴ�$�2͋��Yl7l�کbB"`�%��:<%t�6kB]�5;s7d�V�=���
�*�K�2���F-G�L�\f�^�T�go0'��f�x}|����T�o�M�٘���3��6��u��t��G�T�
��<x��w���:;!���wUa�)N��|=ShJ �����~�?P�����TךF�	)�(�(��?R���V�h��ӌ�;u��g~�?'�&8���"��jF�ζN�5z����a��@���c�d�|?跿g�oI�S��\��G��bג����-���mH۠M���w�����W��˖��k]R����J�2cA݌lH	�/�B����j��	cCą_��VN�Z�\�k�6ˋ����I���9�b.q��b�q��u��G�#����r�Mj�3��)��h�KJ� �2��I�fD�̝�&;����s��R��S.����s��c�Nfip˅������"WorNM��2�M�\$�5��a�ϭ��/s5�/��y�
O0&�RV�!*�eK���9��/���\�z�P���d�Uc�Ea*�2Y�(9�S&i���0I�������
�x�v�QU5j*���>+T���ɀ�U=��;����7W53w8��o�\�'� ���eʝ�H�9�l`d�5�q¶ϵ��cʅV�����+Of��C����͏rQ���a�=������k���f�P4N�D�P$���kPs�d�6{�ؠ�MѠ�Q�6M�U'Q�+r#;}mm�w���Y<�C�Q�t2S["���:�+7��r��p��]h�3�����혙m��V-�(����7����Ƥf��c:��t(=r;[����0z͐S�jr����,^֤`�o�FY���{%��ӹ�6'��;�{URj��ϕ_�(~LP��F#��1�l�`��P�q��{l���b��b<4�_��#Q�Ϝ����|��]|4�Dݸ�Ө���)x�|o$��Q�Dly�N�K���q��{b�k���s���p�G�u�B�}��x�e���k�_���q鐥�|9����s�F�Ԩ�n��LKbM��,��5��_���zLP��B���u�#W��t�u�a�}FܠO���ſ;�w��U�פg���҉�I�̚L�d�\�޼���ǣ���>]��η�6y�Rg�X�;�7^��֕v?�i��h��A��,'�~5����a?/�l~z�O ��"\��
u7ϧC�H�����Dϱ���cW>�o��`a�IԎ�1�EݣXrKk�?r�p���'����V�ԝ@�q�S>��*�m�b`��6b��>y���,����:�S���.�Ç��G�[�U[�v�b`v�KX{�T���&��N`��:����lٖ�K��Y�
�����Ej�ͻ�^,��d��6��W��Y?�x�w��!��� �ݦ;��[9�@����@�_�\�+щ��xr��-\��w����]c�׭;G���V3���N�Q�^�;�]ӋF��C��ޅ�{N��|��4�O�)��/֋�D�^|L	���>uJ�g��j���(s�R��Cw$p���Q|���c���m܂W��̷\�4J	���t��8���|��B����L׆�_!���������^:��4�ϭ<�Q��R|��6�䦿����`��j#R����*�hߦ��/s._��l�m�_�T��	r���$I��
73T�[9�M{{h�f�t;G[i�A^��=@���o?5�eAr�N.;�0�����P�!�1;��3ԅ��$T/�_ԟ���Y3��׾�ob�Ph�3����M�����$85�3ݺ��Q��/��O�y�D<8N��S�~Ï���Q���P�k�B5vr����Sx/�z��w�3�M��oG��;�"��/ҋN/��/+�,��A�^TY��_�������I�;1�����@��ջ�����>���W��"��/tR�R�))�B\
o��7Q�hu�x*����o��'�R/�=*"
����Q_l���9N�L���/�r����[Yv���J~��.�^]���'cpw�ԍ�l�w�w�%���	�X���%~��,�uJ.��&9z��^+v�0&�	Y�@r����V���NƏ[ŏ�:�M�I��A������@�T3��Tj���c��I=!�����bR\"ye!��"�ʰY��FY�2y�_����V}�g���wY�T,�a%rn���R颴e�r>��r�\C~��x��)�3��5I3L���F��h9uv��W�:Yɰ_$J��"\��nY͑2(��Z����
�&rUJ��2��<V�x��x0�[���u	�����
vk�>,½���D��&����\y ��S�A<��臇�}μ����G�OP�������O��K/�n��8ʽ���yy_ l�D��A; 勴K�6�I{w����/����K�y	�Q/��K/tTȆ
����n+�˖1��{T �Sw��3�;�:#cPw�a��~/!;���	����z����*d8��*ʬ�k��.�Mvw�N�#!����za��*i�p2!�ǡ�
9D-�>��C��QyX>�C�<�ɬ �J/��;V�k�JB�5R�̷FǬ2�Fǭ2��u9,��0-�~��Ǹ�/���Z��%�������u^c����L�oP�7q'����=z�e�mR����C|?�.��(cN�ݵ����jj���N'��	��~DKY��SIK4��'/-9�+�Y}������<��I4&��\�n����~<#��"�Vk���C�n�E�M%+t֞r�!�_PK
    +Q�H|O�+  �
  "  org/bridj/CommonPointerIOs$1.class  �
      +      ��mWE�����	%P���X5�@}n"(؍iS%�n�&,'���&��<ǯ�'�-}�z|�ѷ~(�w��&d7Zx�3w����sg��� ��`X6�V�n���m���4�����,�b�^����A��X,��j����BS-�*l�|b%�G��p���|	�TQ7���jziiͶ���gϴ�2���Vm����#�$���#�f�U��T�{����8
__g`
�e��R�Y^�Y�����aȤ��,�2>����Ee��l���p�)z�Si6m.L�2��e܌�5ܢ�Y	I�Tmw�J�a!���e��F+�M��$������%änjϩ|%*G�qַ>��C��k�9�N�DWq���S)�R�H�(3��L�W�]�s�����Tݭn������E���;��-���<�.����2�1�qC�7R?�h;�ښ��Qڤ�iY�ٸ�t���1u+�E#������m[��M���h{��I	��eP�c
��ĩ����.����T~�ˑ��;�Ÿ���-c7��*݆m�P��fCm�TKW�m��?��/O��Ѳnh��'u�3�=�e���E�W��W�������[�<mw_J��U�R&��u���]���������i�F��92d�04����l�ё:/���[5��o���W_B~A�	��g֙���}Q�h��:����)�k�bmq����S|��z��9�)��3�d�z���7�]h��Ң��[H��g�!K�!_{�F�$��q �D�/�!y�1�����{����\j̥�����7�ǆ��ƀEe���w��!>�C8����C�|v�a�'�U|�$��t�
0?_qpF���{��ܐ��p��==�{Ip	������s�D�O<�����b:�g^���1�\G)�Q�u�BO.9J9�^��%$�2V�M���&�Į���p'g[+=|��7�!�>d�|ǇL�����Ϲ��>'��aG�+�=|u�;.��+.	���'�c��T�M���}��v�`�PK
    +Q�H)���  �  #  org/bridj/CommonPointerIOs$10.class  �      �      �T]s�F=+ˑ�*�8q�>m�N(�ǁ4��� &L�&'�QƑIa����[^I�L;��[g�Qge�6��ԞY]߽{ιg����X����,6\kw���8�Sǲ}ӭlzW��4�\�W��]�K֭�^Z-	LETjP��o�o����5h#+�m�����<Qlv��{-s�/�{m�*}�-��J�mI�R��+�eyk_�╷K�����eQ��M����+ҁ�!5���d#|,U�C>
��4̲��ʯ:�0�D��4�����Ul�����$����+:.b>��q��9v�󒪎+�*K�u����r������.N���v▽k���U^��ǂ5i�v~[ ��m�uh�lNvw�J��ؿ7��L�Z�G ��wd��$[��H/�$Wh�7h�ш��'��7�����G7����>�.��%,��`C`r��4��å:Ҙ�H�_u��5%��c���2-�.���IN~�1V�l���A�t�Lr�jچ�2��#j,"��G�Bj�9tẇV�r��i9�e7��+gW@�ض�����N��
�#W�I@��T~��B���{�'�c�q]��1�3���0�S2��$�d4�i�?f��{S8���#2��r��^������8d�Q�B����-��6.#D��#�n@N�+'��7e��A�_�"#�O��*0�r�@GB��&+x��Y(��4>ˡ�xGֹB:�Q��;F"C]�����1f��'�|����=�nN����]��P��~�:'p;��^�X�4��1�� ��U��6�������Y+����|F��6�u=��*���Q��V;�t��O��C2��sȰΌF�6����l��.���B���PC�1<�#��S�!�@0�Jg�>PK
    +Q�Hi���  �  #  org/bridj/CommonPointerIOs$11.class  �            �SmO�P~�(��*0^7A��a��Dq�n�b��o�VFIiI;� �_�#�����e<����:�ܞ�{��<�9��~� �W3�YOWL�v�������P��b���LFc��Z5�n�-�/z=��e��!0�w�/�'2C�7��a ��jc�a)^�'Қ��Ӧ��)�Fz�㑒-�m�5ٲ���� B!��
���W-���?;%����^4|?��
<Xe��%�#]j��J�a���l1��#�PGJ���S��)!�p\'�.43�Df��hl��Y�Y�E	���p7�����a�1�G�B����醡_�k�)�T��m�o�]��2CP��,k�
�s�KX�
�Ԗ���d�xɾ����U��]�s����؜�W֚�v��o_���#�pwA�&ݥ&0ɑr4��QS8�Q���l�rESv��0q9I��*��������n&���u�qlR���o|��.���}��1�ͪ���*7��fX�^�4���T�uŴ���
9���+}�`X���`0��^��tNq�Қt�k��Aa�N�ha���(Ʃ�Œ�7�1�lP<�3�ZiT���6n�"�S�/���6q��gs��T�1�����F�t����"E-��S@���%ryO�o�y��?!?c0"4��Ľw��G=���u�yt���$ڦ��7�	̻j^o����뻮)��E��4��ܮk�K�D�;�9��K��յ�LȺ��\Ebh�ə�+z�.���\�}��آ�@c^ڍ2[�PK
    +Q�H[��a0  l
  "  org/bridj/CommonPointerIOs$2.class  l
      0      ���vU���褡�GC��`��aJ�6�FIL,HK5H�Xu �,2�5Y�����x���./\z�C��g�t ̤��̞s�ٿ��{��?���'�{h2�f;�0���ܖq|l�OM�f�j�^���*w�P9RN�\G�۹����y�)G	A����w�j���%H���k�����T[����N������VG��|�.#�h���jí���I�/V�.���{�čU��Qj!�p�#�a��vY̗ӣY��	S,���������V�⡃�r�,c�F�n1\=TB�A:Q:=�ڢ"��XI��n��s�ư��_v��1�k����rV��B�|s01]g�tȪsŴ6�w���\_�`�&�F�L[򆖩�WyN>$5'N��(�`���^�ŷ��X	�5#�xҲQg`�&n�q�.�g�\��6N��%������a�Y4M�!�V%��j���ńk�"�"�}J\��E���	��k�/K�� �2�*�_������m����j�8��^��,>�"��.����e��_T�C�e�<��T:u�ԔFG�����A:�bb�����qC5�HdWk�J�g���G�O�{O��%���~����i��K,�k���_�ݯ�.�ڿ_��F�l�;���m��1,Mo?V����\�uմ_�������ӏ��`���@��h4��_~�%�cأk����u���*n]�u�ǭ)̐��d�bn
�4��!>t��!�{F*x܉lbsZ���MН&]�� e�@�$�P|n��jߓ�>=Q��NH������X�����Vc.5�Rc�ʭ��1���!>?`L�����|�BCSh�d3�_�(���#.<��#x(�lPƇ���s���>�g����a���Q�p}�p�.7��=����#=�+HpNƃ��o��&������}T�~Ǖy�'�eH�������(�*��S�Rĵ����u�Y�P�S�H-�#��&��G�B_���:dW�L��萩�2�9�1��D�Ů l�s%��o���N�Knp�.���G'(��g��B��}�v�1[�?PK
    +Q�Hh�g21  �
  "  org/bridj/CommonPointerIOs$3.class  �
      1      ���R�F��َ(&|(M�Mٔ�$��.-���!qZ��	��ld#�HI0�:�W����8�^t��>T�g�EV,9�i�{�������Ͽ�	�����5,��(�i��cS7�*U��$0e�g�/v��S5�Q�v�zhZN~=�0a)!�0��6wg�L� 1�tCw�V� ��Z���jgϵ|)���Qm;���H ���0ĜC�f��󦍒�����(|�+��]��~j!�0�0���[i̗3�4����`!	�)���n8�V���cJ9S���w�x����JXd�N�ΉVi�z�&�H�$�p�L�{@��a�j�?��8�^P�ʔW���P�L�!i�a��&o�oq�������R�}�����wyfS/�D�Ȑ��OZ-��h�%�6C7s�%��\ě��W��C��$}�5.����3G���hF�9d�S��R�2o��n��8�^�x!���U�x����"gnRt���c��U%|M;L�U�{�_B�s���6?�����&�X�I�Au�غ�\�N5:���C�M�SW-]mt�P�^���-�wtC{tr��,1���mCuN,�E�:G�!Y��cP,�Bm�~ِ�L�H
���j�K�G�M�j�XMm[w�e4;��퇚sh0�%��,���l�R�k0N�t���N�b�K��兕W�_�x���z��[�o)��	\�x|4�i���ƲX���<��(�aEzR�=��
wlyq
�z�����}�"�iч��&7�2$i(��k�h�Cm�)��G_��i�o=�!�b]�v��n�VS>5�SS��G�c���S>?#tc�=���'�Thh
������]���	���	|.�	�Sƃ�Dh�ާ�/� ��rp��������7�s�!n<ĭ	��E7���"6�������bjyq.���_;���J�ϼ£�2�}Ei_Q�W�F�_S�(�Z�� Ξb�=���~LmPKl���	ur֓��ŷ/]����!S�{:d�|O�L}�u��3�
8W�����u������<:1!?��Q�􎹇���s�Pa�PK
    +Q�H��/�)  _
  "  org/bridj/CommonPointerIOs$4.class  _
      )      ��[wU��'!�)I�KC�-Ŷ���VmK�B�(HK5HT�d �L�̐ո�ѵ�
~_��򡫾��\��a&5��l��g���r��߿^ ��aɴ�ن���g7̃�xlꆣYŊ}�ư\���k�}�P�vT��-9Zn=�0��(!�0?�&?�p�t��!����ΰ���,��њN�z�D�G66:�m�R5aD"�B�!���6�����$�OWO���[�ȍ�s�Ե4/�y��ɶ�0�P�U̕R�U�7	���{�J�e���*ȸ�7"�c�!v2���ҡ��j��F)xh2��$��ɀ�pݫԿ�>1L�Ʈ��JU���B�}S���1�dոb:���2x��[������(%ohY��Pæ�f���v[-���+�(
f�fv�I��E#C5q�T�w]H������c��_	v4���1�(f޲�#��k���W�4�$eFH��*�
�֩p�#��Sp��{C�^L�6	b{ �J�~J�?�'[����~J=P�^���L�rZ|�������t	6�]��6�j��Z���hU�`X8�H�XlL�uC{�=hh�X	o�mCu��w}t�̿�ݽwƣ~��_+�����S��sgv�������ȶٵ�ږޯ��옶n�jΞ�� C��߉��U���O����U��/��3K+�!?#{_�3=X�9�Ĺi��)n���ǭY̓�lY��b�Vv��֠'��s^�T��L"����x��E&�M[.2�k���2
1��dA�${_�'r��'��x���=��O3�2c.3&��zw�oH����� ��9��P�5�����P�$���p�xv�aFN��X�j��Þ�M�ӧ�.�����
���޾�\n��y���~C���Gp	'み��;�2�x�%�诇������s��ېt%]EIWQ�脢�"��!���g\e�u���i ���
urz �J�����:dW�LS?�!��t�4�\�Ȍa�	¦�Sz�>v��[r�KnpI�6!���A|O�@��П;֗C��PK
    +Q�H	�zZ�  N  "  org/bridj/CommonPointerIOs$5.class  N      �      �V�SU��lخ@�*�5��MQ륡��&RRK
��I6a1�fv7H^�錣��RG�}�>Gg���G9�Nr�Is��������}�ہ��� �0f,���F� ��-�e��n'���u	�a~���m.�hGZ����Xb_��-�o�ƺxK�1L��_��{+� 1,���bX���z����X�Z���V5%�q��-��e\�E��o8W��
���_c�����X�o0���.Exb����u�2�
wM%�h�oIs�}(a�A�N�Y�����L�*���AL�E"� ���0qs�e7](8\�/�
'�U��B5�@«ґV���e%��.T�kx]�,�Ƚ��e�tFzF�tI����ǔ�寮{�k���s��� ����R�ݰӞ�K�E؉��-\�yz�$5�&z�l�R�R)xB]�&EMÊ5<��\��T�e�v�|��ۚkX��qN/sC��N��i�,�yæ�Ty�j��娆�jjζg�,�F�R���������:�:�j�s���ضn��*9Z�����)�h��M:d�4ݖq�r�����6P�͢���ؗm[�2������v�}Dt�Ӭ�@�|w�\�O<͛���Nh�}�		w��� �
�v{�;�{��ca�� �Ty��>�I��*b2��ݫ�]W0�K���c�����i�-�6x12��0��"]Cbcx�0���aV����Q45�b���EG���y%��s
זVnt����@'Ù�s�|g�5۹ ����iU윾fԋ�j�J�C#rWw��<]�I������;t��Q��/?���#0|JV>���Htf��S���=#�u��!qn#t�[���0A���V���ie���¾�'u�s�G���E�_0�ب!�+B'�J���!�hy�X �&ߋ���z����Fo4
��"N{@pN�jx��w�ۃx��6 h��.�#���@� >A`�`�}+Ddi��BD����w�|8��)V�lc�=v�c���2>������'�s���5��K̙�Qu�"O��w����=^����{���7����"��i���x��:���S���q1�WN�i�C�S�=EA<��s��-��V�'�0�~��)~���ej�u���N�4d����Ӻ_S���P��:�zC�B��u��:1L�`X�%C�'x��%\��%�:=>!���� �����~�X]�?PK
    +Q�Hj�z�9  �
  "  org/bridj/CommonPointerIOs$6.class  �
      9      ��oSUƟ�����X!�vC��U������*T��	��L���n����+���}!�qR�o�P���^6��R���{��=��sw���'��ìi��uK�;ȯ����q��G�ʛ��[�R�����z��۪�ʗڦ�V
c������p����$���n��
â ZZ��5�|���V(6�۪m��2�H�0�qg_�.W�uP�{��0u���``en�d�xFCbZ��p-���J6T�Ax?T��P���4�s}W��f����J%[�1�Rx�F��J�c���vG�l�z�&����q�\x@��a�g�>�|����=��U��V%����m�T���\5E+�����%�v���
�+�]�Q��+�*	:�ҍ��I��Z���玖Ye3t3�yR��iC�����R	|H�[X�(>U?v�Ә��f��}�e]�,��!�L-�6�4�|O��=C
9�R�V�ƙ������ܼ#�ݒ���b�)SJe���Q��dl����j���/�I2rx%�><�G�1�K<�F�a���xj����UKW�m��ߨ[O/��#U���v�%V�[z�P��E�r����q�
���kŵ��ح�7e9[[#	���G�չã�&�ev��V��Bo��i�F���{r�04�}`j6����c0A/z��a��:��K����ǐ�=�z_��1��D��ŭQ\�|���B�,��0N+��=�W�w�NSD��w�T�ù�qL�]��+^>�s�I�>tW�����%I� ��]#������.}�iH����i9�b���v�����i��Tn��[���|~G�~��Ih��v���BCChH��&�_wQ<�'}x҇'�'�B���,����;xW�y98��]��������7��"�_�7z	�7�����߸�-�ss��p�������|�1���!�+���2��6q�)E��"��7$�L��1���L��H���ׄ:y��5��G�\����!��{:d�|O�Ls�u����q�$"t��ܛp�O.��%�<xu�B� �r?����c�K\w玹r�1�PK
    +Q�H?c\�9  �
  "  org/bridj/CommonPointerIOs$7.class  �
      9      ��]SU��'6	����b��H��ZR��iSAŪ��	˄��n��_�O�-�I;^8�3��o��ѯ������6�(��g������ey���? XB�aƴ٪��d���i�1u��YŊ}�Ɛ)w�x���z�f�����v��-�,3��,�e�u~��g8:^��0����°����Voj�Vv����\�M䛪m/g�eđH���־n3\,��II{��"��i>����ܸ�0�K��� ��a�kh-E	�q��	Ʊ�'F�;$��ar�.^mU�u���*�LA�^L�.2${KH1HGj��U������	�����2.��V !�d�׍=�>E�D�p�fB����f�s�m���+����Uf)v0�J�R�t�%\��y�4��F�P�8Ex�]��Ç'�(�g�f�]I�&�ĸC]E�Rɷÿ�T���\yHT�[ڳMM�h��b�wղ���W���R=��%g#���d@�ջ�U�qh�����>��%�[��>a�̔R�=%E�8����Mz������ J�<^K ���Dަ	L�M[�ys�I�YS�۪��$u�_&��N�e��n���%F�z�P[m��\��Ўkp�g������@����i1����T����:��~�f۪i��u��4m�h��Z���\4�r^���Eʥ�f�я��`�&��(�������C����]��q��oI�ŭs!��8���lY̍b�F>%{���'t�b���w�Tp�C�1L�����x��i҃�U(��!dHRć�s���~�gdG�KOT�i�=�"��,v��N�Q�5�Q��ʭ7����>>o��f?���5�-4Ԅ��|j<�u��x܃�=x7<�����KO��=����wP������� 7��*�_����q��t�1n~����t�Gܤo��08�G�voҞ���(�)J��;�)J�q�`�����1���,�S��2�J%�!�~K���\Y�|��Y��!{:d�|W�L��ꐩι_�a���.�J"B�x��
�<��\������s�J����U��#��7PK
    +Q�H2u�4  �
  "  org/bridj/CommonPointerIOs$8.class  �
      4      ���rE���e�.%�-V0�"�#'�B$|	%
X�`q�#y\�Ljf��*^�'`�l�[�*6�`�
(Nk:#E3��������}����o�p
âa�sS�;ȭ���~��t[5���M	�!S�����r��:��έFGU��J�a�'VB�anT�`�8�/Ab4]�W�RCHSmuԦ���W�š���bY�tMF��e����p��_G%���Q��uV����B�'���d[��)o"�O"I�)a�a��DЪ]i�,�H�һ2.��X��E	��#��U+-��ԮVFW"��$�w�>����S���>�̕(}��L���kr�y�q������%nt�Rb���B�D'�2d�̳D��:rg|��Z���-�ꚑs"i��vl����P<U*ǻ!d�u���`�4h��`G���>C�4WMS9�B��bVԲ��^�F�)
�So�-N]%}����.�]	�ı�8�R}L	��;�\���~Eߥb(��i/KF�&PW	��˘���}��ƞʥ��ҩ)��4:j��Mxr��X8[�t�n����b&���u��4^y�K1�~�~z�1�b��v�Ӏ��ULW��:���B���"�F�l�[Z?�z�cX�޾����]����f�M�ZX��N����^�`�Ҩ� ��l&����CO���8�8���w�h��4����(�FcY��`�fvh�3�'����xΫ���&"Z�~��N\d��i�EFq/�e�x)�����4�~Ƈ4��G�D�/���80��Z7vF�s�1�L>z�P܀����ΰ_��]Zy�	M� �M������<���.<����Q�l�Þ��&�uzz+�k��!�am�;\��ܐ�y�!�w�����$�_�'���f��x�{l�_�����G(��!�:J�����$�����C��W�?b"�����p�ɹUj���U�N�8�.�p�a?n�Cv}��������!S�sC=N�y�'��NID�a��w�[r�%W\���& �O���w��w��?���ۡ��PK
    +Q�HD���  �  "  org/bridj/CommonPointerIOs$9.class  �            �TmO�P~��(�U`�n"�"�E�+l�8A�L1�2�ߺ���ђv#�w�_�#�����e<���X;�ܞ�{��<�9�����w �x�0��d�P�Ɍ~x�kotUk(Fvל_���N����JԏJ1��b�!0L�b/��2C�?��a0�jjc�a)��'�uY�%e��T��#%�����e�L�J��%������5J�}'+��X��*��`�a��5����0Ԕâ���\�e#�pOJ�4uQȾߖA(�0��M�5�"�Nm5v��L�,Ds����b7�	ˢ[Ag��n�}&���_ժ�	ٔ��-�g�.�X�!P׵ZI�7:咗��&�-���T4w������5��]�s܆��9歬3����ߺM	�	G!wA�&c�R	���Hi�BF�*P����l�r����0y1I��Ϋ��yXV;(�5Mn4�7<tx���ڥ�������iT��R��U꺩j�WJc_�2HYMS�PL��~�_�U�&Ee��≙�sHg�	��v�q�:7�a��)�"Dx<��?�X���0N�-�y�磕F@�m>��}C�]b�f>�-�<��S�y��T�0�����B�t�����"E>?�Q�C�~�%�yO�o�y��?!>c(,���½���G�����yt���$ҥ��7��o���<�"5m׋�)��?na�̪��K�Dη�%r��/��T��31L"e3l�s���ǧx�\�p���`� @��=3��j�Yrh� PK
    +Q�H��&��  H  2  org/bridj/CommonPointerIOs$CallbackPointerIO.class  H      �      ��]SK�߁ȒuEEQ���$Q~K"NjbJNQK�6�l\�����?��B-�/����(˞�q��)nf'�=�>�=��~~�`%��[�T\����;�ˎ��c�w���hT��Ф�1�r噙R�1U1�Q���.ox6W.gg�{��o՟\2V�c�*PD0��Җo�ŔD�Lð��D �[m�	r�my��&"ǒ)Y����yV�p #q��A��)\n6x�˔_4y��#��!V��T썣G)��Ԣ.�v3���L���s��&�3��;���\��v��l:��kM�����U�����v<��t�mW�CoR���]�z�2M�r�b\gY��i�*�]]�\ˮ����B�8��z�DW�Be�z>�-�f+����H���>���'Ω4�	��;�@A�A�50��0|=�˰ǯ��P����^�9�� ��.{�ܵ<�{�^qj/t�=�K$�b4ڜ��!�?�M�F��R6KbU��7�V��2-��#�x��m.[$TC'E��V�6��K��N�������k�/�E<�MF��t�,��o/W�+-c���Kt�d��[L��;�} �"����*�m	-�`���Ex��l�z����O߿�W4�ҿ��>O�:b��S�w8��q$�����d��?��n�	����7���>�|�i���k�c�����Rǥ�K��7��_���g�Gά��F:�z��5$�#�&D����%�󘤄b��%�@%B(ua��+�eCB�%/�/	�J1�s��sY��)W	Ԑ@�bw�(n>$VCU�QW)JP������h��MИ�"h�TZ�Q;�0�v��h�J9ɣ�&f%�&}OG�i&pKj>�cQHss[��rJ(�H�����A��(����[AO�tSPK
    +Q�H@�2^  �  7  org/bridj/CommonPointerIOs$IntValuedEnumPointerIO.class  �      ^      ��[S�@��K��.G���� ^�V+`kg@x��`�2i��pƏ�3���W�Q|�/�x6YRڦ(�a�9{.�s�|���#�I,1L��Bb�ж��r�T��5�T��re$��kJ��n��Ւ#���R�3�meWI���
����lr6Ws蘤	�
�$C��L����k��ej.Abp�g�R�;]T*���,�4�lH����k�,C_��,��0�"I	�c�m5_T7���5�qq&�>�#(Ç�.����k>�z:w��0u|S��T�!mnm2k��d;�zh2�p�����͜���Wxo4��8���8[g�PT
+�)�<�0o�KV(^X����q}�%i�f�/� ���u�C��o�{,K����p-\KD>J�vr�h,+c����
U��P��h6sq/�*��"^g>:�pK��;|����4��̎#�I%���	�L򅰃����Ԥ*#�!��.u~E+�Y5�8�tyK��˛JqM14e����_�:!�3qЛ�tu�Z�P!	7�f�.��.����w�������
׷R�����3��VBj������(��G_m�I��o�C�y�����%������"��ا�>i���m��l�9��쾵�����FѾ��:���O��K��hNE�}���F�;D_:�#���>�F�	�]�9��� ����/[� x�B6@��S/�qc�V���rBBH ��n�ޢ�r`B�֚&-���~"�_���fH�&�G#a�'���jd�&���Y�$�6�&Y��L��|��ả����Js��.HN8�	'�p� Rs��S� g�;��*�.h@���PK
    +Q�H�nC�  d  6  org/bridj/CommonPointerIOs$NativeObjectPointerIO.class  d            �Uks�F=
q��!��@��֏&Nx�i� 4&�	�>[	Jmɕ�4@߿�_:ç~�L;SSf�~�j{VRdǒ�����z��{����~����0nZ�5K/o�f�j�4�Mݰ5k�XYRm}K+�mj%�ߖ!I�0�ty��j3�Q��K����C!6��t��m�[�����ɐ*RB�V��^�j�����1]�7��f�m��jtL,
�\E56r��^�!',T�7��=%�X��S���Ѯօ6�lE��� ��QD0���S��� �@qW	��_��J8�*H��+��X�WX��iتn��-��յ�V��{
��D�"�R��n4[�jW�KZ��MC�k�Z��ҍ���^)k��	{Rn6�GqoH��d?Ҭ�Z�iF��6.D>��P�
�xS��vDz}��Ȝ��0�ܩJ�aXZݬli�-�m��d?�H�M�5N��z���:,'�KQ��[z��:kq�e���M9�ґ:X2������5?OF�m�cAƻ<�:=��/l����F1�9	�]�mwi�H\�;Q��{
��%�>~��y��>u� a,|>�t�ǆ)�e\g���s�.�����T�k��h�`5��)A��4�p��\H��Qֶ��#$�j7	�q�2����TW�\�c��'<v�+E<U�U�&|K�-�����T���h�"�)��V�Y����8Ş/K:� ���R�ád
>����j��Äx��X]+���
�X�_�zϚeM �%���֮���vo��<ClQ7��FuM����^�nX\��S!��Dw�N������[Y0�r�4ZI��s��՜��p���B����s���L&�#=š�a~�!w�d��X�N��S�q��s�����Lc�&&�r��ŧ����C�qy�8+�,��
g�6��K�E�Q�����;���C4Am|V<�sD����p������ߣ];;,}��y"����b��,t�Ep� �%�W}�{�q
��1�f|MT���� ~�?}�_�9�0,���<K⸸�xf�3G�y���,��љq/�X6)
���7q�� ���s��6�:1��K�G~7�<R���Ze���8��k�����UtFb��>��x:�(7q�v���9��u$|	O�X�����L�Bk�іqL���6����C�V���]��{��90M�U�x��+�(�lr��/�M|���2*�V��UA�Ӫ�F�~�#S��&g[�mz\��Mlw����>��ѵH� 	����[g��w�����z��?PK
    +Q�H���U  �  /  org/bridj/CommonPointerIOs$PointerArrayIO.class  �            �V�STU���.W�!�R��.�j�&I���BB(���w��ݻ
V�V3}�C/��LM�S36�:9iߚ�?�S�A����ea�:6�s����{������z�>,1�e��ؔk'�b=�t:�elǳ��`v��v����T���#G��f,e:����9k���X�R���^�GF:��a���
��a#�=<CSy�*T����2�9'i��Eۙ��?�����ɠ%��d팓eL�3�{�L��Ҧ��^;MF��]ե�e���f-��ƽv֜JYI��2�c�ܑ�y��@��PךI�1.��o+'b�+��bC��@�v��k&9�N�z�3��L�L[���d%������:�Dy��e��h��c'�a3�X)�����'�xB�a��F|�P��O�Q%�\'������;We��}�._���C`G�P�vi`CGYbE���Bgۨ�0�r�th��&��؄�|���:���!O�i�9[P��D��l�s��#���6�>�Ig1)���p[������_dP��))!� >wR�^��Aeff&�-Ca_5Ǒ��*f���#�E���In{����/�L>�����3C�Me���W�N5�e>
�CTm�c�dg���z�{u��n��� V�Ą�q�Jg��/��~�;��MkN��&P�´5�㨘d�������l�F���Q�if��hw֠�v�}֐�e��*L�s+��aϥ�&;9��1Pq�L���-�h�)�;���7x��Q���e_���-�g�i�U}8���P�N���e�+U��2iem�Jj6�^.+*6��.jȁ:�z؞uH�R�JO&iq��i35j�6��#|�(�c�ʥ�,Wބ֫�Đ÷��Dʩu�G�!����V����ʉ8,m8�s��c6OCO8��
J�,⽂��@-|`�D� t:���}-t�KC�>���YÇ|ܒ�[tZ 
}���`WK����Vߨ����`��]'�������ߦ5B�
��J^��O�I@�xd�-��.���	���t�b_�Ar���P�G�D�#�\�E�nV&*J����%fw/)�o��:*%�!p�-2e���r��M�CX��u�{�ҿN�H/�6��n���X$���s5�t��E,��`$����e��,�p���.�,#�#�����%&��w^@��k�����*���7��֏H�c�	1�)����sY�+�I@$���"�V�s�����2�i�*`��I�U���Hb�.��$�wD�p�/H�K��c�T]&:+E��tH�!�^��|���		a�e�aQ�JZG�W)b$T`��,�c��,��\���J�KZ����s���
5�0>v�=�I�2Z�Z�b2ZK���J�=�h�J2��.�̱��;�y�� �A+�I�n���"�@�&	�k�#-��R�� i�V�MhlI�a�h�H�خ�����آz���ģ#-��p��xt)[c!�"��ü�yF��b��]�>�N-�Se�� ji�,&d�6q��W�`�T�l�g��ٱufA�L�o%��P�jT�PK
    +Q�H����  	  1  org/bridj/CommonPointerIOs$PointerPointerIO.class  	      �      ��[OQ��
uik�Wzx�E@-V!�ѨO��%˖l�|�?��j��o&~(���V�Y�d��̜��fΥ�~�	`���]ͮ�Fy=;W�بY�5�rt��T?/��EcXȗ���ږ�55��]Z]�ל�L��ǏϷ�Rn�~��	
B�9.s5��`R
Cl?.�ڰʺm�V�� 	eD
�2t��pf���驧G�
���6�zŤ>eK;����}U�)i6�����<<������ �XK��fv^�h�Y�lmC']�^�4�3�nr���Q2(�� �@�	c'B+���b�z�i��@���9S�ש*�p��wVEGzс��ye����ؠ�k6~�I�I����,pn1%12�i���u�*�:O�I.ʷ�$��.��]�ʦg��{b<DR�.���6-�"�撥��Il|7���R��*�����D����}CAEu������*��iw�f�؞��I��"��x�d�z���H!��әY1���4l����:O^[�̧�mh��^�:�{����#Z4,�IccU��eTzqx��~?��Xuَ�mfᐩ�\+�Rk�k�}�נ,K���ב�^u�?]�����>}u@%+]m���Yޠ�F�X:�=��{��c��?��41��'?!���\:�>Rh'�sЛ��H�ȓ)���>�|�4��|��� ���zD^Zaed���L����ϸ����x�M�ţ��%sGS�BiZQ�GM�n7��E���+�ߒ<�]D������Uzڅ���_="��h�l!�ã����E�(���yuZGP=��U�"9UEP��Lb8��&f�3�>��;�I�]��b��*|S�#e�LaNh>�h�W!�&�/���)��"�Z"J���J���ݍ%�tY����PK
    +Q�HݓZ�0  �  0  org/bridj/CommonPointerIOs$StructPointerIO.class  �      0      �S]oQ=�����T[k�@売E߄��CJ�%胉.�/Yv���D��&U��(��.E���>�;Ùs����~��	���E�(=[�J��,�����f�ɩ�=�� �1�5�I�&��{C���zk�ّ�0gp��V�U���
%����v�1�\�&AbH-FN�6a�:>�K7��n���#5a
�ΰ�?�P�2d�q	)�P�;:�ޒ����2�2���pWvW%l1$�*��cN��Z�JC3���4����w����:��/b�2�؍#�2�cX�M�t��p*�|a�gO}p	�Ӻ5O\��lo8��Z�^�;��ʸ��7�}���!戛.��L2e]��jX}�ϴ,]3��-��A&t��<H˙R-a�ɨ��)S�[s'6�q՚�:.���4Mn7�q��[��0�=.m��uʓؠ��~����t�t��o����b�+���ԇtgY���3b(S�Šv��Bg�T@�8���k�p�i�����S���|��	��6�9��<�#o�4�´�?��HqHq�bŏ<���E�N�N�?PK
    +Q�HW���c  O  6  org/bridj/CommonPointerIOs$TypedPointerPointerIO.class  O      c      �V[wU�N�f�0��\������rQPZ��mm�,x���05���	T����.߀%�%K�����.��]�/��Nr�ܦ�X]��>{������L���� ���>��-����и���س�e{�;9Sؕ��b.�w߬A�=��F�:��,�Q#����a�kB����s�����i�HR �q�@,%��;7�ټ���.xn1�9.�+���Q`������.�m�ԄG,��F6&���ORm�8��1W<˱5�'JS4l ���bR�&l��Fl؛� UO���DOmئC�Ch���G}Ѫ1��9q2H��N�xDF>��tʙ^M�&�4��O�u<��"�a���IR�lm5�D���e��H[��s�kٹ�E+�(K�W�5Q�:� �	�7l���Y�^�g���,��q��2VVL{�����u
����q<!A	h,ƴ�lʆ7G��I<%eh���Uǈ4�i�d r�%}�u�yS����Y�s���
&�`�;kqn�t#��ɠH�(xi�eA�'���:���g�8&Y�sF�h�d�Idt�(��/"���li�f_g��'i2�{��nB+�uV&/�D������e�>5Z�4<3�΋���{t�p�bVL��CLq2�5L4���-�欋fz̛�f2G�����^��(xC��x!½�cQS,�6���m �6�9P�e��@�kє�Z7��{�jb* O�M��%��-R)��p����l���@��};PB�pS�pVV� C����̉5�0Eg��yA�c��نWt�)4�,�2��1�'ג;-/�Rg�V�Й�ls���`�����e�tWv"̪�+�@��bk;�*sE朢�1�YT��m�E4�S\/��K��|꒟�S�F��<����.-wF+��%n`����Ɂ��M��Fl��v͕����g�y�6������-��>X���y+at�-�}s���d������y��3�(ƉG��OV����_��ע\���>�~@~��'f���f�_��7��
��ߔ�ϩ)��X��O�&�%�@�z��[c_b�������Z9�P�z}E{�"�mG/I�
��+ɲ����0��J��{eM
�\�(��;����2�_���>�9�����w&���U��7KX�FS��}�Nd`�!;�%����v�U�^�����?
��q�)�+�*�FzO�����>z�L.�G}��B�O�p�w�g�yD���M/�(R���3qW���k�=]��d�b�'���բ�2�	��6�k�P��=3���Y�Wg�{B��F���_g��ZE�V�9�Wju��y�
��e^��%\ll���i>��� Z3�+�k�G�{W����ɹ�@�PK
    +Q�H>^�N�  v     org/bridj/CommonPointerIOs.class  v      �      ��mSU��7.IS
[��BED�(�BA,��Hk���$KX�٭�J}h�U�S�Z��:���茙�/��rƯ�x��l�n�I������{�=w7��� ��3�q��G3��[�ƌB��/�n)f�b��14���rT��|�bfM�ZZw�c|x����5%���a�ʶ�%�!�lq�Z������KO� �ѽ�1���ɚ���W=��-��z}���MS�)34U�1��D[��2}>9��Y�Z���w��Ԃl�늳ݞ<��N�y���'����5�A�v�6d��	b��I�,�S��(�����b��ן�8�O��8�OPQ���E�[��4A}���db�L�QQ�91Ep�f�y���VT�@;�WӞA�VLR���d6,e_�3C��]��#\+$F����%�͐�7�yA�A�9�����֊��Q;,�1M�u�|�\��:�L�ו��$�m�	J��}٤K�[\3(������ZS"��a\@<�:<�Pg��E�����TTs2��	Zv���T�SSY�������wc5�X�pf�R���'�� H�]��99CȈ�����9^�_0��FU�{o��'�1�2٣�8�SQM�V���g/�.L_^N-'�W�X<kA��j����\���ݏ�B�̤����N�q�B�Д�SUj��8���)���>}ݎ��A�*�Ƈb�7q+�4�}\dwǧA��	�:�U`�ٔ���+�6�;�tr�j^���IU��9Q̄���E�TeZaJ�Q�+�BF1ݑP�(�Ye^&�uŴ�D)ҬԦ�A}���0L~��ϐ�����<~��9�� ?��ϐ���gɟ��i�3#?��s��=�9zA�2�O��Ii}���|O�ag	�H��Bv`-�o4ba+��D��_+LK�8{�d/W0����ɾRƕ
���k��^/c����$ב˔�� ��V6��/�aTН����2�
��Һ���26*�LK���������ts��]�'�HKw6���������tw_����{b��^� �X M��~��3�qvq��؟Xa��
p;p�������'�{���5ҿ(�A�C�M�ͤ-�GH!=J�(�1��mv����p���.W�]����j���:�?PK
    +Q�Hkt���  �    org/bridj/ComplexDouble.class  �      �      ��mkA����$�z������ۚԠ
Az�`����$K�p���^�[� |��C��wŇK��bgvgg���?�~�M¦�'�a���΁����@'�P�A����c'#s8�ʑ)�!����p*N��\Eʼ 8���G	e.�\�V�	��府K�/���"�:��ǜT<a"VBAi�z?/�w�����%p��.ޗ�A�L�Ɋ�p�vs������ᡊ�MZ�4R���;�;�m�X�-q뮚���?�=�c�-��H�+��7�V�*����P�g��Q5�5WxE��tē��u�XQ(Q���v�(������Þl��K�xS�[?��2�}^�4����Uβ���I�^�3���)�>����{l�y_��õy�pQ;?C6Nq�����ޢ3��������R��>�畨����y������9�O�?;�D#�PK
    +Q�H8Z�  7  #  org/bridj/DefaultNativeList$1.class  7      �      }R]OA=Ӗn[Y�|I�Z?h0Q ƤФ��"/<Mw�v��L����G��?�YM�1���2�]�&Hv�g�s3���<��2Ê���/�nyO��6x(��.���6��.��U�|��
'4�d��&ߊtK�T4�fX�i�B��Q�h�2���r�+ú�� C�s��6��Xl�_�!qR��]ǓJ�����1�ߧ���S��s�}_S�i���{0�K'����1q�9dq��$�f��<��7R�'��ۓ����%JѾ+��	k&V� *��0Y�g­�>wd82��2���^��+O%oy}X�K����͗�aHU�K���k�{�܏�E�a�.�hz-����k������t U�@���$5��_�x��*�R������y�`
a��G$�^������7�F��wR���z�5�c�A4�/���,�1�<ְA���xA��c*\ E�p��^y/�yO��!>��)axF��Av�NT-1+C���|�pPK
    +Q�H���[0  �  !  org/bridj/DefaultNativeList.class  �      0      �YxU>��d7�m��I�m�m�٤��RMK!}�iS����(��I2t�fg�TZ�
�S���B�@�T
�KQ�>�S� T��Lf7���}b?2s��s�=�?�9���S�?t��N�fHT���szu5vќ�J���+dCV�դ�!I���]-���򜸜���{�5�-0�R���ڛ4t9j��]]��k�(�h��2�Vɉ�6��*��<���5z�-Q��B�ٕ��C^��yt
KKT;����y�D�i����0��W�6)� Ѥ�u�J���m�WM��5��U��2_&ҁ�iN�&�y���&�a}j���VwR�Ӥ6쭗�IE7T-�\�&�޸��Z�|���r��P��!~�BS������hF�8؎�_;�֋�	�X ��!�S��q�D�P�j?5�,R&e��Ǖ~9ު�����dcTb�=�hJF����D��q`�}4�5�.�	���BPzi�����@�j��0�1o�R
�N��Y���旇>.! ����V$&�`.}�Gg�GaX΢�����T���
y��[-g�ͧ��Ip�j���g��ߙE��b�
��C(Y
͔��2>e6E�J0����&j��ق9�+�� �8��R����W���~�g��H�D��!pJ.?���}TF��TA�L�.?��d�DeиZ���%q����j���ho[�iT����%�~�S�T� ��݉A���>�z'҅���םH���4�PbC�.3��+Q�9ez�w*K��b>�2X��r�ߴHN�Z��K�$��P��B�}�����-��U�TT��^/Q٫��cc@N� |���Ay�:���lAQ�Bm�Dc�(�fK**XTC4���|cޠ˔N�*�1��JD���O�4�C6�Ѹ"�~��}]�� �-Ҙ�d�ff�DL�ؑ2:�j�D,���� B$1�<���^��F�w�3��Vl�D��d��.�_��t���`$*��fY�O�g�h7@0���ͬPd�����5� '�����f>���P����V���r.9��רz�M��\�Ru�S�0n����I�8(���AmXY��P����Nu��k���:���|�|�nc���V8����>�k5�w��E��C�PV/�������E�t�-&?}�������~���}HݻE��_a���n�;Pa�x\��F�꺼��p�5'�� d?�C�jC����}���y�a��f��L��Q ��U�M��rگk���.���<��P6f�|	e�}�{�Ü.�b������M����f3�ݣ\"�E�A��5}�	]@�͹FÆ��#r��Y� �6���	z��<�j~��Z��Ϡ��ȷ�v4Kt]���������;
�:C�z�!�!P�Da�:k�1��^����rf��Oy��ph�oG���fp�y�O�2'~]x����?SԼߘW�o!��i"�0H(J��#���t]ID���3YT��Z��/�I�j#����6Z�0G�������&��?p���=R,�����Xѱ/�ЏE9R"�N+z������맷�����ST�����i��&�׬r>����hn�9�	���_*��\~pO�Q!g��V'u��Û�aR��{�(����Ώƭ�*�$QPc6�;�H���Z�4Q*E�&�ITܩ��L�\xi1��8X_-�i�2{����(�Bi��PV�{ݚ�����3�s�"��ϱ?/��)\/E�6ǞP�W�(b����b1x�XAf��?SCr����SK�Qe�*�H"��YV�M��b�˸D�/���.Ǹ����ܱ�- Ħr�\It�Q�Ļ[�K�#|?M��T��ߜ�TO$U�����*���L�y�4�:�R�*�Ʌ�`�056=N��ct�5���k�)姦�C�4������є�%��bЌA���������y���͇�'��u��p�!�~�6?hn�/F1b�
�KU�ǔ�iK�;7��x�7���r:��Z:=�*�s�h�,ǧB����kp2�S	<{�|M��r�0�=��oe��Y�NN���|ws#is%"��;\WA�=4c����f@xԥ�b��~��}9��mpA$12(��=�<{. 0쮌u<˞sa˗����Ӵy_��%yΖ䑩�Kl,WXX�@�-�b�9@_�N_���aZ3��O�eAo�D��z+[�my�wќ�¦�au��*���
!�Y~���r�ToMӍ��1�؆v1��	�d�[�g��x��B)�O` ���[v�h��1�?غ�!Ŷ���6��6�/���2�@_��d�ɡn;uX�V[�VH���V���}	��RZ ����H�+,g��6�r��������	_wSq]�6o��'���|r���Y���:���<W���=bb6c^#������-v�l������-
���;��p�*T��QE��]�r=R���F�r���N�[`�Y%���z�]^�.�,��,���]^3D�.�X�7�6���� +���/�. C�E�8HwrQKӾS���Z��lK ��[�r�p�䫻���Y�Bl�� ��"n�@a��	
Q���$Q���Q�xɔ\JM4�]����a�p���m�uz�#b�kJl��L�c2~��T�m)|]	o��n���P�nC}��x��	`��m��8�2���?�yfe_w��=�mQ�ʭ��Un�H�C<��Δ�v�"�2|�����TO���;+�)+���(%͋�Nh������oB�=�ҽ�|��D-N8b��8��z�\Gϭy�8O^�����tV�;B�,�]���Q�ܮ4}�5�`����8�ǝ{������Ӏ=:"�� ˂�,̢4����#(LGp�>���0�7�i&$<�jq�gwДڝTR��JkwS�=���h��ܵ@�G-���'-��B�&?��Nn��/��蕖�@�1�TЫ�Eiz-�п��][fl��Z���u4qb�;��3Q�ܸ�L:��)҅>��	L��L��-����$��<���O�AOC�:����shs�G'�l���.�J�7�8v���D�h{5��*+L���o:� �Q��|��x�զ`4�' zo�$�{/�]�W����GW�&nC�N��/����j~�ޓh+_\������\�7�7�5���M���������V�7����~��V����L��Ɲgu\��yQ�$wZ*��.(�k�J�~Sh�X^_hU��,�Mi�8�����I>ɟU�͵��Z�ը���e�SG^i��@6�5�I�ii�+��ѳ|�do?F��K.)(�>i:�����2/p+�I��PK
    +Q�H92x�  �    org/bridj/DefaultPointer.class  �            u��J�@ƿi���hk+"^�f�`�jC@OA���7�7�D����$x�|(qR��3��?�}|��8�6a�ԩk5ϼKy'��ܖ�0R� �؏��L<	/E��ęL�$����̆E5���C���
eB{|4sac�A=�e�Ղ��r�G�$���VNpӺ(�0�D�3���sՉ�ӄϏ��~�
y]=�R���T��0��ڙ��N��%�b��#6Ϻ��9kM:ǯp^�h�����X��A\�-����!k�7GK�~PK
    +Q�H��qM�       org/bridj/DynamicCallback.class        �       ;�o�>CF���t���̔,}�ʼ���d�Ĝ����lvFF� +��ĲD��ļt}�����k;L!Ft1vF4S�@�X
r*�5�1���f<gpfz^bIiQ*#�V]!A@e\���Eɩn�9�l�L� �������� 4�cb�b���L� PK
    +Q�H�,��  �    org/bridj/DynamicFunction.class  �      �      �TkO�`~^��Q��_Ԃ(c&*(��e��&l!!~꺗�еK�P>��+���H���Q��3��ؤ�i��9Ϲ�����	`�Ӗ]I�l�|�ܿ4՚�����)�1�3G���z�&լ$ߗθ椳�vԞj%U;O3D�Z	A��[�k�A:U5ǲ/�}Y�<B�q�j�f:��� F�C�&�2��;Y�@l�8�aDd�p�!�T��J�T��Q:K��]�R�u�8/�>���W1��uŪm}RK�0��!`�a�_E��&ݼ��9�V̏�,"����i�1��m�t
��h�����8QoۑG��k�����>�3L���`*��(s[�c���s9U7xYq,ţ�h�]PRJO�� 7i����xp]ܻ2P	1,�$�[�=��G���U��cyFZ˘?�|�x&|�i�{���f�۴2�a��2��t�5T�
��h����P���U�YG�5�X�uY�D����0��M��Q+q��*�Su6=O��UZw�`5l��hf�yZ�����hG� (>%0���$#�_��7ל�3�)1��$��4�Hf�]����D1J��+i$�'�xpu�҄r���,�\�It���֚x�r��_.��7�"���s��4���[��&�� ��@����!�6v�>�!_ڇV����Âd��[��}��;���=B��x����PK
    +Q�H"9zuQ  �  &  org/bridj/DynamicFunctionFactory.class  �      Q      �VkWWݗq_�+R���� �DS�B��T��N�ILf���>�}����~ծ]u��[��������DH~�b1�r�9������׿���$~�Yv&����b�ʲ��d�h&�2#Zұ�e�@Ϣ������	M%���K`os���X�_C_/����O�΂�
k�l�L[�E#��m:z�=����E`K�2�]�N���t���5��K[�M�$bd���rM�*9�j[�y&��k����"F�Q�4�1���:�pV+FZ�M�.}#�9����m��Y�C���)��./��-н.��vFw��|���nH5�	�
�b�د`�.�᠂m薳C�Z>�]8�o]t������7��������n,�  �#a����Z�p��
Xfˀ���!�PqLA��:Bd0o�3�b�֒�Dvw��Q��zfW$��T�gv��g�dV��9/���9ь���9�� �A4G��ҕo�׉����M��X=��5'�&I���ti�g�Vo����|[�ӱ*�$���B�q����I~M�:R�iċ�x���%y�Z��@�����K��,<��ַ�ڬh���e���K�氽�0�\�ƥ���&�i�Բ�Cv���8�1n���D1חt;b���R�>nva�<�4e��E%ݷqG��vSS�-�-I����-�]v�8ؿao�����5=���K
�"�ETw˘�y�y]R��$]0�������xҕW�C\��TY*��3�ae��꼊,��1ܨ*e�)�hEC}k�EE
e^��h:c��Y=���B�3 �G���'��L�k�Ș�S�y,��;aQ�s�mH���O9��������	����\B��+K��&����(�j/,��9���;c�1d!J�4u�\�^�!vg7��q�U������[�7!�{d�(�z�ǽ/9���n�ϰGr��@	V�S�+<,�Ȱ[u�����y��+8����~w	�_��������%����%\�w?õߟ27��yp�Ì���H1���.&�)��$�@y6���)g2����:f���Juo
Ӝ=�\���S�9C쳌v�Q.0�(c_d�a�c�ť*-_�v��$D�,1{~ƭ�~�������i���j̞j���ʬ/��q��W�gߔ�e���]|TE��k.���?�.��G�I��2����rqp٠�+�d2؄�`�٠$���#�ʫ�;�y|̨*|e^%s�U^c�aгơ\)��0J���D�⍜� ��(��/��go�p�-=���+����<R�Y-�~	�x���Y@�眳�'�=R�lGy���+[��{�^�z�ű�?PK
    +Q�H羵  �     org/bridj/DyncallStructs$1.class  �            �RMo�@}��qbܯB[%N�i9 P�^*!��H���^��u�v�� ���G!�vC���Ͼy�fƿ�����{��]-�Q�7U�~�'^5N0�����W��w$��@~!�c(U,t���6��P]�:JHvV�2PbXw'2�{�(�1�l:s|���r�PulgICǂ�[�������9��\O�*���7��P�+�^�l�B����R���!ߴ�f�����JFug��;�Θj�ڴ9N4Mg��n��h�X�ぉ*2X�w��ȪYx���-<f`c���|�:#A�X��n�ƊR�%wq�\��T���+�u����g�r_�'����M$$-��p�=q.S����H�ᅈ�B�:{����D�c�h�	��sth����6YFv��;_��&�V�.���t�i���P'T�|I6�3+߰�O�|�P�^����n�cO"OɳS?A�Fop��xN</R����Y$ėO�@	���b��Uq�X�PK
    +Q�HP҇dL	  >    org/bridj/DyncallStructs.class  >      L	      �X{|W�n��d7��l��Ш		� ��<H�a!�����t�;�����Y ��V��VJ+jA[�J��U�4$EK�*
��V�������o�����浻��GvΜs��~�q���K?`	�+0;nFݦ�h��U�h��d�J(�;�]j�Pc�@[�N-l)��9Ys�T�8���%

���G���ݦjT67%�
��/���#P�^#P1�������u+ܫ�D`�������$Ϸ������[5CS���L`F�\�,�V���3C���3�kB����4Q�F���Z����N/.�
0W����<C(�\\bś�=��b�����:�s9��mD����I݈�#��j�q�j���z���c��Y�<-�}�@�j$5fZ({��x^��4T	(ZL�6����B�H~����8�`1��jVC4jjQ��"-�fD�JYUu�Nᤥ�������ă ����2ˈMB�A�az�+���h����'�E�V/�P/����Q*��7k��S ^T�̆����A1=Pd0�D�w<��Te.Kͬ�{�-��2����~��R6�������M�7r��0�㾶*ע,;O�Yf�&l�x�1�"�&#��҈Td9���
l���s��팈��;�f$<.�e���
]��v`�\�Ǣ�2�e_��5y�c�/������L#O��a�O���bL�E1ql�Wg�R�	��n�CX`ָ�6J���.�Yqg�@mN�37��(z=�΄�w���W�z�������'��	�s��%��j,�O�"i���?-��==��_f嬪�X�bR���f���ٰbY��J1�b���.9o�jFe/��ok2Lؚ��6Z:5M�Mڞ~��E�l*ҙ>�%����=�)>��v�$��;�2�
nf�U��=N���߅[��N��G���� :�+-��I��N����G��^�ou� ��>,	y0������������v?(�������8��]8� Ƹt�&��L�`�j�%���ò����]�6p�q�%��l2�[�*�V�ý� >N�j�/{q.��Y�i�!-�z���ÿҰ�/=�<�aa�6
>����w��S��!�pH���{��`rL�$ئ`�N��X�Rca&ܺL3�ȴH�q҃�0"#r�����Ԟ�N�[_��l��s��쒏p�6H��쏏2c;��l�4�_�cn|_J_��0�E|ō3R0��޸I����Y)�9�^/�/lV_w��)ل<�ƓR0���x�w!3�)7���Y�W�ٷ�xFJ&L���$c��n<+E&�0�f�3����aOXK���������?ljlFc�ҹ0�=�D�;�b�xq�@�e=���G9��=��ă��S���Pr9�t��<~.��6�D�;țvV�!�g�G���e��㠫��/g폵�s���l��T�N�ҫ��J�V�NJ3���I3M�e�8A�TM]��!h5�Ǵ�ɾn�WlN�d5:���i�Bg��/`.�0��ϥV͉��O�a�E� x���f����I��� �]��|�H*>���r�J*���q-<�K��*��ab^����Whs�P$����4��g�<������5��)�\:��"�Q�WS�F�<Q��w�CXt.ql�0^��j��I�a�F�t
J�I4��M������tP��Fo\�_�:xu�p5�-�n�:������F��M$*\�J�Ʈ�p�8V{�~�۾/���l�|�w.���x)�丏��'�G3���\�u+(s�����ȓ�_JL������K�����`5-��:Zk�F4�vn�\��ퟰ�j��UDr���v�6/ŭ��>�Ł�_������~W����pO]���JR�G����)R�zEQJ����}�0>{���6ZW�+�)���[��:*/�p��-!��30N� �u%����>��|<����A���_=
�O);#���>$���'��8���u��J	�t@
��R��������T
K���;����m��=����F$w]Yyꠞ�~�X|
�u����yz;�~,Sʡ�7'��5���|i�8#t��v��O'��bL�¯�k��F,�o�Q^�R�[�@�cԋiJ�ƨ��a������Z[#��~�l\.���2W6�&���ζ�՜�^���	�Ɉ�8G$�'�u(nş�Zen�/D���")Yyv����b��j[�7��7������ߴ��y�!~9ob����
~�m�t@'e���"~ۉ�ո��G����A\�	G��ҍs��)h<Q���r����N��A0���[�����}H���B��R��/��ۦ\��R=��M������~6f򳺢��?PK
    +Q�H�b�hm  �     org/bridj/EllipsisHelper$1.class  �      m      �PMO�@}�j�����p�z�x1�T=h�xZ`�%��l[�^41���2N�	�̼�˼�7����� ;��z]#�c����ex&ԝ0�6Þ?���S\����=�o�x-����x0�q�`(��o�bX�=a/�dX����͐?�ZFG�j��b���h$C�m���MԒ�W�`�Tk�g(N�6VJ�ڏ\vǢ5\�� ��h}������F��Ib(�R����+�73%��G��ڹ
b��2mm�
B���"}���Z���a(B�Ӵ����3�a�*�����p�ȠB��"��%�u�|�Ta%����Wf���'$^�����lq2y#��b3�<�-�QަHVʤ+�}PK
    +Q�H�]��1  �    org/bridj/EllipsisHelper.class  �      1      �V�WTU�`�0�@T|�$j�! )(8�A�����̥˽ӝ;(j���ʲ���,{`o���ʖڗjUk�����׾�V��;��Z��s����g���ٛ����	�_3,׍`ՠ���ZUU	G��N���!�1,�G�*UւU]���oJ�d(LgV
Ê�,�����P���Me�{u-bʚY�+�Q�3�r��%Jp2�&�RHW܈0,�\�	\�t��60Tν�8`�k�^ծ��ѡ!n44�Bv��)fC���ׅ��w"YfH��V��))/�j����u�RπofJ�:ۅX��,g(��g	+ȫ 7�xJg�uaV;�w��9�'��P0{C������9f]�݅�X�D	�Sʓ*�c&O�x農��k&oQr�
��>�v)69W�r'JqC�IͰ�3O<*Q%60�B�GW4S�^ð�ǑU�|�����&��"��p*�t2
�uTd����B�M�M�}�����Ʌ��gS�1,JQ�C�A����-9Nn�ɭiϬE���v0����v�ޑf�M�e���-9N��]i>�dH�_�,�8�ۦ��ŢY�U.kzE��(��П�
K���o�e@8�'�
��
���Tz��üG�+*B��m��r�&k�c�CN����]C䃧c�Kɠ+v�	��鵓6"��N˚nvB��ά�D��\��/�����(Úiդ�<(�ۍ`t�kf�!?��N!=D�jZu������hd;qD�����ۤ�uk���Z@����GeC��4�r�E�A�����<N-L��`���f�P:k)~:���<5C3�mͣ���<ΐ����9j'Ԩ����$MW�I�$�������6%���~�<�g6��5\x��x	�0���F'�����b�ޤF8W��~։1���t#�h���[����m*�p�nf����w���X�fQ&�
dv��=����("sLʙ=ˈ����(������k6�UkD9!�Z��V��lF�"˫�pC̋�x����O�xgtd��g�5��M�ծiܰ��#p� ʢ��81���%�,B&}i(��W$Uї��Q6�«�
���E,A}�z����»�l�����M�8�;o�._�ͭ�5��#�"��W]B~y�*)t��;37ge���jˊ�j��b;����ț�����,G�-n$�n��v���k�6��x��w	����-�G��?`��,p�����{-�_����z��l��qrt	����=�!��,�cI���d��i�<(ln����8�?��O��t�#�gNĥcx�Ă��'�3�8���f�p!����g��+�$�s��Q*�G-efoRR��Ѥt*)]HJ�'�o��/I�Oʺ-M%$�N�ֳ����`=T'�Z%�Ç�H��c���N���i�|B��g}���-QSg��*A'6P�VSQ�`56��ln�f�u؁-�"�؏F��:~Ҵ>�m8��8�f��i(���j���y;�M�_с߱�����؍i�N�t-���&j	��.�� j���O⁔���_�H��/������R��C�	+5\�oI���C�%�m��PK
    +Q�HS��    "  org/bridj/FlagSet$IntFlagSet.class        �      }R�NA���"���$#&J�
�b0�=@�p`�K��,�$����d���=��Ѝ^fj���k*�����y����ۖ��/ѫK��ʴ=n���Z_�D�f�X5��r�Z��*5�vܘ��]Ma8�;�V|�(B��?dQDq�y��b3��HY7u�B8<��sza�����Th��ba�	!�N��o��ab<�/�	�rM�k�&y�끐�mk��/!9��<�b:�}o��Š�S�AGMa�mȆZ���ǇI#Y�My�ܷ��U���3��X����v��B�ï�#/u��_���\�"� �J���bs*h�l���a޵���f�K�|b��c&r	,.ZA��
���,�2�`�6�=��@�㧱:e�3k�q��X�v�e��s��K1ɵ�A�PK
    +Q�HG=H�  m'    org/bridj/FlagSet.class  m'      �      �Y\[�}���2��#� �vL��O�m0��)v�L�5��U��$m�-k��׭���vMV7���;i����k�u͚�[�-��u]���=�~�ܣ+�{!^�_����������?�� �D���Drx�@2:td��Xd��Hy!v7�n�89Y�ć׶�'F�{[��5m˚�?p�L5udD��&���n��۽p�8�"_ ��X#�	,����-��4-�g�x�Ii�]���̖Xd|����ZMQ��ܹ���J7y�P��>�턗��["�#��on�HEck;#c\�4s�ن��t�N�T#�9���	��i��oS�������@ 7��*(���aI ̓�� "(G!^ 5��u�(NQl_�l���J��ƦY�W�Y3'��T4�bu %(���
̛��u�ΰ4�;=��� ���X�E��)G���V�Qы��-:��HbH`G6DO*�� X_,k&i�u�)���я[��|ζˋ-�&a���D2�{r�S\Sk
�[�hm�L&#'�q�;%�.%�$F�q#���x�<v+Z��c����xd f�N&Fr���=�+ϴ	Td��'�訑e�}~t���F��G��f�88�����_^�6^jl�&�� �Eu�G�W`Yf�-3�#����Q��u�M���5�I/��G���b'��!�#ccF�>���#��)-�������9�p�Ɉ<9 PJ�x"�3B����@,:OER����y�]�QCZ�.��cXZx��v�=!3.jjC��)��pD��J�������Än�5�;�L���d&��}c7ұU1{�0y�{�P(qʍy�	����śr���<��4Ę�J��pP�U�L������+���~$���dj$2>Ғ2�AFMQfSG">���4�����2�۳m"w�"��~<��x��)8�2��T"���ʆmz����Hjp������
����A��%y�_Nkg�y�+<�'�a<MnR	)&KJv��u��7x;R�e�Hp;q��Z�D�ZA�[�m��3�2+���NW�gbp�5f��s���D��F"�3^HV]ӗC��d�g"-�T�a�;�Nh�t�P$>���9�f��9��f��/��<~��וx�s���X`�//����\C�'b1eI�7j~;���f�艎���\6���į��
{��Nf�'�Ȉ~Ur���^���)a���Q�×���hr�f����̰��;709��
I��F$eXm�j��֡��X$]��k�n�LV;��_�˂�,z�f��ƱCu�@�jo�u}ߔ��A���������zb�!b�"�P̈��r�ۇ��i���^����2��w��2rICv'�w���4��3N�L#�-�8kM<��g�C}�����/�tC}�3��H6�Y);�\e��`��I�՝{��u��Y�M��wf��������d2���m��������y�+�����@a�8ަ�4r�^�IG�tv��u�Ǵ�J�N��Ʃs2�p�|wy����\�r��l��Ǯ�t�L��^/��(�T	���H�Y���P@,�=R���>��'JncQ���媒[I�Z�����`�״q�k쏒 Vbm)*d����� ̃�DRǐӆ���URT�t7��e�1�ƍ��hjd7�ƚIY�W9�qLD���$�+$!F�����Hy��$��9-�Ւ�I�b���zyk�m��wu����Z�/k���H�K���;#�G�a�K��L�~+}J�c�?̓1��B�3"G��#�O6��/��az�Ão��6{�`Gb0;IFe�TZ̞d��w�����#�g*��|��G�|�nnnu��B�ba�%�P�[�Ŏ�V�쩩U%�k.'������?�@[��]`V�dw�I��j.���d@�9�����}g�}K�9�ڴr���v5	~���+��1.����v���Z��*o����2��h��~B�� h�lg=��=҇��4��ԙ�� <�����Dr���#��IE�1�jmH ��_� ~a>��V���-�\�{1{��Z�˰�gٞ2kn�̇�D�4|���4\uU�r�T�.���<�MX��Ip�FޥF�-vp�3˰\�/�j�]�ܵ��2����� M��Le����]Deq3��W���K��qs^�:��Qw�����^ƭS��Y?��]Sh9��A/���~�����W��z�ݞ)�n����.�M���2��/��[��/��048z���G�g
�����jO�#%8��I�&k=U��u�'�+�)E�{��p�s���$���Ҵ��'Yr�	k�I�A!���l�[�����`#�b;کK'��G����k:[���peH��I��#T�*�g�q������x����g�uO��z�r�2s��!��Z�z�+�Ls+������;h�>�?��4�J��%�%<>�e`LQ�&L���,��j�N�}OjG��or�O�OM�W�����d�m2#��w�ۯ�׵���,�ω�i��j��GNc��g���w�;Ma9,(wwLbG�59�Ć�x�r��M���8(w���qT//�Nv��:y�L��?'ْB=u��|J��ۭKK/\�n��OS�"DqS�*�i��Y\�*�|�8�S��`7O�W!��cs�yk�y��m�t���a�s��o#�0
�b'F��	z���n��o��?���Vʌ���9阾bG]��X:��e�]5�{�>����[��ɲȒ��N�_���_����Iv���&�_V$Q��J܅|F3����ʜi2���g2�����=H?�c|UE�1ͮ�1�'���=���cY�g�wO�O��S�)�}m��.<�z���u��z�h$�O��'[��Ou�N=�}����+��E�y&��-�EC�dʛa2��eE�S�<���5L7W���e��+�#�_���_"��p�<ep
Gd�|D��!���K�c����8{��*��/�l�+L��\·�q��������@�3o��L��b�b	Cڄ�K^_�75�YBK+�g�Γ%!������)�mW�-����(�T6���+��0�r���(_��1��V�E��s�v�kR�
�|��|������ċ��'��m����z�鬾�f�/���%����k���}���f����$���`��zR��`����B���V�K��[�D��Q�)�i�Gy%i�j&A_��3� �e.����
<�lzm�W+5�kiރ
�*�}�����y������Z��0fe�:^Y�f�?d���S���r�k�+{��[��mj��ԗ����K�e6"�«�ˡ�ޔ�jfvܺ�q3��H:���G�O�g�g�͈׻NZ�
tf�C _d��%�����	�_�tt�@����yj!O4^E���N׶�v��r�ғݕe�
�f[V_�f՟�<�=���߬�y�R��b���%�D	}Hjۨo�CX�
V�2g�t)�P���Hߢ�79�mJ~7�;Z�.��^ݒ��-�����Ŝ|�5[��}
�	[5;u3"�-�MO7"�Z����"Qn��K�.���k���Kb�A�����\��6��6��5�m8%���l@璠j/��Y{ ��2+�3k˭���n�{;q�[�C�$������B.�!�X�%6��,�b�F>�[���4�)ɱS)-���l�ev��\cw�1���ƾ�[K�m(��j������)����bIC��qK~Uy~��<��a��Y�*[�E�'V�E��k�X��އ墆��fu�*]5(�eCWg��,�M�U7(Ցy�)Ub�^��:Q���Ck-�U�P�Mc�?��lTVXTVب�����Q�Ң򔨟ی�b��f�����Tj�;t��K8v�/�u�(�I%<%nauȍ�r[|��Ƨh�P�P���G�_�G>�t������kC~i~��,Z�ݥ��[��޴�l���Ի�R�T��re�e��|�4�{uZΧ�}�!�m7��@�ZOw�jޢ�a/�j�r57Sm�r5�ڣ\M:ѝVI�S�T��Wl��.�)i�V��r�IkW���*��u��FT�[�뱏'z���ؤ�������M|?;v��p.7k-n�!���DU�.���kґ��3�g/UZ�f�{�/�4l�4���4t�DF�>�ˉmbӌfĔv^� ��c/,�,�y������۱��V�]��~-�O͜�%�h"���t$��-W�,�����|a��Nv뵍j���D���wC6i���gPK
    +Q�H�Ү\�   �     org/bridj/GenericCallback.class  �       �       ;�o�>CNF���t���̔,}�ԼԢ�d�Ĝ����lvFF��ĲD��ļt}�����vfF4�z U���9����>���51����K��S�2sR��X@��������b� �L� PK
    +Q�H��@  �  $  org/bridj/HeadersReconstructor.class  �      @      �WYsU�n����$�$0.�%��a&�-l!�	&�(v&m�0�{f�Q\Pp�}�����ŗP#�˃�ZeYe��/��Gߌ�����@Re����;���s�sν7?���7 V�S�y�=�����݆�oة}F�J��v&��lB��~\���@xo�Q#�VP**��B�
�P��!�Mow������3�}ƣ
��i+Py�%S��Nv����!�x
���>+�`����v"Ϥ�x�CO.ڑH��
f	��L(�-�sfi�b&��&���e=A�b��2�(K�)����)o�����@c}�����a�}q�ٕ�V��6�^��D���[m[��)�m���җY���zjЉa���r�j�2
	�[����ˢ����9�%XZ�ŨG��+h`B�T�q2��s0�F4�c9V���#�Ǿ�������j�9�:��y܈�}�.�V@0�n�H�\���V<N,�Jn=�հ�^1�r4�8������TQ#!�[�\�>l�P��l"��H��V�ڲ(���U/��b��3�I�A.��~�����I�waw9v��z�TL��툖�4Lfh����4���KB��9fwK7fy�Cպ�_�=�i1N)�-ǃ2!s
��i�������A�d�cq=��S��z2i$�M�ͮ��G=Xt��p��"!N��IK�)�U�fԴ��L,�A&G�����
�)I)�'&dy<�4	X����&O�!�#RD�%�����vc8�㲝�p�z���İ+<�t�i#*gO�sZ����N��V`��;bw��	��qSi�>-d�O�}x*��/����=�&7��b��w���[lG!Ͱ;}$Z� ���q��ݒ�b�Sp�0�4\�pi�eh���q���FQS�\bS[vrPO�rٙC�h�p��Y�������
ﺔ��Z�L]UԊ���$�/_R�L�	���z��Un"�m$�t��xW�#�v,��t׺��3v�r�`["a��F
P����+������0��__�5��t���;�
q���>~G҄ ���Ԣq�!���u�?puױ��{:�X&)�ex��h��wX�|�ؘE5�!NcP����RF�%����_�#��b{$
�@EcH�bO	z�buS(�Eg	mvF��v���|9Ѳ�W�ސ���|u�jʂTeq��`8�`0�[~��q���Q�Io���Fql�]��1�cݐ�V
֓�ڙ�k_�[WIr�8����ᄧx}�K��y��z��Ps�y�y�'�m`R<˫�rIY �N������,�zyP?�g��[�,�ct��<oXxY"+0�Kx��3�Y~e��D�^����K<��?��
��, .��T���K��E}�/�h�)��W���Zn� ǯ������bU��x�%�Y2�.#�B�M�Ӎ���<�+��E�L]�\�b�f8�:�W��U��jƽ�|�%O�p���F2�1�O�w��^�f6�V|�V|���;��N�ɋ�_�������vt2����K����
����-��~��A?r��f�����ȇO�]H6fG��3�,��f�^x�W���PK
    +Q�H���D$  �    org/bridj/Init.c  �      $      �W[o�6~�~�"��hV��q���u�ځ�6@`$�fJS�D;M�����[I� �x.��΅��r���ڽ��w"��8�{s��n��L_��R$C��r�s�����Na�C�B����j6�~=_,�>�����q��c/�W�mL�;o板��ϼk�E��r*L����K��Bw>�I��������D ��.Z�+�r��5k�c�m��L/�ֈ��0B���A��
����8o��Х���B�7��1�"4���d~�,�>����%'�!��b"v1/0>�K��f���4�/�h��6�����ٍ�h�<�a={:���?�3(��������6b��]�����0%�T�����B�5�j�)��^rKg�cg�O�-�Ɠ����g���x�Հ����;�')p|���#��x'��Y=t�Υn�y���M(R--�"-r�?��3� ԕl�""ő���l��v�@,	�ɛ�S��$Uv���w�"�$r�ڵ�ڠ��G≚�C�x"bF�Y]R��QW��F;.LP'5e%��#���KdJ�:?��Q�L�`����=W�R	]qi%_ے�5S��B�!w�3{'(�!a7pO���(���G�( ��8�w�ħ!������;�J� 襒��P��Li:�(�0����W�t
r\ch��ө���JA�b�	�1~PM����"����:�_�r�,5�tn������|�l"�c�j�3I�#�B�&��Fl�:�'PA:
���M���YAA�!S�>�D��~;=U����Lͣ�N�.SK�I�����ٚݲ�b�S�L-tQ�`�V��hw�0���;�}�R���̲�Z��Ȕ�)���Z�z��棞t��N�غKTM�zgX>����d50Č�b֥���RA��}�r��b�YNR?x�^�*U��������O����.��q���x��/.P.���0�D� Y��R�1T�,5��8C�pi�Uj{�����L{!��Z�09�,G����)�瘑�q�(����A�Z̳�F���r����4�r��x��nS�J=���F��-�<��� �"��yi�ɩ���>�dEhX��Q�;J�=���p _pWUR��X(!}̵��0�(��l#Sp��s���b������L�I�-�U�6+�rF��<>���goj_Ֆ�5�p�a�жS�i��搑���'�9Vw���Q%&�a�2^�[$,'k�0�*���n��GۆpLHv��� �m������-��l�`��槶'�PK
    +Q�H;��   �     org/bridj/IntValuedEnum.class  �       �       ;�o�>CnF���t���̔,}ϼ��Ĝ��׼�\vFF7W+��ĲD��ļt}��M�������RVjr��� �)Ռ���XD�iag`cdBq�H7#gpfz^bIiQ*#Wp~iQr�[fN*P9+#;01p�If.0� PK
    +Q�HM!���      org/bridj/JNI$1.class        �      mRMo�@}ۤqb\ڦh�(�@�azN�K��)Q�r_'[w#cW������?��x뤠69��xv�{3�����/ �x)�����z<�g��CB`c"?K/�q�}&j�[(	��/�%:�U��H�L�V�$xe�k�X-T���]�2���]��P��/�tظ%��pca��WMT�t��c���:����2���Bgd�oL���\��.�nY��{�����>�m���7&8W����Jn�H?�#5<�d^$>jS|k�"9N�1����HFC�jD�1T�u�Φ���3��e_.�Jk�2������fZ0�كd���[]�GQ��8|��d,��ƱJO"�e*�k�p�\5��_{�<zA�������u�֙%qw��T�L���{�2�>���|Ã�5�R�o��s�����/�q��SF��.���0�~уK�VYhӗ�,�皆���\���PK
    +Q�H�&F@�  |    org/bridj/JNI.class  |      �      �X{W=��U��eKNq�����$�`cЮ�����P���ݷ�س3bf�F��j
����M���{��7��������|����w�y��{���=��{�p�ca�l�W�vf��R���0z�>gϻ��9c匨F첐%�j�X�^�0�v �v$jG,�$��&���َ��x����Cd0`a,�g0D�Z$�Gω�Yؕ;�6��DF-�E[NHi�y� ��":�S;JzYZ;aa(�U_Wea*W:��],�r}���T;ؑ����yD�B�Y}k��xlky�Q�]:�x��vN���WE�f:W�m�J��/W*�H�-��_�BSŶ�Þ8��Wl���wUk��Gjt��1G�Dzi���U�6/����0����"+/rt[#��B��������;�	�(\=�a�ӕ���{��(}����ʙ�v{���P�G��H����s&��s��D��I�C��M�b;4[
���_���Q/LR��� �w���!���drōu�3�b�攊�3�4���H���؝Ӕ=�rږAH9�� �0	ds��bQ�o�9��D j�{8�'�'���&e���f����}���!�ʲ2�K]=mˆm�ny�D��"%�'�ް��� �]�cO���3�I,�)�W���[�*�8��a@�%E�P&W�q�eIiӒJ}$솤e-�dg_�
Þ�ٮ,I0|P�i�:�ɞ`H���Ck�7=�=$E��ҕT"oz"�H!�!
[v��]H�!�X%�>`�P{者��+y��9`�,ĚVa��Myg��M�`�i��!أ��M˱bM[��ÒiZ�"!��M�|I%�L�& )�R�i5�jڴ{�+K�i9P=�f��ё�Z�Y�Kӂ�3�G+�H�0�#I%q�CLjBF�&EYԢL�v&�4��?Н)�v�J���}��K����9���fyZ�!��IZ�ur�q'��.�c1jR�2�A)Ϻ��`�v�2MM�0�B���;���W��S������������_���z��e���rBD[~M�E��i@>.�Q�vS[/��L']z[��؂YX�<���'[�W�B+*�;�
[h�C�)t�	���y'�p�:��vΗ�($���$�>Ŕ��Jܡ�H"e,�ј����6M�M9�M�A��=� �_]i���ԋ/\gӓ^5��R3�������WC�KC4�ۺ{� �!O�?'�(,_��ٴ%I���uڵ��lil������D>�V]�"4~];��A#��QP��ׄa�A�(��2
~M�Yا^�Ǧ��U[}n�,;�Xi6*4~k�`祎n�TӋ�]B���'��#�t�@�t��f@��������1��~3��%G�.zͽ$D(B\I�}�_�a�w=��gZ͓����{�K��9���ٿ�w��\g`S���
�w���L��>��d1�Ye�Re/3����
T�J<Dه␊H�:�^%y@�)�,�z*T�ud�"q�7_�#/��ww7Bo��&�;�(�?)�u&�c�1�X<N���	�^�lO����x�Ó�)X`�<
�����湁��T6O��S��d'd72�I<�AN�� �x���ynb�<��s3�g�,<�A����\�RA�AjRg�l�y��<���2���x�d�c� !�Dh2�9���<;���A^�3�K�Ry^� �`���*6�-l�[�j��a���u�z��Aވ���� w�y���y3��-l���m�v��Aމw1Ȼ�y/�� ���l��y>�������|�`�O�S�i|�A>��1�ݸ�>�/(��%e�L�߰n�\T�+��k�}�f�U3.|��l��o�׍���ߤE�o��U�,���*�=����`�?4��H���Tٟ������_�W�������m{�:��w���&�o[Д���>�r�m�7}��:�VY������+�?PK
    +Q�H����q  �    org/bridj/LastError.class  �      q      mUmSU~nB����-Ѐ5�$Ph}�Bi-m5@����n�%,��l�g�����������Jpd��O��G9>gw!��������<��?���'�K�R8U���9�,��f��sӶ�vJ�́`Vw�m�:�#����Ж/��vô

����-�,[
��荖t�8:�ئUg ��f�6K���+Ac���©���u��H
���
=��lC/d�y�� #�%�)�O��؄i�ΤB(�ɤ	1yxjQC��h��nG ="��,)p��
�[�Q��镵)��`2E�N��X�Q4��
�m�T5�VIF2��Q���G����pNv�L¸W�K�&�s�u#VX����"
�(\4['w7�x:�:ʆ�vD%�Qf���\�R�5�(����^4�zD��d���W�RAxx�%ɥ�rcx�0�F0���lƤpo�����x�t�[[�t�V�<r�&�)ܐ�7N$���.!]�����=��d�\�3b��"Ȳ�N���0+��0����lC+��V=�����yV�eO�q�D�[s���jX�'Q,b�A+���u�ֺU��ز�X�;�\\~!�9%��Kеj�Jk�����7���.��s%���(��	&G��;�▕>>U�*�n9�2	�y�h�N����Ҙ���n��sA,kZ�lu3g��Mt�\���-�dph�]pt�d|����������g�uym��|��܉�ԃ��|ҵ!�)q��;y���j��]���w�jorMxr��ߍ��Pu$X�GA9���0ØS���ǹF=��N�����r�p�v��ԣi���r3���\_E������C#�����_̈�a~����#��m���|��|�H������|���
y���;���3�_�����CG�r���������s�'����>mr�����`��
�o�]��
ȿ�toe�1�����Į<Ax���5܊��Eb�0�ᾆv{��!&-����QW�%o��<�n~�[w�R�,԰¢�_���7l�OI���i�d㏠�F�pW=�G`9޷���p�K������^���]���rS���+��!rF��\�@�)�	��6k��p:��H��_��	��\�.��PK
    +Q�H��3  �     org/bridj/MethodCallInfo$1.class  �      3      �V�nE���;��9@�PJ n� �I���P�8vq��ƥ	�n쩽a�vׁr�D �} $*qmUUU��WH�!�@�׈v�ݸjDe{��ؙٙ����; �Q'��N5����Բ�jv%��fκh'�# B|K��S�nUS��[��E�Nl͝�I��~�"�"����3vEڶ\O�<7Y�ͺ(^�t��M� F�ل�a�nY)N��g�V��]2�]o˨Zs"�#t����d�s�+ז��$$��$$mJh���[����seӰ��}b��K.�]��kYC�����N	]���%LLLn�`�f5c$�(��0��(��,!&J�Q�G���s�r��	۩�n���iCR��?	��<�Høʟ����V�a���="��?��)��/E�ῢ�i߯�N�������E��i�F`F^�Y�֛o(�M9��K^3}N�ozłm�B���Ud^6:���N�_P~Z�<ݬ�W�ӐQ~�Яf��G���ɨ?��蒊�e�hl?]Q�U9�5۰<�˻*�a@���RXT���ɘ�����s���O`�>z܉��z��a@m��x�fuד��0��>��(w�e�&]k�[�M��.�<�堡��ߣX3\en)�S>j�¡��'e�Б�+�s o�]J�c�=��B���X�oo
���
v�)���3Vٴ]ê�o��e	'm�+��(O��_�m�\�qH"x�x
O3�@�ڙ��n�Н�c7p����pG;V�Gǒ/'Yv��e�]�L����8��P�`ߓ}R�=�R��?%u4ԧ���zQ�P��Z�Y�{C�,��P�I����P����y�|}�k��u�ݼ�rs�X^d�J�eW(M�j�?��G�YD�?c8��q�	���"ck(0qe�
v�2z�
_3^�7��x��;�k�7o�.~a����;�}����o����@�HP�i�q�Fi����Y�9:Cg��D��IP������<��6,��l&`��V	�����k��{��{�d����%6������}ƿ�t������N^{�i�4� �L�T�n~�=��|����PK
    +Q�H=	�A!  �I    org/bridj/MethodCallInfo.class  �I      A!      �{	|T���9w�̒�d�d�e���$EE�B E�$�̄�I0ںԥu����
HBE����u�Z��[�V����e�dX��>�?���w�=�{�Y�{<��6ў�|�!����p�	#%Ś��ȔhK�I��=!�	F���xB�)�$Sy��2�i��Q���IL���ӂ�pG�!M$��d�rN0����r��ɷفN�0�S��vJF�#1�#M�c��Y���e�0{��J���@������hX9�ܧ���xg�ĆD2�."(c�om��1��p�*�Z.�+�ڌX	F�#��������t�2�1�i� �G&��i�L7��M�-�T��퀏�N$ǀ�~��S�S3Ê�CM�`<]�	&@�tjZ34����na�l�A�C�J�d{<���<ܵ���D
���h�Z�6A�2��C-��4��1��[A�,c䬤�-#������m�ŗ�͡��p4)�,ln�^f��P$2��`�5�Q�E@����'4[�	KÉ�C�P<ܔ��1Q8�1"1�X�x�=Ki�J���`c$4��%��7k"�����V|||!$�
'f%!�&M�aF�=!����D�aB�dbn8�h���la�P�9!)�$�cKS���x<H�|�_L44��Jlg(.�$&��-��`l8N�cڱj�U=�i�-�o	Ӣ�t��A1�z�Oݜ��k��;B���X+�nU�v��Tc�J�s�t��P�hϠ��xA3=4�fe�M��#!��b�,X���/��-�KGyh̓�1׬��P�ɘMy֌�u���cd�c�W�x�k8�'�|Ū������/;�;�,c�R���񩦓�vͤ�s�'AN�&&r�,�Gow�ѓѓ�P��
gj�cΐ͑��h?�=�^ȷY^`�m�P[(�|�)��Qe�z(�b�OUn��آz�JX4ƴڡLi��n���K`�P�m�lV�����N��It
�^	YH]�fWR}t2��S��i051k��rqa>�<)j�o�%�������b�֌3�7�gB3L J�h�Pl�6���Ud���`��\h�漙��׺���[-�P��������{�D��.�	/���F�f]n�HӺA�k���t�EWS�̳.4��h']��"�� ��C����W(ߤI�g,�"�n���]�$��Xt�A��/;�c��������ek[�=p�ግ�%�oL���7��[�SY�}��C��*��ټ�Qo���N�[)O�.��IJO�P?W���VGX�M=����k�%L��NZ��j�=M��Pn�z���A��4B#�hjk�0c�	Y.�`��4M���ƙ���ɸm�X�	M#Rَ��h?3n�	ri�l�F��%G�����YQ0��-�=%��v��VVUo]�=C�
��Y��U�t�/Ћ����~����C�q�q�
�*$^��3��Z�pPؖ5�AZo"S�L�B�r����B��_�L���氪�/��/��7#�I'5��d���EQ}ԗ3�ǃ���O�R��b3�ڗ ��^,��>����slyv���D�NLjmKvZ�5�RH_�7h��[h}z9���I���j�E��p�@G	޿,�`�~�����=���L��H���j��i��ִ����x�~�7>�-�DZ55eg��"�4%�%]$�J���8Hm�^{�b���l�f��p��.��������NhG�^;��D�y���e<H��M�"��&�6���v�1��jl_h����<`�A���H��@�x'Ibr��[��/�bѮ4L�2��Ƣ�����ߔ�.���ݱ�ɘ�aq5z�t�뗸���k�ΒG����<p����S���l��{��ͣ`9i�����tv,�
��j�6���l�r��;�<���;��L�Q�_]5e����(�m#�y��<�cG(�9'o�%B�3jy ��[��P����1�SmFD�&�L,��n[<Y17��6iđ��>̢Q:���-�˴�[��ia�AƢgY4޴Pl�e�Q$�l��[�<W����h3�|��!��Qr&�dm���I �1@��%�x�`��9f9>P��I���b��8�G�7ba %��q~s����-�߲���a��u'@�nm�hg����kK�/���`����Lh6}t+���(6�Ǣ+)��ǟ��â��	O�����gЖ�lJ�;(k푲5:u4�e���g$He3,0sr0�i��Ŋ7�':<��A�Z�@��f�Ar*4@Oh����+g-	'�AE�$�R+f%]�?���	9N��C�b��Iq��RL��>��RѢ)[֢�E�� ��~X ��~�������X���4i����F�Ȥ�_.������K�r���7�D�Q/9��ݖ$g��}��5����9-�.!z�&czj����S��w�݂�+�1���Z؜n��_������q
�ċ)^m�؉�C��,R҄��p���:I��"�͑'��^^�9� �s�I�'f��z84���D��Y�g@$��E2+���"��Gu��(_Tk��S�VC��v;C}�[j|EV� "�.�p�P�2[�d�9�ɬ�@�vF��SY��婱�B'?��6�Vr�JB��g�g=�Ay�4{ތI��|�_����f±�[C���ɯ0�fݟXk�4�c�H��1�oO����G@ޟr��~q���ům&���~���h�:}��fM���BdDdy�!cn��	 *ȿ(�����0:��W	��`|a�l�����������a|�l����?Β؜X���w�������!�H_$�"�i�)H�JR�����C ����PW��Y'ӳ���4?��'!~`c��`�����dȩح� xB�lƫ<=^�g�*6
F���V.A)
� �c�
�����NU�V�z�@B���ʡ�R�®�ل��AY�߰��$	��V�	1kn�!�g.�m�@�����\n�����1�$~b�]�H��V~M+d 6ήgX�)��#��Ԩ�q�6���*Ek�SE��PjJ]�lXPF
�ng��iPPx�	�i����y���8p���V�xh�y6�C��R�/��M�Q���`�����Q�C{�_�w��_������J�:H��f���7�a�B�Y�Ĭp���I��V���4N��hxq{(��@���W
�4j�ǳ]�!j��NR�"�	�������%���p�4�B���Hp!rK�0+<"�=m�{\����7K{澾�$��M��TH��I�T/Mo�w��G+���{�Q�h���P�o��&��c&u�:��Y���7�f|©�p����_����"�L�l��dM�٣V:�H���d�o6QeI]$����R���ɠ�����mR�T�Q�¢(1�@��Ģ�'%���o�'��;�t��oi�6��YF�T�fȼ4�nSsxm�Q����?��r��S�=4D!�(e*��Yڍ�v N'��b�ڛ�F:�+�9�i1��d��d��-�׍���~�~��r�o"1�4����h
#VI�s9�N1(�z�Ͳ�码��da+�n��<���\�x~8�tJ{.��aM:m:�R�K��:"gm��3K]��R��ԥ.�r�nR� ��Bە&��^�Y.Յ�D����.un\��˴בQSS4��.��T-iB$\�������Mz,�bq�7��AP��R��B�-W2��!g���;���;�3ƥ�/@�EI������}�`� ^�+���Kݏ�!�(��v�k�����T�L�2�II�x�,v�ӫ������f��=�@O	�a&
�����c�9
5AA$](�ǥʙ�� ���Z<"�)9
Q�m�zB��&06 a�	K3Υ�,_f4I�@�y��+3I&��]u��G(������|]�?H�����NJٜ+0���)�����U*.e�5��Q�/�5�QU-���Ĝ�[��L�.�п�b-{��-���(��%vŗ��&�s�����}�ӏ7�(9��@1_�H��IΫ��G����f�ߐ�|���ɢ�FL_c��6E�b#��(lN��7;�P�oM���ߝ�ey�f�5S�lN0W�?S��д���P܆��;��y��×S�ݖ����u+�59N������p������}W𿟹3m�s��g��o��z�Y��xShrX�Ś�n�ߌ�.�P��kg����R�+K=W�*O�gw���j
�{��{������ē��=m�(���}���;�N���������]ɧ4�y���}g�������}�}o����"���1M����4f"rjj�ҡ�db�/�6`:��j"N�\V?���}󩀎&��)�[��l�!��]�C�(?o�;l�/�8V�ۑ1�PZ i�n���	m<�>�_O9���{�l�`d)5����.��������c�����C�T[��!
��W0R�+�0��'-�)�Y+�V̑��E��8��Şjb2������x��MI��pM/������N���U�;�z�4�f��@�� �M�zƀ�ơ[��o5��W��k{M�D�'7����S90�1F�<��v�n"��'v�<����.���t�ر�n즛��nZ�ǻF畭�������ek�v�&*ꥇ�ș�������˨\�=�K��uu�cY}���=�'q=��y\/�z�[aEDX�����;}΍T�9�ѻL=�Am}�K_Ի|�u���$����*�~�����y�����R��Gm#�2P�W��#��}BK[��X��� ~f���������a��<�'�꣜�V�@s�����Oi��v\)u�v"��A;�7�o_�hŁ��\혵�d	��I��#N�\�BwN���z��Ō�ѫt>�Gb���;��~������R.�+xg��+�*�����#2�3��s��~5.���MT��������?���*������+�p� ��O��z����`��s�<�Ak���J7�t�+�b���a�\_��W���C���g�jޡ����c9��û�p�&r��n˩���z˹J��+p�����#����*�ռW9��+���1������fZ�+�(UYɭ4 P_���>' =|@}�j>��vH�3�}e=<)5{+Jr��4�g��}E��^��UXt��hs/6���(������D%�&:T&*ɘH�Jj�R��wH7O�,���i��1#�+֍�bڏ-#W�;���Zc����l��35���GwQq/'PW+
{��V{����-F���p��2�u�ٷi��Hu���Xzm��ŦkF��隙���Ԥ��i_N�Č�Lϑ�!O� �CG����^>���S�Jy1���=����v]"��k�|*�&��Ӂ�t��	�nI��ӭ�	��������-�.�+>ɭ[�<�T��gb�B�S]�g���Fk�9|ZE��:��V1������iI�ǲWQI��c}�4��:*����o�Cᇎ��)I���FK�v�Z>����N����
z��Mt/=C�ы���J�Ç��ZZ�{Q/O��<���6`�G �Gy	�����|-m�{ѿ�����8=�O�S�:��ߡ��zV��9UJ/���E5�^R��O������Co���Mu<��Z�m�w�b�Hu���T�T�E���s� }�^�/՗������(�o��?!�s�2�	�$ֱ;*p��T�7�L��P-�������}v�tg�&�[���{���j����w�>̑��KҀ�p�c_�1iDg�X��ˀ���v�c\�������0f�TΗ3���+���,gקٙy❩,�N��ev�8��/���!K�}e�=�!���ʅ4��i6��<��1\FAF��
���tCr�n�8i'�{�)oB�_�׃��9f"RMF`�15��fE��#��|�js�SLށ��#�ܙ*�O#y��m|���\��7��9l�R�r��;� X��(h�}+�i��-(F�u�p�xwL����$�2Gz��^^;v(󪀽K���;1����	޷�BG�uQ �ǃY�!���:*�=hO�6�C43�:�쿐��{yCN�i[G���D��u�t:?B+�
��N
�rI����<_�F;�+��͐���q���y#ܭҭMp�H����?R^F]�����R��,�۵ȿ����0�_6� F��g_��@�fg9?��v��s�͏=��ջ+�˨��jI�rS]9�pU׭�o�]���R��:v�Τ#�������.*�at����4S����w��h�<���H�I������C�(�E�]��<ח꼟1ȹW�w����uȘ��g=�9|�j�j%���6� ����ϕfy�v",�2��d���̐�I Ji�rhH�@\��K �Rr;zT�jU��Ct��X��C_�v���%�S)��n'�U-�5���G�y��H��zԾ]�����Uc�=�ɔ:@�)OF2�u �@��m�C^�)��V����q�\��P@����J[��نH3�{�������B_�u|�j��,�j�0k��� �H
U�Z͎��^�xn`=�|�g�Jb��%+׫ΔΨS�R��Q�j�g�:�a��9j����d��T��R����G�K���Ju&"��Ρ����-TI:N�V�c�!����E�K�[��(�+�	i��%��^1�|��. �o���P�4D}�.й���Uu�������>�Yg�*G�,��Q����qL��͇�D>��x-B���`3��Eg�l:��R��j�(Z���z�O@>�"/@�z<}��(U��{�Q��P^���:>��p��(�1>���s'x!��o��%|w��|
_����׈����|:/G��|&�Ff�#�#��=�M|.�����dv�|�+�K��/U�|���j'�R��W�Z�R{�25��Q�Zu,_���F��u1ߢ�|�:�oC޸\-廰�w�+�N��W�?">����y��"��7�j줆W�s�<�ٯG���ھ�l����\�Z�.�Eq"i��#X��H\A\��:q]�k5�:)'z׻�>
�+��.\w�و?�������2��K�ri�H�
i����F�������?���j��F��r^+D����	!�L���m���Ҿ��"���[o��o��)�	ҾI�1�7��9^:3�㪵a{	�������S]zv�%��[`� �������V��)�Q�����٣����Xz�Ǧ���M��7x� V� ����f�G��yg������ҁ"�Q����,'֋�Z�cE��G�]t��k�<_�#����CL����H�>kCލ�Y�Q�E�"=��W����#%0��ES���>�0�P���<q��{ԓ����/�[����\���T���`׹>�&r�<�:���4�@
*�R���ћ��7���$�nՃL]�f���B�o���t��z��Z��GMi���*��>��V/ yTv��h�l�/ZRS��T��%ե��U�p@a��z�F��:����q2f��y�sĜ�.:��ϿG�{��H�"�u�&j�'�$~�~�Hs����i:����Yx���:~�n��.~�V�kԍj��*̷PY����T�|�����%��^��-���ʟ�����	J����A����;�?����p����{��x$��{�O��/�σ=N)�<�|>_�R��˔��R��B�IY���%�^^�J�[��:5�7�
~L�j?	����ߪ�{����jW�W��JP���h��h<�Q5*���b5B���Pg�=�F��0���Z�Q��}U��O=��W߫��� G����G���(W�C�!���R�O.5���Pۓ��2v� ���h^��G��MW��¾S��u�.�\|����p[ͥ|u�t��X��!�Z�������id�i�i�h�71y�j�&@^U��>:�Z}��.�K��cF&#�ikȈyŔ.)R���	`�D[��҅t�=K&��[g1jA�^Wi�9�k�������-�L�fe2c	@�Ro�d��Ro޳U�:���|��lˬ20���:��r�R���(שCe��J��̰Y������o�Τa�l��G]���[=�A���\�)]�u�_ ���TT�jKB�OQ�b5���\��6���Ȉ�M I��<�M�>ɁQ�7��;y��e��f���rG����v9��J��j�M-CV~-ժ�v-H����*
�z<_����R
SK)�p��C݂�H���ʹ)[ߔ;����p ��x뛲h�������6E��fn�J�d ����ڭ��-�%��LZk@[K�s(�/�.�^�}�ۼ��Ң��3���C���H���zF��2�.��S��B!�g���2����CG��^B|!Y�x�� �S.p���P���N��PK
    +Q�H�4g�    ,  org/bridj/NativeConstants$CallbackType.class        �      �TkOA=��nץ`-> ��JA�m��b*|�ڤ��tY��k�[��D�F�g���lC�ä�d�;��{�L����`E�Y�o���_��}h�=�p7h͔��4��������1�T��!/8�m6��A����J�R�
b��yQ�0�߶
��7ä��Xg9/�l�]3�=�!ۯJ�a+,�z�-E^�˭3�|���6w�Z���ˠ��^V�m���Or�m����i:1�D71�M�sɓL6�sW;�}��v75c�$�a;JٞJ#�m�Y���z��^vx�U�����')���$C��$9}�F��l�VF�P���鸇)�g��{6���L�K�fs5�F�L��pM5�Bס����!XP�ґ
�jX�vI�`�v���A���H��ɝ�m��ɤa7]�}z���֦-6�-׵|i��Z[��q���kcB@Q�ƁnL�84.��*cH�:� �	MQ��A��N1���SZro���q�[�D�DVKG���)"�>�g�����.���+���o"J?@��O�`��]�}!����y ���B��A�S��H=��� w��c�KP�K�(��K�/B��F=���Q�w�h�,���Y0"��$+_�	�i�Y�N5E�B�V����H���PK
    +Q�H'!
�  ,  )  org/bridj/NativeConstants$ValueType.class  ,            ���RU��� ل�d�_�
�M@KiK)MJ�,6B���E��CX��b�A�x^�W�ngZG�N?;~w�+�
����9k&`�!���s��g�sȯ����
&�Fmv�a��n�y���t�mN���KOy����qd�Z�]�]�[�|������������H���(��5#�(��V�e��
Ξ��|��o4��^^(:v-�����^u���-/�#�����#z�i�k1��������Xܰۓ;3~�i�X��̺�n;�c�.o�7\�,�i6�H�|�2j:w��|�c��xɬ��92U^)�_��{xʃ�9��d���axg����(�Z�M{�g�I�E�S8�$�Qqb��=���H�m�v-�=e���h6so[��ͤ:2���3
�l�N����F��7m�]R0��7�e�Y\�י�u�}�Uj�jI�L��"���c���?�k*��Sg�KYR�`HHYQ�dHJ��BcФ|�"Ő��4CZ�'*����U���/EW1�0 �jd�RQ1�0$告a�a)_�a���b�aT
W1�0&e_�8ø�/�
�.g�h�|�U�ፒAW�?`�jXe�a�Fu�fn�����N�Q��?�6l�7DCys�"��M�d}�#�9D000P�
���?�@���C��8pܧ6��~��Q�����N6A�?1/q�&��)���#�f(>�l�����C�?�7��!8�dr��s����Y��a����W���Dz��r����y����,D��^į������_a��\��r�[�M!�=BV�"Bք��Bn��d�aEMn
��d�=a�jQa%a����ma�i��{�1a��}�Ņ=fh	aUa�ZR؞���	3�h)a����<�aQ�ty��n7�J��U��WT���FCw4�I��{����ھM�����<<&�=<!$<T	I{̓IHy���x޾%�tOA=�S�G����W��+�Ds�������;,�{\�X�3\�k����7�'��5;�;��{��J��UD���PK
    +Q�H,"�G  �    org/bridj/NativeConstants.class  �            uNMK�@�ׯ�m�U+^���xT��R��7�R7n7�I
�,O��?J|�""d��̛7ov?>���a��۹X5���H�R��IRa��:�X
O3��H���*���z���ҬC_h��q��$4�_�pP�::��{MB�%4.�Q��zt<u�b���	��A%��Qi���x�!�Q
=V�@�I~�#e�8[��(��8���Qy��#��E������!.�c��9c��O^�~aR�fa(Dt����j�p�5���Y�6c��õ2���a�PK
    +Q�H���;X  t  &  org/bridj/NativeEntities$Builder.class  t      X      ��{O�PƟínt�&����d��B�L�DȌF���Y[ҵ$~,Q?���t��[FL�G��<�9��r����� �����k�v��=�3��:Ԫ��4Ү�B`�.�dٕ�qy�VWvh�_`���z�I`�"��!���E�j�����sX�$Q�ݲ���Z��i��*<�t�������tF�MBDN�����xkM������dS+��_��m�Ц�t�%�_(VM�b,���鴤'A ?�u���$�Md�͠�&�D]1�K�U�D͛IԢ�@x��o���E��a�8;��	�.G��.ۇg��!�s)X��Q|c�
ø�"�Ҥ�^��FV�߉L�z�e�c�$��r�����t�@{2��*��ϸ��ҭ�@˚��o�Ҟڋ>�T�r�~�jG�s��TPqe����1�o��ہ�z�|��\�:߱i[Q����:�����9&J?0��S_1���TΥr!�K�����ʚ,V���>YF�
{�f�:VZy�я#f�fV��ԇW)g*��8�Z�O��=v�O�vW�lė$�Y�J�����wt�]�=ߓ(���J\�萨�6��Q3"�\B�PK
    +Q�H`j�G  �  %  org/bridj/NativeEntities$CBInfo.class  �      G      �P�N1=e�� b�X81>6M�\hH\v�B��If��b��𣌷Սc����{Ϲ���|{p�:�^�� ����穜�k��T��s���c(O��{!Wc�6��aj�b���"��_�6��oW"�F�``]�l"�5���B*�^2�]�5`�����e�%dQvPD��*��h�F�t"���?�9��N4�V�^4��ǒ���������S ⟛�]4���F���q'�I"4�u�~1C�f�^4!=��]!�Q� �Թ�W���������a�
(�l��1ô��m�crLxB�S�?#��q�a�N���F�/PK
    +Q�H����  �    org/bridj/NativeEntities.class  �      �      �WYwE�j2��I!@Yu&A#��Q2I�n=3����{z�����( Y\	��������x��
�ԯ�g�$,�]}��[����W5���ݏ V�{�y��ה���@S��C�Z�1C�(�ڐ֔�̾��=�(���׼N*	���iY[�H�t[�4%�!p�y�cmf���Z`�7��͚Iǰ̌�̸V�1�M��f�v��%^�;��2������E�kn��C��d��z��R\k�����,bZ:�В����@�ӒƔ�^ƅtۍq���i=% �p-�i8���&s07� �f��^�e���y!�G�
ӫ�3��"���
������op��ϻ=�J����etvQ���NWs�)=���҇t���u̮�5�
L��UA#w3���:�����=f�Ӻ[�f��,G����4��2���P��y�����F����I�n�[��~-ӥ?��ݢ�6����ঃ�+�S�]�bz��R��_3Si�Ft�X��j��y��!�*֢]
�b:J����P�A��2e��<:�3e�}�Ne��CV�n�C��zF"5;]8ŊHR��S�G`�T�T��;�yZ�L���>bU��T6�Y�%�.�(��2�7U	X�^���̅��$px���R�5z���ג7G&���-O�Q�:�d��߶��m��t2������-/ndd�HUC�4�?���Ń[;���1��9Y�h�đc��mm�@$�u2`�S�T����A�[��s߬�_�`�d���B��mq��Q��AV�vH����`���529�)�*�xJv�Ӓb�L>KV�����s^(�K:r�^$v
V~h�쩾"��U}M`�JX����*�$	��e�ػ�`/(o��Gic�f�nÎ&2æ��p���p�e����*�˦�u��|my�<�d�d��a�\�=R��+x�0�ӝ.m�>�w�U��˱<��#R�G��mKFl�"����,9�#|"]B��TV��ң��B8&Sp�IZS�����A�H���դ���|���tjr�-�t�@�O���S�`����X%�t�\�m���Y�qcV����E�ۤن{�|�K�a�]�m	��K��j�Y~�Idu��A9_��������H�0M�v=�,!Z��WU���g8
`�3'|�N��U�];O���$�m��o��DG��5��e��s�������0\.uݎ�a�p%��}��t
�@�����q��b���o��p�ц3X���9�,o̡E�H8�S�g��/?�5��;������~�R����_��FO��o�~)�Q���PR��m�V(k/�veCEY�(;V�1Oeyme��b,���2XI���ۃ�����ó������,sx��U������b�o�[��l���YY��<��7Y̷8��,�I�@T� sћ�c��"*��8�P�/��rx<��e��Eg�=�g*���;}6�6;�6/�l^�ل6/�m^�����,-���ۼY���U�S�=��8�����Á�1�k��çè�1Ύ�4������-������p'd��@>�rt_H}���W�e��kB��
�w�>�H濍}��>6�~�~�@8H�0�	�	�#�Q��s��'�)F�c���yȡ�� �n�d���NC	� Xq�%����*�i����|�q��W�j5��PK
    +Q�H��/�  �    org/bridj/NativeError.class  �      �      mQ]/Q=�ok�V���?���sE����x��7�6kWn��g��~���6݇�{Ϝs������;�mTE_;��Vv�v*u'��uDȶĝ���sj=0N���	�Ԏ�T��^V�Grh�9������jJ����	��nG�����?���K'�~��_l��\[r�#���m&o �QBl�>�"�/no�g�����,�&J�&�?���9iL�^�3���,!�]�P�����y,���<aۚ'B��ށoG��{!�MW�����P�<��4��!ƙ��W�H�2��/ ���� a�o�|�qNU֟1���8�uQ�T)�b��g#�m �*2F�絇xT)�!w��B~�	��/��􄥇os�L�2V8[�}�lq,G��PK
    +Q�H�@�;�   o  ,  org/bridj/NativeLibrary$SymbolAccepter.class  o      �       ��AO�@���"�^�yR�l<s"�Fܸm˄l��f[I�k��(�В&��wx����}~xFH�+�*J�Yfћ�̆c�8�7��:)�8M��b�@� �Y���Y�qZ)�����n�.y-�5BM��p]�'\�oU���O�W�08�,��%��>>)��aA�͋��L�O�݋�eɥ���ƾ�-�p)�CP�3\�E)tѓ��ǅ��PK
    +Q�H�'|g  H/    org/bridj/NativeLibrary.class  H/            �Z	|T��?�e2of򀐐� �aO&	A�4���&$	�Ơ8I^��d&�L P�K�Vi��.���v1�ne��*Z[hm�j�j[�u�Z�v��|��ޛ-L ?~�̼w��{��9�����Dt���ir(���5�o�U����w�u�ְ/�W%f�������;+6���ۢ*e1����c�ݸ��5�jkӻ�zX%;���1�9���z����j�Q[<Tr2�}jR�r��&=S�i���]�zx�ޡ�x&g���Ӭ\�\�+����*Md��0�:}����ĵLjĐ.�d��E;�Ϻ���a,]�4���m��Z��o�C���AC�k�Qԯ��Ժ�&�ρ��koo	5���k�ɫ'�T���1�>}dy�Du!�SwFZvX9��cK#L�c���!���E"zX4Y��Zz;4z1Ի��G/�3��Cmm�6,�k�fc���2e�l�h6��F%LS�R�J�.*��΢iNRh�F�i�<-�h�ӹ�O���T����� �|���h)���۩GW�[>��$��-��B�B#7M��.�%��E;B�.����O�H�i�'��5gH��V�����A��~x�{LrS`�H����C�p�h��p�S8�ĎP ڳ�ak��ƶ��;
\ɤ�L������Pi#���ͺ�]P�"m}��O�'���a<Ǩ�h5�h+}��0NZ��ѡ����x`~q]:#ˬ�]�B��1G\���w0)^�\t�����A�qRq��j�N�pH�}��z������=������.�ȪS��숆�I�B"�e��4}��[7m�x�㣸��푒KJKZ.-�Ļ��A����;�ފM�(0��m��n��Oq���B�ݴ�E=�]�h[�d���<Vu��=z�M����\N������ZD*}N���Nq�F�е.���c���tKd�d4��t�P��&���*}���í����M4�I7��,`(o�/��=u�=#<��&ϼ2OG�'���FB����	��8�'�[ ���2���1P���nwa�;p���!���R�Yk}�K���I��������Z=�5:hr��o�ݨ�ޘ��8��ll����/�6����p���n� �� _�����6YVi��L����[�:n�K(�;nl�׉�-�L,��`ٕi>C^�?�;G �H_��"u�7& ���v���F4zJ<y)=e�#U�Ki�9�,(���A�F��P5}C�zjp!�C��ܡ��F�o1�@�L���j5z���o�w�,)�V��{���B��^?4P��O4S��7� �t�)��'L_�_a�}RX�AqE=������
����^2P����a�Z��/%:��~�1��x���_K}�ټ����	��JJx�~''{�J�������L�zWwHF��F�>�"�*�.���q�z�&�儍��I�R鏰dX�
��G%��?�;9�6��v�O��Ϧ����"��K]#��SI6L� �{j�)�����x�E�VyT���#���(��'�P���6_���5H�0L��]t��NJZ�<t6j-�N�.�Z�U��U�d�8kHc'�r��hV\X? ��Z�x�F/ʓ¹p6�<�Ak��Ȃ�C��8�ē �Bz)���3,���n�	3է9'��TTI��kz�����ԻLO-�Bѵ�Ւ���Q %y!^+�.�������L�&.��|FZ�h�*9���g�����8Ӿ�"��cٙ���4�yAf
���\��yiż�\�6�Q�<�,*�2-:�g&@y��|d�ݾ@����s��� u����/��>cT��^,+�xEn�>��C�Q�<�/NAqIK���������Cr=,v��a�4��e�`3	��*_���b?1��ja��^���S��B#v��.�x-���5�ar�k��x߀D�X����Dd��5�8���N�"i�*_�u�"zoT�F�6�7�t!(�����~l�&��H���CUZ�e���SŦ�g�v4.g#?"�����mz8�l�h��D�6� �vH�Z͗n�R<q����p�hg�]���qJ��RT�q'�E4*�2Q��Au�1����L8enm�2���W@RĻ�ޙ�׈X�g�2��˘�*	��g�غk'��.�	K��*��d0 A�D�%�:�%�ܞ����o܆���X6���F���C4�h�?��*��3�Ec^�������3�����[~�o�!�oB���g,]ڝAJ�A��A�/G�����j4S�]��1�JV:B�.�<�����oO������T��ş7�0�o��B���ߴ�yG]M����k�|7�����_�t]�=��P���/�A�����m���хm��{�[�������T�y�X �T�x�Y6}U���yH��i�œ�kk3.�G�1�g�5j?���Ǔ\W��H���*J.���!w8i���.�@a��8�G�O�mK?%�)����Qt��̇�h�������K�r�+ԓ��f�7����\��:�[�n���Hh�=���2ԭgX�~��+���n�m���.߂����8|3� �x����"�F��#�X�_n
G�K��냟�K�?��Y��ڏ6�n��/�Q_8
<�vj�+���-�2 .��1��7t�����$RǤ��HSh\��w�kp�=�p�X�q��o w�����e\�0z-�Q���d�"h5�5�R���p1���G�ᔀP��q�R������k���+6�J*� �b�����Yf-����W�p0���hh��k]����x�	lY求Ho�Z���¼z2~)+>m�%~4Y�)Y�n��Cb�CW�ϕ+�-����k�3U�1� &����H��,����)�z.���5I	Q����������w����zȡ�˅�x�hJ��P�7���v۪�?6)S��+ Ǹ�W���r��L����Ngfƽ֭Z�(e�"��QΒ��F7�	H��0�w,oX��L� ��\$�v=���L�h��@-�0e��hu6�w1j�V�.��Bm��6_��=[�Cn'�A��G��F\�������^)^
�7��ߤj��q���]���	���-ZM0�����A
و�A+�<���wH�M�)�̕_`���h��tG���I�"|zR�g�N�ϓ�w6�!E)��A����;H^��5R����s��#��[h;B����Q����Z�\:H�1������C��R�O�!�2ZG������$�P�'9�M���8�G���&P3h.ơZ �vZB�R%�P*@a�y�FǁD�
����'h�#	4s����n���o�%sbq��iw@�zj0+3(��9#��Jk�+�Q��+r=O�}Z��������#{��7��V�G1!���G��P���҆���9�u��*m�1��\�}���6wv�.�u�(���-�-FWT��"C��Ru�n{���t�1�xU���D��0}��J�� }:�fp��/��p;��s� �!����tA��ܮ���{���$$��U��9G�iZ]��� �� -���P����נ�g�e��5z��&z�ޥM��6U�M9t-���=����a(v}��X6L}=J����(B���Ct�T�Gm�8=���t�bp'��!��=PC3��b���Et9(���nZ��)LP���	w�o/v܋�}��]GWBҫ��v�\��,������܏�݄�}���N: �#�5+��iU|78WJ��a*`�K��_�#W��.��!�f�+���1u|>^XY�͘���f����-*��%�vt�&(�q	4$/ZE?>d�DZAO!�mTM�oĔmh�\qc�kn�gAw+�s�;�w"J�����@K�b���`|1�cDE��s�Q!����F�漟�Ϗ���0-J�������B?���bK�����"\]�<�ŏ%$�$�%X��K�Cqm�������H,���F�"F����d���u
:>A+�Q�a��<�{
��y��_���`�:��}�=�Heߟ��(�o}�C)Ǯ��a�DH�ह�
8�8��~5B����p\?}�B��}A�<x���e�y�'
tz��⬤��	`w�M�=$_0� o���X�!�+����ۏ�T�*fM�8���c�(��G�1�X:��3�&E�j�#�'�hc(B(�^$٦ �La�!ކ�xL�঳y*h�R���?��O /!A�T��r8I�z��i�>��N8MI>{J���C\�{깡4���\�S������n�0�fl�I���"�r�3�h��bl��o���lx�;�l�W0�a�Q���i���a�Ë;{�71U���a���<53�j�T�n5ƗJ8Ng{�t�CI�yo|ޘ9̾>r�s[?��YO�=Fv�c���g ��>���;+����rQ%���H�Dr�B�#�Y�_f�,�4�ষ���8���9�����r�y2���2���1���t��^�G�$nL.ὼƜ�S��|%L=&gQ��*���~�W���s� 1G���.l�H������5���^G���@y����H�o��xû����I�<|!���?����W�?X���gx���Y<�m<��<�qbTa|]k��|�lC|�ã��6��`��~���v�U�O���2ʹ��eJ�L���a�Wx -d��fh>`1�мbH���)��ۅ�<���~B��Q��!S'��	����~Z\w����y�ɐ*e�]�3G\�T8N��|o?M��a�_���RT�9�p�P��\c��Lag���`�,��l:��Z�t.��
?h)r�+�\��:Nn����>�쑗�!>4�-���f嫖�8�T���Xj[` #њ�mbN���^��2(��f1 Rn�,9n��"�bQ�Ȃ}�Ȇ�I�	U>�A�g���A��QC�49�˾b7Q��8!�bS��-�ʖP/��h
�o���ʙ��0�47�UQ��r5�z�� �'�ϻm�a@-�K*�W�L�/vێC�i�f���X*���,@�m@�c�C8�������_�^� �.�������2�T8��-���ZZn�^��j:���I��ՠ[K��B^�L�!���\��� ���R�Hky��E��7S7���P��R����|1dl�����%^�(���.��Lt��w���x�Ф�ׄ�k���=��!��]��p����O/�e-�.�.�}�~U^�}�$��hI�[��m�җ����ۭn�d�uպ���+�N�șB4'=���8>���T4vs�Y�4%V�_�Ͽ�'�7Q�,����ng�jZ��B��v��Wp��o�gs��Y��}������x�)���%�'���Z�Yc@hC��;��͖���T��#@E1���ۄ!�d@Q��| _q�x'�MVp�������'�T�L�*.x�������(��Pr���^U�)��%�HlQ<e�~j0V�8L��Y�A��s�EKߩ��ÛoE�#n�7�#wR>�����.��W ����x���&ދ��v�U���J�|݌t{�#�q��t�<�7��|�~���?�m����|�H����y��m|/��A~������fD�D%�J-`L"}I�2�4�L�3:%�����(�fo�2-��-�dv� ��~D��3b�L�y��km��cٕY�l @	F�M��$�Kxw"����Wȅ���ÔǏ��x(> M=N���>�h6�ȡ̉7��ǉyJL����q�M\!�v��x��-[Yd�Hy���N@�F� �|��;����PK
    +Q�HA�48�   )    org/bridj/NativeList.class  )      �       mOI
�@�v�����ԃ�W=z
*$��!L	����(q����������=�0W1�<$l˵<	O�"��`�%��Yʳ���DD�Y�RO��2e���!��j�ާ�B��;��5�����2�BF���N���A˗q�u�a�O�����*�
�UA˼O&M�Am�*�zNUt�yPK
    +Q�H#@       org/bridj/NativeObject.class              ��[S�@���{B�;TPEM[h�"X
H�^`xЧ4]j���4e�g?����q}p���x��^h#L�{9{�~��n�����6�u���ja?�%��!���c�ݗ�dI֊�S��a��frcOVx~��楄�Ӳq�ڧ/����ɝ�e���� B-<�NA��SO_�s�a �p��B�!�n]��:c��iCȬO�Ρ$������2CT��u�l�R�]����"|b�9'��V���3�%7�F�2FED0F3ߨ���&�ߔ�"�t�bs��ř���`��.H�*t�a�޲To3t+�V1��b�F�����Qׯ�t��5*E�s�l�g,�-�ܮ�˺a���;��MUׂ�f�u��m!�8��]��mU.֐�!�Wa��O���ve���9����� �>Ղ�m�#����-�)�1�jQ�ͪA��e���tE.�ʆ*�K|�j�Q��%8=9�jY=�sñ�ux�{|.wE�
�R�֫��7T+@8�i�Ȕ�J�W|��Tv���%�з̓�S�i�Gzwd{L3^�]�o�ŧNp嘦^���^[�U\�QM��Ӫ�4;�n
��%{�4�L@D�AX�9=x�����	v��<���uA�	��!�Y�0gg0��h�`�2�Ӑj�@B���4��I~�xi�.�S����'ƙ�g�M�۲�uj�3H��Xk�;�C}$��O�{�b_0����;xqTW��Ց#xh��� E�ٛ&Х6ЯX>Tj�`���	�"��O8 �PK
    +Q�H%�8 h   �   %  org/bridj/NativeObjectInterface.class  �       h       ;�o�>CvF���t���̔,}�Ē̲T�����ϼ�Ԣ���TvFF��ĲD��ļt}�4;3#�Vz ��\���Eɩn�9�l�L,���$�XPK
    +Q�H�D֖2  J  #  org/bridj/OSGiBundleActivator.class  J      2      �PMO1�Ǉ(� *z1F�	c���DI����{w�X\��[п��ă?�e|$��u�Й�Ig�o�/� ��N�4�'|��}�j_��a��Y��H:cs B�/GR�2ꉖ�W��!M�I�&�iqc�@={'�����ob�D�܉��;%�k�N�X�#�<!�nuL��~]�A��NZGثy?��4�S��Q���g�K�m�mbg���2�H����%OG�j8�*���@]�Pa)��}����\�q�o������X|�!�U��Dd.2��+��K(M���� ͌Չ05&Sˌ��c������PK
    +Q�H���$  �    org/bridj/Platform$1.class  �      $      mNMK�@�צ���V��Ѓz0�W�KQ��޷��nIwa���<)��ѻ��~ ���,�fx����@ۄ���hlU:�.3Q\;��|�57"ʄ�Dé�"�Q%4�R�嘰���N�)��cBugwb	�<����������v�	�H���8�C4˲���&��t`���Ub��aI��@iy�����t�+���<Un|����JO�e15)!<�Z�~&�\�Q��Wa��=��X���w��[7�`?L�k�Qw�3��w��Q��=�~w���-}A��M����R>�ːK�q�PK
    +Q�H���  �    org/bridj/Platform$2.class  �            }U�sU���eCX �7�5)%P�ETz�ִTB�\T6�I�u�[N6%PЂ���|�3�Ff�q^|��7�S���&���d���s~��������o���U���(�s�,L�G,�-:brK�
��0���eإ���ϻ*-�G*�m�,�"İ���S�خ��W��r���ߴxy�����d�3�mσ�%�������ī��u�����4D��\O���LWj0,�C�I&_u}��SM3l��Fu�)�E�z��^�C�l�!�ߴM���eX�
VjX���Vix-RZ�h���bmA�c��f�aU���; *�`�<�Y��ӝ����t�B�K���笟����W��*qw�ܮkK>N��m��V�1��<Qi4`~�0�ASh��t�,����f��HK��J�?U�I��3�*K�'k�;yBË���cX��T�x�"�4��8{�7D�\p;ϻ���=�+Q�]���o�Rq�����Q��u��k8Ȱ�i�.$ï�^IGe�2�n��<s��My<@���������r���*�)�i.rN�2�(����q�q��VL� oq4�QY�	��c��ibF���o�`�0���M�u�5�ʢ��yb�8NH'��l�����J���.�i����9Yp��S��v�y�^a�(QPb��o�u
���>���ʺ�B�ˋ�T��u����#w? ^��&C���L���O�)��Q�W��&E��p�ޥGp�!�i(�P�`��Ƞ�u\�bwtfAM�ڤ�dr���b���*���3�)śށ
���i�h��c ���؜�a3�)�G��2c�|�2�㢾�:����Y�g�-�L�qwܡ��l��j�2/cM� �����h�!�4B�+�пK	�)I@�֕��ۈ�v���Ԧ�H��`�-=KO�Є�l��2��rG����X��b��w���I��xɌ�v�װ{����``_(���uv��5�t�9�"��D��Wk��Q��������w�	��A�$��$�v�������7�����;8��N����-I5�b|l6����r��D�w'���4:�bjl���w�?���"Nb��������R�>�Ytc�xW���9�*1�ǘ���t��w�xZO'H
�!?"D ����$�u�#������'��x��l@�"�� ��CR9�N��*ѫ\�!eY�2N+W�W����&�5�{\W����N��[<T��������q������$Eɻ���PK
    +Q�H2n�9  1	  $  org/bridj/Platform$DeleteFiles.class  1	      9      }U[WW��`�z	�5\4�X��B���
��ҁ`p2�N&(��b�-����>�k������Xײ}�SE�Gj�3� ������g_��퓿���9�.<����L-�.Z�7���!iIO���!j�%#f�|��̢���(�yiD]�m�D�@u�;����顸OƧ�qF���#��ul>�ЧO'�����Z�ʓ�mz��Ѷ�0j�]C uo�d����E��E�?
��~u9ϴb����ڮ
lۨb�@���kx�+�m+�*Q���ь7�ф�Dc�}{�FvL���䯆AK5�a?��}u�K�Ex�s+*�������T-AD�hD��6��,W��%F'�+��hf�錷FL�j��5�OY�^슨��L��Di'7Z�Ӷ�s�>G6�Z�C�f�X�0m��"&<״���&٭�����4f'�M�+��L��֯a@�!Zʟ��i��v�H�6��W]B\A7�a&���$�ϑ��9ו��4�rԴ,�B�w$��א����SC�8�s9�3��$A.j���=4l�T�s"y�F��s,˹I��r�7���d�����r������I�@���1�[^�/��"Q:c9)r&Z��;[P"
�_�uW�G�s����~e;��T*|F�x���#A̒U�u����#�#1�!��[�āhB��ĢB�Ɔ��9�H��߬%eF��(s6>f��&<c�F�5f9QY�ʼ5���@u[3��u[I���%m^��4n��22Y�Rix�K�e�k�K�<�{���tl��ޤa�ؐ��ߗ:ݙ5�I�5�yR-��� �r��4�͖3/M�&�y��r.�6��[�W��ڄ�sg���R¶�;h٬̢�<�.�.TA��]�T�sM�yʹ����+jb�����	v<�M�q畨G����Tq!5U�R�L]��Yk�=z�Sx�=��m��k�x�**������]��r?P���v�(�q �p�ޅ�Ky������yuw��X3S��B��F�8�q����m��7~A��^��+�S5��a`�	N����ˏ{~��Ά@woE�3�M5U<��S�-Õ{���u��Tv���㾱R��C����Ohy�Kt7^�\�����b3�X�X�U��u��/�,�a��5���p��6M���.�Y��
�;l��+x��<l�Y�n�q	7�%Q��2K��A��'���~|�] �8L/;�)P�|F]%� >�>��%��!W�۟�N=N6@�#$�s{
���b=b�"Χz�Y���<�Bǒ�����Q|&�p���<�P~/ƙ�ߢ
|G�h�B�PK
    +Q�H/Hda.$  .F    org/bridj/Platform.class  .F      .$      �zy`\U��9�%����閮ӅfOJ[C��j�ѴY��BZ$L�I3�d&�L�d�(*(
�J��d))�S
AA�EA�AP��s�{��I~�G�{��{�g��s�'>��!":�8�)?�^�	��<3�u�#].b��;|�|�A_h{ec�[�EӨM��f�q�칫�A̿&�G]�Ô�6�4~�\�;��S]�ǔ�6����.%US,m_���P �og�{���F|�=��l�Ӥ|&���چ��7�4�n]�	�ڲrm͆���P�\ROk�SO�u�g8�{�1�ʠ/�����Ii⥽����]���v�#�4�i�o�cP�X{bO,��Dc�1w�в��d���;,,W��"��Xr���P8h�ŏIc��%ff�8+2Cs��E�:��@�jъ�HZ��\&��n�����LX2�v���L�'�*e�4�=z�=Q�&�!����D�Pcǖ@�=�;Zsf-�yW��[�quKcݪ��5jW7�Ԭ�����6�����=�b�t�zE\��&&��E��Wsa/$�E��Q_kP\*g�8�r&��x�E��T7e�h&�o�;�i!����X�g��cR,��h1SI�P��#q����ݤhiF�n��}�.:Q����C1{RgHc���'�SnZN5LD�p(c��d�J:M(VA�!��h�ȁ�g�Z����\H��I�EMCȗ��}ǝ�G�x�	�"�ҟ<�.@5Q����T\tb�'=�6���I��'9ܸ����-Vw�%/�5��Y����M꠵M�Y��P���E�@�p�?�pR���X���q�V�4�k�?���-j������ü�2��	����M�q���{!�7�l�[hv���0{���9�;��N��@ AN;���M3ԅfuQH����ݾHH���l���wK�--�j��qc�-��#�c)�n_�d�D�I�I��V�tAF0�˺�3�I4�Ģ[�`�p*��%n��.w�e'y.�����{�dd.�m� �
�C�P�/�ۂ��_{��S����t	�+��LDu���l�&զM����|5}#��N߄X�J�7��H,7��$�Z���qE�X_�9��Έ��` ���4��� �3-�]�}�ߢ��M}����\t�M$6�U6ss�D�@��4-: `���������!�`�Iy�hĄ$��gk�.�t�
F����v�Đ�`����'UuԢC"���`�&�������3L ��0�\����֢#t��z�0�谶�D-Z� =$t� 6#��E?�~i,zT$|�~�45�=�[�����,�M�sA�c�V�����$J��H����OQ��#�02�36N�Ѥ�xX@��!��/�.,�K���Рv��Hķ��߸�y�T%e�G$��Ӫ�ZgR�H/���I���.z
��E�̴=૯����w��"��3a4i�?ҟ��� o�c,z�~/���=z*O�QR�����b�@�#l��Ȗ�? K ��t�O����6��AP��^&��DB��-�X�� =�j����ν�6�{�?m��a�2\?d���+;�5�M�E��_���;�:��:�7�6Ŕ���@���w��ѿL����p�?�Wd�2cuX�+������y��μ�gs�����S�����:��6U�~G��J�u��dє�upG==�5���d��Cz=?�G̟Q[�H&�z_P�W;�h�,�N�W���
ɼ&���D{B��/�g�]�$�x�]ZAcݨ�����Z���n��S ߲@��ۧ5a�4�}<���
�c�m8�3ً�γ����,�#��E�윃L�=�i�<�_�
���*�3.F r1���7m�M�ev�Q�e\.D��`���;��N����B7�ʋŞ�&���*I,�����h�01̘ŋy	���a�m��x��hȨ�sx��O�O�����5��HI=���N����r���,�l��5!�8�T�Ю�H�k֝��qdς�m���]l=�g[LS&ط(+:|=��f_�G�v��<��ye���7�MWl�]����vņ��&oĐơ
�M�l�Z�E�糥2��-�
���i�W^���	�7}Bn Zj����"�A1:�Ns>BEy҆&Y�q+�	?����4�ck�=��4d�`�J	�,�Mu�� ��BoQ[�'��m�{}^A���@4��/�#�.�J.j�db ��e$��w�z.6y���K(�_ڳ�陸K�L��N)�uK�Dc2>�e�66��ѵR5��Q�!�r`x���M��R�H�5x�m��F6�n���D�j�/�5_������Q�?ko�2���Rۣ^H�N��y5%�P,��O����Sb�:_�!�"���$i�/~n��g𗑴�E&��ҹi̸�͗����Vj��0<��N\�G-R����]tS(�k�ˢQ���?���u����J�9�;6D_��d������R�fd�N_��~�?ԦK��o��7�Ӭz_[cb���ɷB�U���@��~[M� �l��n�	56�|dvM��芦U`��&�c�-���B��D��+->��I���f�`�RIޟ�έ�4��@ ��8J7��@ ث&��i�l[C(���:!(�!Q��G ����j�ɨ�szW��=J�9��R�.�2�	)0}�]��&?�䬊]]!8��O#�l1j����m���֘n�56�_ju�D���t��km�&h�M�f\M~��v��_Y4`�V�4Z#�����R&��+;��;2r���f�jվɞ�?X|ؖ�xU���g}�e��&=�*v�pX�Q4�T�����^*�a�߲�Җ���5����ҏ��_n~W��0E�L�|җ܎�^&a�C �L�[T�r�#�X�������*ME�JoE)��@wg8�G[���?H�Pߵk7n�	�"Q_�9�b�4�k��WPnJ�Q�Z����Zx_�1&�;;0�"�m��S�Sϋ��<����U&Z��n2�hԈS^�Cg��ad�����Գ��6'�V��p���F�#�,oQ8����BS��B��h��Z��9��h�y���bS	JI'֘r�5	���U�I�ſ��*�NIPg&��$��W�
*DY�B�	�c,"���XdO�w��P^�
DP���@�t�K��G������T������e\��_��q���U����W���V��Ad]F��0\}�M�է$l�;��
IK��Jxpп=��{Lb;�r 2��H��X���5J︱�J�8���[nt��З�	G�NV�*����$�m��T(��(�AR.���{;l��ԙ�,@��`�Y�A�m`�TD-�Y7�j��:�fA�}jk�����S����GA6-A������7�ĒG�.Ւ �_�[���v�V�&�
�+�S9����<Ց~�Jc�)'z��?�h�
Q��ӭJ�����R�]��H &Ysj?U�:߭�
�+�-(����0�#�z,�ą>{�*�L�8���R��<u!�br@�`�Xe%�m+2�t3��pOLl=���r������@$;��;�0*��M~�"S}	ؔ��z���]��՗�WdǨ�r�v�C&K]e�j��T�e/�Om� ����t������W�m�G�r���g���H5�T�BE�"}�=������T�43%vC�����������dG�����^|���I��!a��&{�fK�m~�����
�Ҧ���V��C�a�?q���2�{���{.0�]���JF.�eR����1�=Rڄ�]�r٣�PW����Rqe��d�:$��R��v�C(���M5�� a|��3�Z�I�>^�=��W>�y���b���j���1Ra�F���� [����!]�$��R����Aw��~�T���ʞh��=V�&AJS=��;���B�5;]*�<�D������0�	�E�����(0�-V6�T?r�n��-��t�����,��c(��̍�f~���d�,����Z�z�.A�g9`.�;�1�zŭ~�~7��b��<y���U��I��� ��vnD�	y�(x�����'�����Jm]�#���䛲�_3v�v����ZH�ሥ�"��?�??;Ra��wC��p�� �WcG�\Zb�gQ�<�v�w��k����@w,��!Cy�P0,�զ�ڿ���z_w7��`\�&�n_��<w�����R��4���O��5�۞,e��XO�2X��C�Փ����/�8���Ab��[N���o_�v�'#�m������X���'y��
uLtO�Mgjho�2�[4�W�C�-c�1�m�2�:�RV��b���p�?h���sWE��KZ��@L^��x�+`�1W�O�d����meL��+:��ir|h�4T��S'��*ל]�[Nk�o(N'��ۣ��I����~Za�,�E}cY|�6�Q⦸���>�Je�[4�&�E1*-��=v�E����=�	�&�c�Y�?���&�cp���-*��PZb�1���&�#��px琏q����
c%��@g�݁�j\���>�:��9Lc-��B�Wl�mjZݲ��ve��-�Woh�mlhi\Ӳ��aU㖦�j2�:��t�f�
��֋]`+�61_(qn�����G�)[�?5�ׅ���j��7�?9�A3�Ѓ?�L�$�ӝ -?�{���a�_z���>��v�#���ݤ+�j�jC!D/��,R�ED�u�Ɲ[�&q�L����Y�Wx_ ^���}��\';�}�,?���i4�7��3Ȕϵ��Y���7G��om�:/m^!劽4�b*I�S��r��x�;Yo�����o��O,��)9L�Rc#�[� -�O���
�WPW`�*:�a0CS��/�Ӳ��cM��Ǜ5m5�
�0&?�������1�.=X�8���\%�T[_�8���~�*^���kϢ:j��E5B��w 癸S���BU��<��J�ƌs)�Z`@�ڪ3�@6�1�>���d��%q:[$s�ҹ�������G���0��w�Ⱥ#?���]��>�ճ����ѡH��zh���b�t����zi���)�QF;17�;�(;��.ȷ�6��q���]%��g�Ѥ�<:�@���Kpw��؜io���zmjβu�Ԝ�6՗5�?T�eTeOȞ�u�*����:� �1[��o��<�fs���`�3�B�s i����2X�r�n�E8\ls
}	w��]Ξ�B�WȞi��˘���+`�v�S��n��#_�K��g)H�Q�1�<\�±��*�����#t�AC8�����8���.�)a.�f<v}}� �Pz�nU��-�o�MC���܁;ۄ�!���&��q6F� �F��=����8�����������b���Y_�hٱ{A���H��T:(�L[�}�������7�n/�����MF�VX,w���c\l�"­��L˦���}�I<O=B+l���A�Q?5$|�q�_�}�	�'�|���?����[��?\���J-�� Z!L��i��B��58�p�_�/5m=K��1��~�1M�Q�%,r8�&���p.�E%�RΣFEx4��2�-?q��)�|��ۼa���M~���n^'8B/3՗�ט�hn��������>*ҐP���ߜ-' !Nom駼�rۺ�Ǐ��P��-zbyb⻠/�j��� O��Y���J�l���zg��ݢm[�e���=@w�KD�O�3��3P�3I4-��T�"����u�%�MA���_�n
��$�$pU��hG���y��P���y"M�ITœ�t.����鴃gR{iϢ��l:���..�B����	.�_s�R:�y����C��~�.j6<�~yxBS]�C�˧O���R:}AuVAV��Vgd?N9�)���<[��*�QeN0'�n�悜	��܂�A>ž��GiksA�a.�v�ӌ꼣�O?�r� BF�j������*)p��k�5��(��\R�m� m=�K!|�a��Ah2 ����|W�Wq�-���
�W�+��=�w�偶Lg7��V#g.Ր���+a�5t�FX�}Z#�����W�.�y1��]�}C�`_�3���R�00�!^�RҶz��p0e� o�]�P�M��_�J��i��pj�>���~��N��wb���w���E��݀9��N���\� M�
rM,�s]C��d�ǧ�M6�R*ה�T\�s��5Hɥ�q'x5��ĝ�ʥ������i4_�����T,վ��Z�y��E��GY�f�&c��7yxǹ���A�J���|N�R�^C2�Ε��S�۔}ti�}���|O��������99! bd�DX{x�=�0�p���&I�O!��~� G����8�A��&�5e����Ɔ|����\�=�y�>��(_��K�K�+Z�+�Z�餔%���Sf��*���=�0�oӻxNU%~�D���]����1���o8���Mm�)�@���=�F��>x5��x/���(/�<��F�Wh2_	��� ���6���]�	ȿ��Gg�>��먉��W��K�FD�Mt=�B�|+�� �÷� ��C|���1��~�� �����<Lor����]>J��\��[�(C�\�L�,���˩q�vM�}�������ȕ��Ѹ3� �G���$�e����L0��]ݍ����~$N(���I8}/��]'��$8ݝ�T�p��9����}�灑x<�&y�sx�����7�0痘sx�9�4�9̉'��v渵���C�_$�|�u�9�J� ?<�U������,�Eq~t}����h��]���O�<��KR�eip�kwoi��Z��?���يi��-'�����g ����>�gGP�2��WIՎЖ���J��f�	�+AeQ�>�I�s�̰��Pbo��/��ͧdI�<����99lN�s�^��I����������Xqr���U��jRrs��Y����8�����:X�q�/6�9�xƫ7�_��7�����wy�o6I�����a(����,���h�9�,��� �����f��w��{Ǡ��h �+M4�uj��5�B;��α��!�Q��#3K-GN�K�j�Q��D͡��jS�(�
�
UDרT��sUFϫ���:�>PX�EN�݌�⣄������b!dJ]J�����*�y��H�lN��׵-�JB�ܡ�2����)ǣ8�xܬ-�WF�J��Qٙ���o]�o�*��Gg�ez�[(	�h�6̈́r��#(i�̹c2�ާ�����Iy�0W��	����դ>�WëKMճ�g�*�r����A��y	��J/.��}�E�S��BA5�)v� Ur,�/��+C�&m�A|�ӛ�;�o���=�IxhH��b��P����j)-T�i��$��S��
��U��nS��n���R��j=����T�<Z5�x���>Gm�V��;�f�Z��G�9��:��Z�?ʗ�h���`N��&�%qUQ���ŷ�F�L�7�j��6��3������2�-z�m��9o]��@� �?��?��n]��4ł��EC�̔�7@�m4U}�v�jZ���C���ح��BڤǤ.?�X$�n�-�N����t������-�����I�N��ς���U��v��:�t�mj�R;i�
�gT�.Sa�E��Լ�N���х�y���Z����_ot7��N�:��V5�jU�T�n0��N�ii�Z���ig�Z��
j��j�N�(NI��\jMS� Ѵr�cӰEKVX,��~����oLu���厑)O�8� W�UW�5�bP5Ue��f=`�!��jS����8-�+�Zi�Y`����8=��m�Ѿ�7�J�L��u�)O�\�yX�[�{T��|T�J�����hz]9����*�z[�.�1&��(p��=�v����ܸڃ�Z}F_rʝ����"hפ�0���X�Y��Kp�G>گ.U���:�W�ˠ�;h�v@���F���H}N�묣���u�[E?֮hh�ۮ��c��Z��}u��b&����}��w`��h��O�껴N�@�F:K�L[խ�S�S�S���z��t����Twҵ�.�N�Kw���C􄺏�Sߧ��az]����~zG�Ճ��X�y�|�r�oŘ�6˦��*�+��J9_{����A��>4��2�%[��t�k���A��G}+���~�6n�m�R�:�j3��7AE���{��8�P?&/��'ӄ/P��0���Bu�GݨK���S�>W��a�r�8'9���9�ok��;��f���9�˻�Glj�N�\�ې95W�Oc4��hk��p&���E	�#�TG2�FU��=��a�����/��[cբ;�k��s������T�H5�%:W�.�2�U��7���&���{��z�^TNhNW �q4�������-�1���x$��4�I�(cx�Iu���ܓ�2A�XW��I>�-�ۂ�2���p�|�>PO��?)G��}��(ޅ>�Mg��i���.V"s(�/ݫ>��=�*C�O%��w8=�"��y��yZ������_:�%���������tQ�����E9�h*6��B#_K�8ُ(���JǑ�ѧ��*����j|��Ϣ\�b�E�0)���`!l{��N>z�W���1�Lc
���2&�X���S�1Y~����ᵅ�۠z�$r���9Ƥ��UodB�12̡ц����c̦���9�%Nz��/rC��[�Kܪ	�i�ޗh.�l�1e�Yh�_LC�	��w�{x7"$D+��@�˟QD�b�m����
�2Tw���i�|��������C���\ǚ�S������{<�5��ιƠ�'�w�/S�4_FbK����- o��x�s�}��:j��yqc�!��.�����1&���=�$��v���@2�Q�d�92�@�ӌ�{~I$�~9nL=D�щč���r�ǘ�{�1K�G�_���\�q�)�Ň蹸Q�O���A�,nT2�Ǎ��Eq�ꐱ8nT2�ō凌O�ǚ7���^=JvV3h�N��n�q�ǨՇXm�����9��Gg��(�x�G揧yb-�0�ԙ�Ix�/����O]+৫`��4�[����)��)5�Ө?��v��ļ/�s�uz�� �O/�� ����}z���~H�a�?���ҟ0�/�+z�oЫ�&����F���[��x<�)��
$�ئc�@šӹ�JG�e_�PK
    +Q�H^G�G!      org/bridj/PlatformSupport.class        !      �T[OA��Z
r���*�H�� 7�H�4`�`��Lۡ��m�S��ዿ�W�D�$ꛉ?�xv۴�Շݝ~s��������Q,3tZvJ��2y��6�ڷ��v>��l ch8��\7��ҷ�"AhC˕Ш��fNq3!�b���2T�IS�����n-�����_�e��>%Ԋ�s�U�/Ma3l�=�y%ݻ?+���1�'	���P��<o�R��������`h�%9C��^��;<x�)��B�>�R�6���"&�6�?0�=i��-�ԥ�.�S�f7ZZ������*i�t��&�P5M��h�s	�8����C��=�1T�ܒ��-�t������#<a� N��D�1Ŷ��i_�/�0C��7�J�n��
���`(�A<%�MqT��%�.�b
�Bw�G�w��M%3���Cj�KC$5ei��$WBSi���r�v��SK4����LM����)��
�d��Jk�F�d2���e򉴶�C�n=�Nڶ�x����3�8�������c������V�/�N���tπ���.�����h1:��L\�E$T���ڶ�vB��#�(���H�B��Ҫ��̈́��j���A#g�9����-��u(��8��$6@{�PWxA�
�7tRbk��vV�hp}hD��*�P)�h)�=p1��m'n��H'S;:��DN�/�"+�m+ ��]�bYc�THݵ#��	s�l�}���4p��o���g2��{M�Cg��������0����S�R�x詣5x�Y��Q̕|����N��ƈ7I�q��@/���ڝ#d��Kn�� PK
    +Q�H� ZM>  	    org/bridj/Pointer$1.class  	      >      �T�NW]���6c����/)��S��8-�RI����23�̘��४�׾���
H���%R��������}Ò�e���Z{�}��|`�%��V��k���¦��f�.ʐ$���Z��F�����U��gi:z�P�mg�ΪcZK���墄��2�ƻɈHP|��#a(�EFLBT�c$Le��C�������9L���'���h��u�iK�8{�={��%�Нe��r]vG�0b����PF�G0G/&)FMsvԺ^-յ�pl�eM��q�qMA�<M�Q�Xea���>+�-5:�$!u�к�լ��JG���!c6�9�2D�
�qSP�(�(�D�k�.Iַ���z�zS�%�P�p7*�E�J�֨������?w|j��Fô����$���qWД�T{ݭ+5�NB�%�f+��Ӕ�!�pT��)ewHƔ��7����Y5�ڑ��J�V;���F��f3��jƼ�����VM��L6հt�J9�k֍Z��9�)e�xt�Ֆcѷ��ע(ľՍwФ��oD�e&����iZ�7�bV5Q�TvTKWw�ڶXՋƗ���@Y7�����f���L֭k$�I��2�VE{���%�R7m��9{&�VVC�V�mk6R�^�r�K�N�z��r���g�u����d��]��p��˟`<w��r�?0~����_�}9����
a���XF��',i�ߺ(�5�7b�x֏���3�9�x��;���܋3�z#��Ȗ��	�����\*v�b�������)|F��ڔR� %��P���� �� \�wS-�4=�;���)"dJ)�`@aBcF�ż��,�2n��#Fz�=�E$}����7�$�$�vH����̿�FqD&i��[$=����0�
r��~mC����LS@��� � �e|���9瞮ix����{��O.���g-1=�Q_�m��S\�,X%�[�m �r"�D"��$�X��Z\�8�nի�1��7����R��?0^�C4L��Yu�5���S<~v�~��%�UM��lW5�Q�a�r�,�HCrS��v���*�����0�	<s��{3�PK
    +Q�H�o�  �    org/bridj/Pointer$2$1.class  �      �      uR�o�P=X�s����pS�p��C4)2G�/�HmI[��W���#�?�?�x[�q�6�{'��{�y��_�����)îL�@8���^��Lk�`k���7]˞rY��<�Y�,��!�	OD�rG���������"��ME�5��z�vfPB;V�0���Ӭ�T܀Z@[���Ķ�J���~Z�֢��ԟ�1h1�����8����֋�#�|$��FʸàX�MjZ��TQAY�!9���Q{��1�:���c��l�H�wh⥾o���5v�0^����o�t�%�w=��|�Z�ϊ����~|���&���ۑ�I���_�8VƕK���H=�l��79���w�嘞ǃ�k�!qL7��gˊ��b	e���M0<$�C6����gk��/���d=�����-�	��~���6�,�H�o�s�2Ec�ѕ�tt�G	e�Q��*J�܋�	݇FQ=Q_1����j�Fl=AxB{2�*''���'} PK
    +Q�Hs@1�  �    org/bridj/Pointer$2.class  �      �      }Q�J�@=ӦM��>|�]tQ�0*��*���th��	LR�K7�
~�%�Ă`�w��rι��|~�} ��&�L�{NG���������`��?p�������]7����m�{}�8j0̍e�0�~;�0�SB&Lc��kb�!(��������I�r�b0�����V�#OvL��os(�j[�,��\��j���`a�a�d~����5l�Q����j]WI^�͵�_��CѕJ��;B�:ײ�x4�T[��P{�T&���A(U�LD��K������0!vhZ��RУ�a�*�2����`������(�Dy�"w
�0b�#�!b���^*/�{��a�4^KǤ1�2��ſ��VTkI�c�����e�M���PK
    +Q�Hˇ�k  +    org/bridj/Pointer$3$1.class  +            }S�o�P������1�1�]�6Vyd�e�d�tq��W����m���21���Q�ss1T����s��;_Oo�������@=)��Y ��K�i9:Cn�^�������1�G:R�E�;�q7�R�-s^�Wl�B����>�ht�dp����j��-Y�2l,��Xc��H�.]�����/��yAߍD�3T����W�h$�)M=Z4�j�8ڡ�E�f8Kz�fkYǥ�(`��
�L䰡�m�Y�Ð�*Lw�H�CZYe�J�a9dU�3qP�׸�#<^���]luh�I��@'G�������u�p{�����������J�_��k�q.��M$��	F��Z�!{Ld��X�����P��S�������sÐ�x@3K�>R��'@1?�4h�=V�.�D�e�l��)�ػS��)*�W���mZMB��R�ӭ��qL+�PJ˧��+���oxB�+T~bM�YAi�b��;�T�STIo�o?UyF��W.�d�Wt4^c��`/��Oz�8�q@1��ee��p�A5ue�t�PK
    +Q�H�Q��E  *	    org/bridj/Pointer$3.class  *	      E      �UmSU~nH�ٰ�H[Ċ�,PR�5��E�P�(h�Mr	K�]f�������ZG�ڙ~�3�(�so����cf�ݳ��>�9w������C��V'J�YٝXsL���pFcYn֬�����+<���2��PA�A�_��O��&'
C���;�~�����l~+�oVdΆ׹ō)�E�	˰���]^����T�z8N+��ϡ��!v����oZ\n1\��L��a��A�9�6������*��^�5U�Ѓn!\f����D�^�����K��W�ގY#r*��гDoP�9𤺄g���0)���n2$��s�� D�L�m��R3(�o
�1�*R� �$�qL�����a��������KU��o�¶4�Ĕ����F��g��ge������z��C�iYK��g��\�L�]N�� (�ΡQ�8Mww�����]z�q��Yѽ4�ۦmX�w\ ��!,P�C��iL|:��3S�z�L�y�����
)"U�-����]C��:��7d���K��bUh�T��_C�#�ױ!t�6�*�
��z�u��ZO4vE�f�|�a-`�»��{׋��h�c���F�ķ��sò��N4��Ӡ9<�T��R2���k�f�&g�����Eǲi�{%��'���ӆY���%��m����g�h�LJ1kێ'!�|�7���MŶ]���iWW���P~mɶ�;g5��AdD��&O|@��N񁢓0�^$�P"�'h��ޯ�OJ���XB�o=�;��+��p����L�:b��� �!\�`BzÔPH��҇$E�4���ә*�Q������� I��d�Y�i$�I����N5	�q����ǲΨ�Q�w�C�3?�K�ۛ�ȾĽ#̽������V��A���P(�u�:�.���,���;n���=�D��Fx�~x&h�=�����c|BaD���IH�`E�P+�>������d��P�~D�+�m�c�����o~>M9Tsڜ|+�E0	���,�]X�����ؖ�Ue&=��$g�~ڂ]���<�Q�,�����19E��ArgT��1t!�PK
    +Q�H 1�  +    org/bridj/Pointer$4$1.class  +            }S�o�P������1�1�]�6�ፅ����t�3�_�.�v�-3�Y&#F|��?�xna.�J��sz��}������ h�9C1P�FO���qH?�i9M�!7旼�q�8�E?2�b(/�	O�P(��yu_�
	�&2��$��5��Y=��p���ٶ��*���5�̍t�{NO�J���>�d�3T����׼h$�)C?:4�j�8ơ�e�a8Mz�V{Yǥ��(`��
�l䰡�m�Y�Ð�jLw�H�CZ[e�J��4ɪ�f�4��q�Gx�
� �"���R!�N����i�^�+�{�x���c鋷��=��ҿ���P�L}M��	F��Z�!{LT_����K����oD4
t�^��PGC��,�\H�rz� ��<Ҡ��X����j�ub��֧���NQv����_q�K�vi�	M�H�N��+�9�4LBi-��V��W(׿�	��P��5f���5K3�\SgOQ%�ݿ�t�e�_^��$�֘���X�b��׈3Ӱ�ߤ�L;ncݰ���Lܓ�?PK
    +Q�H�7A�H  3	    org/bridj/Pointer$4.class  3	      H      �UmSU~nH�ٰ(���-Z�@)�k�J�*1�KZh��$�p��l��:���Qۑ�vƏ:�r<�f!�ɂ:f��={���s7���o ư���z�т'J;�K�p|�Lh`f�Q3+*�W�/'S�k�;�+��VC��^��X/,��?C���;��`c%��F6ۨȄ�,s�[R�d�Q�rʣ��^�3�t$�B��`0���C�9���!l�����6�ų*%�^X��w'>%��a�<��S�h@|V�t�@':tDp�a�f�ѺГD��W�^d��ۢB��T2A�#/��a���-ē꒞c,+�r��C��~ʔ�:B�H��r��p��4��8��S����6����fp����������!h��6L঎qP����_��E�������Z��	Cۖ��ygŷ��W=�H�]L�X����`s�)|*�h�� M��u��瘖ݻK��%��p	��G0GQ��]��J�,��T]�Y�����)be��/Vф��@_�:r��]�����cQj�tQY�^C�#���"u�-�'L%"���^��5sN��z�|�a)�ęw��]�$тM���F���\��r˶]��N4˛S�9:㖸�R2��'d�V�f����ޱ�5'~����$Y��xZe���=R���m<��=���EEP�i�q}��;���{E~O�b朢�V�S^���K��y��ތmU�6�:���*�<�����N����C��`w��f�q�ns�?M�{)�����O�>ĥ�d҄"��HHs�т��q��I�
(��>$)���H�+�*ҁ�Ig���0�f�HN��� �v�d�I���� )}��ty��_QM�k����;:�#g2�w��c���wh7����2o��!f^+V�AJ��R��d�>h�r����?D����c��O0�o�ٓ2��)�c�[ܫ�7��uA�8�"�?#_�K
#|�6BLJ 
 �Z�����G�3}�h�ߣ�Z�͡�#|�~��OR�WÜ4g��n�")��8'��b:GR��-�(��ϼ���iv�3���4AM�I�LrDy'��_+�mq�r&Ў��PK
    +Q�H1=W��  �    org/bridj/Pointer$5.class  �      �      }R]o�0=nK�fa˚��1�t� ��N�`��Tb��N�u�B29��,�?���N�	������s}�_����N�&]O���.�A,Ts� c����w}L�G�T�bE��,�����2p��J��Ͱ���0Թ�#�g��b��"��� ����Y�ҵ���,�Xb�,H�s�7=q*�B��26���Pޓ����rj�����e�TQ@����{u%�1��SI�[�Q�%C�e���D{K(�5�D	��pS�Vq���Q~6}��''G��:��ZP7�!W�{���'������GO�i�K�8[P���<�)��sn�Kh��p�F�L�_#?�d0y#��pL7��P>�"�1��z 0�ֽ�[�ac��{=��FL�����O	�I�E:�5\��>��F�6��Kbi/U��_�t�c���ؚZ��h5�TKG�q�t\�h�E�g��`n�4�1w�0��Eh;������,t(�V���r5�* PK
    +Q�H��:	Z  6    org/bridj/Pointer$6.class  6      Z      �RMOQ=of`�Zm��P�"j�mA*Đ��D��FV��R�3�tJ�޽�_q�Ƶ�h�¥���C=oZ�HK��{�}�s��ۏ�_ ,bI`�Z�F�����ʠ�lB��c���^���q(��	]`z�D�����Ĉ@�]P�cp1�۽Î�������{�?���j�>@��Dbg���]�	�M��N}�f��p��9��L�7�!*�I\B*�$�S^N@/��qL%` /`�U���eʘA�J�\����㊀�n�ak=̽�P���ybh[��"KnKU��G�H`e����*
c��gC�u�i��v��W�M Uw<��{��p{�ܿ���4��<;���CG�[�Hl�ݠ)8�}�����-������`õ;��mN� �-�Vh9>�w�k��л˳N��Z��V�O1Y������=I �a�2�ר�Xϸ0C��9��-�m���d�¢�,,�y�+by�#f������\���0)Ï|�Y��Y)��)��W�-���\��%��y�y=ԍߨ2�*u&K}�z������k��\���V���j�g��@�8�^��I�����8.��PK
    +Q�H�D�\  D    org/bridj/Pointer$7.class  D      \      �RMOQ=of`Z�R�-����j; bB��F��FH]���/e�0�L��7n5�]�t�����M���&.޻��w�9����~���
V���Sm�n���<p�H��5B }�;U��;�g�يL����ғNO�&FR�e�-01 7��v����ۖ��(t�NO�\ޫ����+����pE q�-`;^ѓ���b�t!B������w�M����0D���5�'�!�B��	�eu3��1�ѾK�� Eq�2fدR W��JAq%1/�u�� l㏇��;��R����ڛp�H�Be�4�P
<����Ǩm�6YZ��pB�izrWm�uחO��u?����{	M�߉�B��!Ϥ��4�v���%��1�c��=��m�m~��eX�^O�p��2�ACK��(Z��_��o+��ӎ��)���)��s̾��6�����봋\�*b��^�Q��v�����o�d����.�>4��$��^���o�\���3)�/}�X��)��)]*��[~�w�4,1�@T?�&���ۿPeZU�L���u��Xg�[��h}�ݸ�erUc��ˁ|I������`�I\M�PK
    +Q�H��RPN      org/bridj/Pointer$8.class        N      ��_O�`Ɵwl�6��?ꘈ ���LtĈ8��m�������ڒ�C�3Q?��jb�1| ��D��В5i����9��O����# �Xeu�N��	k��r�p����1���C�bN�����f�`�A=.Z�w��t+H3L���p:��� Ð��a������4J�Y�w��v2$��U��1̗w��[��3���V��\Zg�!}h�=�3Lϗ���ڭ�b#9d1�bj	\`l�i�Z��������B�F�3(�g	ǰ��6T\Ƅ~�G>Wq5l�bH>�����LT���B��0=���U̇TfH�1��fn��4��b!�
-"+���0�Df�����7�F����>�ti�]�F�溼05�÷z/��;��4��|C�o��v}�e�]ע���8�[���~~��M�o��i����9�'�,c�"��7���}����(~�dr�#���8M���D��q�P��a&�ۄ�S�w$�*�+9��D�e1F�6�f0K:�%,�V����u����x���|� o�4���:;4�@z�zA3N�jգH�"+��(zE+t��Y�_d��RxH��B��#�KH��7Q�{<�PK
    +Q�H��&�  �+  )  org/bridj/Pointer$DisorderedPointer.class  �+      �      �Y}|Wu=�}�ծV�$k7�ER,���S�%9�ql�Vv�N����^��֪��`ťq��C��$@>��%N0��RR
hB�#4��H)%!iIz���ьf$�H�����{��{�g޻����;�U[�aI6�Z=�K�]}i6=RH暺��ln(�K�?4�6�o�ۛ�.�:�I��1�79Xظ�ϵ~S���5T�f�B�f��E+W4%��#��f[���c;6�����7��ѵ��� t5��p:�!�^�N������nA:�a�ڢ��g*D5��9k���%2�x!�+h(5n�G���h"��Xă�t�ȃ�={��Bl�R�ޟOd�#)�n�4��fb|�-��X.#7�Z<c�S�¥F\�B�X�C��� ���7�?�?B؜�j(K���>���^Y�X)���P>�w{̏5�NP���UceL��k�h�:���X���ep89�/��T�Ym-�0��p�\�^p`��,���L�N�S8DsoK,�͸D���`�)������"Dh���S)�*S���#�7KvZ��/G*�N�J�q��^M�,�[�]:�A穩�K���A�g¾@C�Ğ��S��ډ+d�+Y���ʢgG&�!#e�`%��&�Jfa7�����T�\Qd5���2�mӄ��6�M�߃�t9L���*H��8�U0��63�\��B����p��h;�9���;@�m0�(�����q��+:߲������]�!@G ��x�^>k���~j�:e���I\70�N3g�đ�'�.�ᰙ����w��	o�37)M�bKJh�~��?`Rb�6��-���u��d�:{��1D�GMͱG�x��@�{LQIN�YREgn=J��P2��>�;d�;MQN��gWvl cȲ�;`X�2dXMͥK��q���p/s��9k�t$3��@j ���p�;�L�+��xP{��R�@A��d��dbD&��;h��͘�.�Ƨ���o��.s�W�yL�2��.K��K�B�<������]�%m����������ޫ{c�N���L&�Jd��Rc�y�vL���?��`��e2��/ŗHp��H�r<�U���A<�/S���H~|�i�������U<a�V����G���|D�I
���T��c#C�<��;v1W�	�w֡�I��
���e��$��<Pm!���e��I�1��N*G:Ɣ��L!0��/[���Z�m]L���<y�d����|��Bi��B��2[L_c�tfuL�o��O���k2��?���P��<3�@�͝�S��X�4ܞ-��FGy�$�l�����{��)�S���ڙJ�.-;���L��	>O�	sCp��'��ul�@2�F�tj$Q��:��K�ݩgC-;KϞZC�g7X�t��ӵ�]�m�Lӵ�m�m�Lӵ�'�m�Lӵ��m�Lӵ��m�Lӵ�'�m�Lӵ���m�L����tE�`Wr4�L�YP7�a[���`<;�L���PC���d�3���y�C,��H��6�Uᗼz !����""Rr^i$p^�I�}��>�7?/�9hVa8��B�h�U5ё��	�q��W��֞Ǳ�q��(ïx�@���r�o���9\�2��_=*}xEv��5m�G?e��[�Y�;n!�#
�#2��["G|M�d��ȸ��:�XHl�~Kk����� �o�(*jМ���[�DYT�M`uC�)�EOX ��:,�:���jX��e��:l�"�F����V�ٷk|�ͷV%�*���)���VҼI��Ot�I�M��VE�o(j�pD�9G��7Y�7a#qjƕ��c9�؅�&��(�]��7a��l�mQ�_�=;SU�?��d��$z����"����M����u��C{m
����`�`�L��Mr{Hn/��{]�(A�EP��m6P�EP�P�&�F(��m�m��"<ߌ�.#��	o'�]I�Nt�ĩO�s:x�x�I��A��l���(�w�n$�$ŹG�hߋ߷��o�n�n�S��8upDot"�Y��l��g�>�3Cq�R�9�3���/���xv��v�����I�H�8�}ɽ�6�a�ىӣ�Ps�a»���GxGhs9�g�s�;v�~�s^uq���y� o&��m�������x�Y��Ν���s^5kq���y'�y��q��^��>��u�_�w��8���7�90����{�� ��fמ�8���7�90_;�I�;Ex��i�!��}L�s�K�uEqV4��ц�f�%̵��,�^�
�0׺��%�{�|_�
����{B���CF�G	s�[��0F��5HY��L�D��B���z���(׻p?IQ>�߷I��h�}��Mc�1���%�V�(늢���\4��*�VK�Q� []��>GR_ �?�M�
�� []��+
����1h�17U������.1�����^$����)`L��!%ƞ�q��nƮ���p)sIQ�U4�qr2n�>���c��a����kp�K�=6��s��2�r߫���:��K�Kh�޲�~7�l�pZ���!�����'ܪ]f��:"�y�G���v���ge�gi����G�����75'Q��B�""� ʙ�B�J���{/7TS2w*w�2���|�%�%EAW�;�R�ҡ�?8U�]*����e�eýX�*��A�85�\���Y�h��8�����w���>d�u�}IQ�U�N��
l��)�n��nE|أ1�v�^B�M�{)�b�l+h{7���j�)|�M­�m�E�͢k��h�|�������R'♛�[g�$�KP*�`���:�CM�Ya��>:�Ww=�94	��侕�^Fr㴹w���Ԝ�q%�]Ex��n���ܹ�^��)�wq�?��+�$�=�� 3�~U`���^^�Z��g���}�9�3Oq����8�W��W-����z��O�I�7��C$�0�}/mN��yx�����8���C�w3m>�����N���=9�V�Fp<��X!�B��[�O�S��t���`Oζ��R���E|���i���]J��Y�"����9u�l����$�$I�,m�#s�`O�S+Nڣ���=N�/��f��<+,=[�e��]U��I�ã�땥w�*Z�2,�����1��K���94G�*�E��?l�&Q5 5���E{��=�K���+�e�oj/����	��#p�L;����|FQ�q�"��,�+�2<i��H�)^�P<	�?�W_d0�|��e�3W$�%�c�'��A�1|�v¸���;�1�=�"�O@���7�[�o�I<ɧ�)
�[x����Ð�>����`\<�C�9�$���/(��B<M�+U"=H�����	|���[y�]����u4�D���,��}a�8b~_{ L���X�dU�7�B,◻`��p��?o#\��`��A���� ��!�p�g�������o�|Т� i��C�m���+�7,�"����n�u�%t�_b�xq�
��Ơx��k��~\�FQL"����3+���)�[ѺB��uD�4�h�X��6���Uҫ1�/B�mǸ�!=���sp�cG��6E?�����)Zo�_�Uz��R���ЩG�C_���
��1���>�yޏ�뜊�܊�_��ʖ�Q ���O�GSϩ�2�C��
��LVG�?ƿ+�[a��M��ċ�|��u�_�tOw?��T�`w�_��;M�S��ĵ�k>���]���A�-0z���PK
    +Q�H�2�h  g  $  org/bridj/Pointer$FreeReleaser.class  g      h      �U[WU�NH��t(0�Kk[cEL���b�(���"j�:Ia�0�3Z��K��/��ܪ)K\�����}fY>�=��o�o_�����������L�.&s�QXIΔ�v��-Ĭ0��[chY�����[��܊Ȼ
N�#����h��:s��}C$ۺu��(Yθ��9S�"C�a�CC<����9�ha�ˆ����b�2CG��zH�U�E�(ܬ�3��p<����ǐ�.����$CWp:���m�(�S�%O���F!��K�U<�X�Џ1�kF��)8:y�����1Z�
�dh*�\�X��HH�q�Ry��5V���(K6
�q�K"-K�iNY�$s����=��-ۥ[2�bOI�y�VSHO5L� ���2��50Ⱥ6%r�b���qzTd�� V���Ep�J���¢���3�]%�T5�t�0.K�#���z�|Q"G��x�J�L\R����q7I�:
�_��ՔV�S��ٷ*2~����]�x��L]���U���Ԏ����.�se9.�hs����^�T,�ŸN���*�a&�iq� Fn��!?�����_���x���G�CHr��L�XA���e�8��&����?��k�8
 ��u���.�7e����a-����EJ��S���ЦŚ�e�����F�)HgzzJA��.�m�14In�6��)=䩣~����Lj;`QI��fm�5S&Gw�]A8�-
;���έ8���>�'�S"�*���)�usA�Y�9���a���jN�5M�^���i4k-��&���SƒX�"gK;/&	R�,K�i� Fc5z�`-]r�ҟQ�h���3���3ڏ�>D�}B��V�WBC�_ЯQjx���h'+�r��?�sZ_����[8}�!���);�~�Y:����{�۷�~����qq���6T�d?���BOW�))�#)_��i)��6Y)���W7�����b�ڊ���G[��&޹� ���c���R#c��c��.������N^��}�d^�"By�D;��$���F�_E�g�+��|_yy��,?�I|���j�*�n@	��pÏ�D؞�����@���k$�h�pr�H����PK
    +Q�HL)�`  N     org/bridj/Pointer$ListType.class  N      `      }S�O�P=w��Վ�@t��N�m���a�@�EL
K�O]W�]��t�W|���EF"F���?���n�!�6��=��;߹������ e<gȸ^�T�x�Uz�rǷ��*��{'G��P���c�dN���t۫��'T�*c��"�YkW$$H�J�w�n�r�n�FeHl�Vc�82L�0H/N��M���6��[:�����c��Z��\~$U��q����d����ũ\~�S���e�Ľ�iS�EV���K�!��{�iV�ݭ�l�F�S�N�r�|wD�1D�#d3u5�����1L_�l'_Sq��N�t�7��$��� )���d(
�$�B�ќ�U���e$T$��D�n��$�ܱ^v�u���s�Ꚇ]3����:o:���h��n�3�m.�Ǳ��Vg�L�Q��#�ia��bB��89�@� � d)�G�a�3n_`�!�'4�Ě���id�e�#2�T��3	~OiT�+��Y��
!�B����H��N�I�0'�^J_8� �!�}#mD<�:H͇ϑ;C! � ,��R�;�p� �â~�aI?���������	�2�G�S��x+A��Y�GFs���oPK
    +Q�H�(�y  +  &  org/bridj/Pointer$OrderedPointer.class  +      y      �Yy|\U�ޛ�Lf2Y��!$iKM�k(I*���2!6���R&�t:�t&L&����V�VZ��"�����V��+↊�B�XTA@�w߻��^�$MM�����w�=�;��޽��<��o P�*�L���zR����%c�t$5�3�IE�������O�X��'��:{�FzӋ�t�&/��^�d��bۈN>y3W�RP`� gq,K/Q�Xm��\���n����f���x�W�3�&6��}��#����vXK����c��̸�gM�x�#"[�]�wC8��J�Si��Mk��L�S����Χda��&W���C�er�{ ��%�
J�4)��db
�5+Y�."W�j��pG#�eZ���C%��P1͇RL��j�������_*ȋ%�Du���vQ�٘#��U�?�}iȍ�"�HzUL��yH���^��D>�����u�Hﺈt]��Ҙ��HQ0ULΚ��gS:�1ˉJ
�_H�W�n�	��'�ا0BtD�#)��6K�#�,�H*Nc>(��ũ

�謞t`z�ܨt�cdQ>���c'=FGz���$SZ���B�R!�nM��˱B8?��w)(ʸ�`��WG*c�]��D���]>���=W���͵`���؛F�! �h6D�$�FT�\C�M:��(��z<�m�T���&���/ԩ��h�ׄSms� %���pzu2�ލ\,W4��xƪ�U]���>lD�a�ǡB�)�e���{&�,��
0a��z�"�%Ѭ8|x?Nn��)렙r���1�M&��s�Jl�>�'o��C�xOT|F�O�5ŵe�A�j݈ٴ�lvb���9fӦM�bIgw��,ڤФ�͇kq�p�.�����`O\�Z�(� �'���E��	7�_!��Q
������ި)� ����SD�C�Q�w�)��G�	}e�Hy�[�1#�����Ox�:�s3(�d?�K��5��W�p?�E��,�W]��#��ώ�n?�=4ʺ=mxO��h8ޘ����׺�7ҟ�%n<B0K��Jm���cܛ�M�aW:�-Rv���Q|�z��Ar�LC�'^�'�}]�bu�����Ha�?�
=p(����E�cq; �~g�=�H"��:u�%�B}_3��%�!%|�t�-�,�hCn<��"Oor�h7��#h�4S!��,H�^�k�VtY�c�ܨsc��ڂW��L���B��"QP�@Gl m���I��3����/͘[;��Ϛ���d�k���{E��T��DN��W�W�o�js�/":�do8�<����>u��W��pSf��#ƨ��{")����&����CY;X�3��Ɗ�.k'��,k'��2����d�˲�!��c�emL��.˺?�&�5\�u�4Mk�,�c�<�pYֵ�4y�Წ��i�X���toK�?��E�^>�
a��oWr0�i�	��B�D$�Dؿ���јB��o��v��(Ϊ89G�<G��C��|������Ӏf��b�GѮJ0����pjW< G�
�(9�h>�hWǠyx�ו����7�I�L���Z,yP�(R\xKt�x�6Ǣ��EK�W�Q�w�}���M�K��O�Ւd�&E"����{��p|)f�U��z�5(�,Eu�7�v]����¼ʲ���5 �5�5��?l�05ʆA5�@D��"��bT+~����N9J&�Oڳ��`o���y� [np��pJ���	�/��p�YnE�_l ^�EĩhW���8Q��4a_l�^�C�q��L�mNR���ߡ=[LY���V0T�}�����+t���8\瀦�:	ڍ�@����D��I�,�;���҆�����\P�&���*�*T��^�:��:�d�cLx���@x�O�Ռ�8]��^�^��G�B���8c��� [�Tl�8O�~���8�$N�I�.�8]�8]&��KpUY�-�)&q���2��t��L�s�y����;Pud�l���U�;'$��H��$������t,=2qf�����#���� �~ڜ��#[9�-+g�\9�>�8W�{��@��f���T�_�?����m]9�3+�����q��WP�[(�m��v��ߴ?��8�-�����3���$w����M�^\pd�춈�[g�d����u��e»�6}��z��\`gyF���8O��+��	s�n��V7�&���~��n�Lef+{Q��-�{����@o��\hf�!����,�Q�l�\h�]h�r��[�r�M�m��(�}�Q�'��B�r@�-Z'�GB��
)�Z�(�3�,�0\���)�ZC�A� km��>FR� �O�f �Ч� km�,�����ʫ�15R������61ڡ��О"��	��IcP�x�c�=��}c���{mʜ�Qfq%��Cڭ��e6}�x�X�2r)N��̈́�8�O+��s�W�G����[�������ޢǾ�u�s8 uڡ��V�a�^�jg�-	8�y����v/�i��Ȥ��n����b��i�Ö����(�"����u��w�+oʜT��T]2�K�d�2�O\u�M��3�.��֥B�CYj��[d.��3˺ń����q��Z��Z��|�NV��4�K�_��n5��gu��Oψ���
�J�����%�j�*��gi[G�Vs�V=(P��yhPq�*��;pՄ�W����iv��IP��Q�V��|�8ԩR��/���9^oE<v��{�M�:�����DuNRgK�N��L���K{0�&A�%�'��z���67�I8^�@M�IP?@xK���Zh�e�=^�o?n9�8o��Jm'���� O�8ϐv���|�'�xUcE<�8o��J]Aq�Eq�Kq�Oq����G-���I8^�uׄ��Gr#$7Fr��f/�	����Ox� �]D��q�D;ء�t�������ܥ��^���Ԫ[eqݴߏoLJ;4�v�x;X�J�r;j�ϐ��M���si�M�S����=0�V�MR�@R�%����A<0���$u��M�v3�}��n��CxX��2�
�;�|���ѳK߇'�?(ʽ���9~��5��V܊~��>Gj�=�Cu�-��p�s�k�ޤ (M�<~g}������snĴ9��y����~�<b�h�l�S���[4ɧy��T�g��<b�ď�ն1��W9OX��͓��l֠?�h���e��iHo'���4Zw��sjW���ye�i"��$�n8�{�݋�zf�C|��Q��q�� .PD��֨#�>�M꣸L}��Ǳ��v�OH�z�B<C�sU �L����!<K���9P�oAck(��΢�a���'���v�{�$�F�����^VŻu?B�X�[<$�E��[�^i�{��5�=l�4|�Ε�H�Q�QO�͛�7���,��l��^\�<a�O�X�	�͟�\}��3�T�E���S�W}��0��M�o�E'2�^^�/�_ѣ(��T����?S�/SѯRѯQ���ߠ��AE�EE�ME����CE�KE�GE�ME2)�`6E����hG�7����ܑ�fG!:%�rL�y�R�:�X�`���G[]Ԉ_�7r�褲�v�	�z�}xi�>�1@z�{�Y�)��k2����?J�пrs���a���.۷n���^���g0�{��r��o0��/����P�9���嘪�̹�PK
    +Q�HvQ�ι        org/bridj/Pointer$Releaser.class        �       m��
�@�gc���Ak�0X+6� ��K<BB��%��,| J��S�²�����q���Cf*���Ųjt��PD�&�½�����������%�~B�D`�-	���^LNۏ#ɋRih�ZNW/��R�b�t�R
�Ny��\W0Q�:M�p��^�����c��j�OPK
    +Q�H4���8  �  "  org/bridj/Pointer$StringType.class  �      8      �Tks�L=K	a[ Z����}�^�Vo`m�U��V�8�~H1�thp8��Jq������/��g7�Zǎ͇={�9�u�����<`�k���{�^\�x~���^��k�W/\��tu�y�ێ�V\����\J3%��?=4�<Ҟ6��_A4h��H��0��l��S�����r���NУ8!�-2�w=uޮ�gP�Z�A�Kx�P̚ɖ�W��צ�s�6áG�Ւx��n�a2��E̱����Ұ��h�;>eۛ�o�����v�p�ʑ)��1��mS��K��*���Ti;�ni�(�0���1E��*��ۍ�/{�כa8�Cm��f�ΰo'S�ΑCA�8α{�dNr���"��=�h�z�Վr(�|]�!���9������CrE��PH���ɬ�4G:$�LHn��rdC����0CB/E�t�;IW=�]�o��A�Ymˑt�՝�<:L�ޚ�����p���-��'|���@^�۝=C9���L͎�n B�P���#�D���H�4F�#3�xp�U$q �`X"�������o{C�a�ք�Y㤟�:�?O�	Ì>��7Ą>�Zyh�Q#�!&�V�1١Y8>�'
�8UQ7q��V�ä!�C�du��%<ݨ2�I����)�1��ܓ1�C�Y��j�Au�o�3b󼢨p�.IzYUCZ����3�^KD�9I��z]�=�ޔ�V&�(�ߖ�NFSC~7��e�KvC�d7��؍� svC����i72tt������p���u���ui�&�i���([�c�B�ZºU�k�A�-1���F{���_PK
    +Q�H�
!o��  f�   org/bridj/Pointer.class  f�     ��      �]	`U��>w���f!�`��@�l �BdI I��@@�G�ѐ`^�/��WQq_뾡�T��Һu���jmm�_�V��U�sf����i�_rߝ�sΜs�3˝y��'��)��$�ѹ����'�����+�i�$AGu㬆�[��%�7�t�	����s2_y��vlޒ�LnhKU7dP���3{�7w�dy1A�� iT	���7@��0����`8��%�!�ؙ�H0,3��5��x���+�i��`Df�]���y�	��o	Fef_ԙJ-O���i��`���F�3�,hMwt6�:S͎]��\�%Hd^(Y"A��@��"�@��(q���	��p��&l��ЄiLM�j@yh�*}H����oM�w�v���N&7�(�Qy8H�e�@]���9e�3zlq��c�ukJ աW�\rĒ����_5��nA]�|]�}%�'Al�����/_��Q�?r�uK._��G ��TK���k~[����(�rk�E���"�aa��f�mI�:ף;t���S]u�˒����E<��m����2�;���d[k�d'�5ُ����6u������dS��s7n���F-��6�[y�Y�������+�����_�x�zҦ����=<3�qi����Բ,�\��:��m�ɦM���%�&�ln�l(���)!��Y�G��׀GdfwZ�<6��'�v[0�U&�E�W���v͑`~Y�9���C��>�2�$P��WY���A�c,��c �q��Lz:ނ��i�u��ق�0��Z,X��m�`NO'H0ƃ�mm��ɶ����noJm፦M�Z!]��=ݕloJ%��iut%6%��Ԓ�|�щ��t*���֖�A՗�Ў�S�G�ټb[�N� �UI�[o@�yֆ�-膣c�[�E��wc+ߜ�H�='�1��ZZ����ѳ�N�8��<ԋ-8N�b�[PG����fߵ��8 D�S���l�yw1�[��TKZ� J�]���$<ŀ�$�����jm;h�l���)d�zJ��g� ����\�#"%Y7`-�&\��b���)љ]�����n!M�W��6l@})d�[���Uɶ�T3�2�[�� ��ʆ��Սg�a����Q��WS#��Q�n'�<z�.�}�Yp$��P�M,�I5"z������e��e�O�9�[p�J�nC�؂ȿe
�3H�9�+EF���f�ߵ��%e�ȂE,��%��a�ѵ�d�m�ҵ��C���s)�2,���!x��<�}֠vS��Ĕ7V�Qx��<�m��\��΀=���S��6cu�ͤ�<�^؋D�m��H5�79M^n�dzSmGs�i�����}��cS,���B�/Z�,<GO/�v75!���<�?
<B���t��5S��Z^'D$�Z�`����&� �ܲ%E]��0��x%�b����(�+�ձ8����Iɂ7�gT���ʪnDIL�%ڀ~{Z氲>Z�����W�� �����+AUVH��
�&���hުj�d�#��_�FD��֎���;�&~ i>���
��������	;�?��ҋO0��s�ͩ�K���Ԡ�7�=��_`ky��ljJ�Ӊ���nG�ɉ�dW2�ђhK�o�ڄu�#�0�x����;�4��J�K�hbV��3�|���Dk����WHE\����g�Kf�]'�����B�����$l5t������I,I�Կ�J���	�l��u*g`#K"fU��<�ecR����-�򭰃T�`I�R��G�jM��Ã��4H*�4���Sۜі�lmD�G��au*��I��h�:��	؞0+aJ8z�O��d���L���r�Z�H�SH����Ѧ���-4R��d��A:`�I�p�w�I0Ix|j{"W��+�u.��-��Q:���0L	j9Hw�3P���kSG7��Ե�ttnfC��p�,�htAjKg�)�L�W��:��
l],lKQh���Ձ������t��-�Xz�T'c�ni���to��������~b{Ƕ�*|�菪Ř�UfѬ��2L�X^nJ�ĥ���&�hLҕ��ٙ<�6�~�"3�C����6ul9�B����!�t�t����&ڿ��[�V��$(�őf+V,%C�R���U@,$���F�uKi���Y��eI�h.2aI�%�
�1��Df^�j���N��IBj|��_�y(�RU��+�-�n�Е`CT�U��<�[���m�;#�%�����-ى�F�m�dJG�1�V�@Ǒ�n�%�D\�:�Pl�=�A�	56'0nI͊�L��:ݱExW)�ŮRZ���t,�'Y�5�)�m�3��G0��pX63�l��h�&�9.m�R4�AGj;�ۓ�[�j��-Ip��#��=Ia�1��a���ܞ�������cQ.�Fۛ��0bp�A�D/QY�l��f]ݝ�.
�2�"T�و]F/�m��.��8��MS�-���#�/#�>CB�=d�#��,|���RZ���#R���ac�6l�?��a�!���[��e���{��s�%��I��q
�QgJgťӤ��p�%<2���VS��t.Us"yY��!�)���Y��W�nlO�5d.�-D�7`"�+�z$�e��+	t�t	��T�B$sx�G՞栖�u�˥+(@�$n�����\%�2W#eW�Z1kaH�bI�b��~��{%��Xd�4����K�$�N[�lmC�BL��~����۠��N49Z�.�&D�*_2�[P�����aJ��0Ɔ��D���Ji���Vه�Y!ʆ�[�+.�)ݍq��e!f_���]֜�G����Z�qS@�l�ʽwX��"P����Bl�D�ɱ^"@���@mx��ͦLgN��ˬ� 3�`�c��qAI$�`������OS<�v a�S���{>���a!3��?���̜��]
11���_Xҋ8<�^�^B!S'u'����ߓ�Mz!L
TPM���.YP7�%�.�C�o`��P��ذ�I�!O��'*gs�����tb��fK��s��|ޒ~)M��o�A��R�$�%����(���4�u�����3�4��,����>�8��	O�5��&��Gp�����|BNF%�µu�7q/n���V�7�O;d�/��G�Ɔ�J\�l����z�]����uCg����m(.����)���RaxnC����\���h#�@K������W�t�dze;�I3���d�!(nM���� 3G�4@\l�]��3)��|�H�5�J@.�q��l��\{���H�[�7��\<�ڒW����C*ż�'�,o���qٔs|S�lVZ�f�&�����A�0�X�}Z��dB��H�=A�15�B,mwȖ<�͌�E�έTK
������?�lO]h����é�4VʭPH]�Z���xƨ�'ѱ�D�C��9���姅,��_*��`��c��O7�_�<AO�*��q�l�j���#�(C�U�r�ӣ(�Q��ET�8��!O�`t�4-�L��S�i\�;S�$U��P��Q͕�8�TÙ8�D�^B�rŴ��l���H,{�.�3�0L���j��8t�sx��M�V@�6�W���G�O�/א �䗴	�ʧ��^9 �,y6Y��І��5��������E���u�H�����H	�6��6AP�S,&���N��S>
�Dgj��3a�+������~�Z�2y�^-֧؛5�f-�[�f�Z?��J-OmN��7;Zu�|�|X��X����ơ����o?��s�Xɷ8N����D��ƽ��pX6�-��"m��� �D�=_�z
SN�h+�&H8�QX���*���¶.��:E>��q:9t#�<�7]�M�;����䰦+
���8�$����쾻�xM�)ٝN��|.�7���k��Y��>bq�.u�~�t�x1B�2�9��ty}9�Gf�]=�(VN�W�B��f���Ɣ+���Ϥ^ٞ!�~�ؖv"9���ΎNS����t�g\�FfY�=!{]I�q�lv���F�<��)S��
���Z6�*��1H�{v�U5�G�ϖ���֎�6����Sm]IZ�Z
��<�ua�ږjK;�����ֱ�T�.���;�ҕ�m�X�p���Ԇ`o_�E���;��C���H��i�)1:�[�üNgoS��ϗ�D[��M7�n��A~Ԃ�"�,Gx�ae�{�r/UI}{��!?A������Ͳޒ��vy�&�"���a��+��>�ZZj����O��朔],�u��H�/��b �0��'�_��k�0L~-C��,XM~"�?@r%�oo�[H e�?��?���~ͽq}��2��8���Dİ�҈�a�(�u���A�G�C�r��|��3�x�M�ȿ��]Q1޲�w�̋�6�@Q��;��o-�}N�*F�R���'��s��D,�(��$���L��=z���J4��eR�3b�%�%�MO�,��U��#�h�p������Hp�(ܐj��L-H	Aг-�������3�
1G�Y7p9�R �T$�s�h�A�Č@{ڍ,�N$7�J+-c���Ѧ���6��K����U
��-EW�8�*&�O!���`%���*��!�
�B#ױ
m��tCmeKWgĦJ�d���;q���'ԵA�؛::���R�7�-InNY��j\:M)�m��d�Q���BDۊ��/a)#�Qd�R��S��ni!��N��w�Φ�`��4���ful{�w����r�8�&H�	��,��]w6�rZf��SB�]���`P��t�2��8�
�����T� �NXJ��rG�L%Ӽ���i�8�[	�l+�}2���$�z�nJv�f{PB���7��a�b0׫�EmIGK�Zb)-yrG�U��v�G�tt��fr�7��Iiw�`0�:����(�����7'6��u�hI9R}���A�(ѽ�9i�v�e62�@�30�z?�@P���?�Z;��G����RY����ؽ�*�̓�i����k����$�ċ��l�H�%S&��J��vǒH���g*�*^2�N���)�ST�co�������\���R�+�Ǖ�J��};)�҄	h�^��=��z�"�j����n�l�� q>!�T('�57�R6c
�n���B�I�([��I4d.G⛎+��.��Ǔf)[1	os#�L`��ڢ�LTO	������2]9���M��3�Q���؇7�$[�s��75��r�#��(��{�,��"K�B�� A�E���^L{��#�>�4�,V.�3��DK�Ӑ���jTvDnQ�"�;�q���#>8�r-���]���ڌ=x�Z�w�pWj#��(dhٺ��=���xv�+�_WWѱߤ�LU���i"�B^WGV[����bc)w�w�o�����:*�6�n���L�ాQ��+[�Aa��9�m��۝ʃ$�C�|�t1�d���$�9�b�<K9�}����GY��[�ׅ�b�&��*�!�y��LV��{�_ӓ�p�p�{����i��<�S�+����E�mߋp�竏r������sw� ��eKy�����հڳl!Qǳ"��5�>?�^�����p���6%n17cN��M�=�k�_r㾅1CZ$Z�;�/�8ħ������M�x�M;`�Q6~_�-I�;r�����lep���!�����l��J?ʶk�:�5r����Y-��v��������\��$[�D ��]S�����S���C�+U�h�~�2���@Pع&��_*_!��5�Ρ�i6�̪�̬5�Ҁ���U�1��1n՚�Ԁ��m�ڔFLd��h�RǦj��:�۔�,u��O�6��@�o��H���"X���FV-Q���ɰ�ܰ�g�-��:��\��-�E_`�T�����od][�X�ST�1�@^sl�����Q���5���K���.ȳ���dQ4ȳ<��L�^2��<K�ԃ��T�C�M���"�ٴ>�(�Gf����V��,�>A�yN�R�q'��l�h_@ޮ�c�P�ȉ�{�����.w�ۺs|�@�^�tg��Hn�%|�:O��e*�RP�B{/�`B���B��#x:�_e�U�j��h��n��κ�``��p��L���t�R��C�#+n������as�9^��m�NB�tt����d����ޝ�r����~��l�m�&�M�CEQ��q
þ�^!�`�_��F�B�J�*��n-w��΂���R�s_8����}*�uu�!�=���pw���i���?���ٔ�Ra\�~����s�jY��:Kݡ�G	��Ku\ݖz!<G￉CX6:S/�[ռ�{��-ɦ֮�-�R6��^f��Q}���vl����ӆz%�N�U��Rw���z�z5r���={��I�����N�y�JՓ�WO���^�H�`e^㕹�Ԥ�i�����%���$E�i�`�E���d[�$�}��~������-�L1L� �rAü$Hq��Zh�KbG�qe�-J����K�|CT.��4�L!>
�, =`z@�	�,4!�ԸRm��%�/Ӌ��?��������hٿ�ٿ�9�=� T���ŕ[�E$�O�ś��0���4BvP���oc���S}Y����b[�$�o����Jp����y�"����!�!�F��I:I�[ ����FXK���+Q?�q���N�����~F����_Lw�x�c�cB�C1�Ķ����E����oޣ����B�oa�1�K��}�q���&3p�Q�+�]�[QOWs@Y}]y���ea�Ҵ$,���I�c�#�[sg�����}rl�^kK��Ӓ�8jA�cjOJ,c��	�.�ç������C�L-7���zK���pO+ ��ZZ!���43<�,J'�I'Q�k�����;Q*����Aal��g�5m�\+�v+d͜f#�y`�i�
,��5�(,sD\���$�Ǣ��dc�)sh�߂�6�	XG�l�G_�椽�S�0B�1$�Dϴ�[�br��M�E~/L#z���Lm
��C,��o��hiӴ�{�C���s��R�Iyis�6��XHt�.r���w���ߛ�������7�������5�x��Z������ah�X[́)����}�aNgڥ-���9Վ��5&��H�w �>ʏ.F���Q�r�B�Q~eY�n"lj+}�٘���jn{[X藊u��F[׎��YZ�vi�X��4���q�.��l�%�44%ZZ뵴��	���0c|Y���F֤m$ڛh!>X·5�ޤ�6{�u:� Z�F��v�1x6"1��.+�?��SW�Y�omZ7���8U����!�<�Ԙv���oĖ��3�g�ڙ�%KK;�����s�U%��?���g���+��B_:_��r\�K� AD1�ʽ~���XD�{	W���Q�Zoi�i��|WX����J�~A7�Yl�vjWS�kx�-yY�.�x�m�o-�S@�ܠ�H�nb=<�)�N��
am2�$nE�i�i��zh��>1��;�.��N���7�]<Ժ��ahYĮ.�^��ik�s�~�L��}y{,�ZдW -��BRm7��&5X�c
����l�O���x�W�H����K�	*{9�Z�OqPy�_P�u�.}��_�k�)����~P�%��R+<i�-��^���r9��f G_"���B�_ /B�����-l���2T��Ob�O	��������g
~����o�4kN,�Y�mio��+�r��x������O���3+�V淼I}l}�/��Z���16f-��j����d��@C{.�L��޳$��}����>*���G[д�p�i��k��a���j���J0:�n#|��T��ӿ�����X���j�վ$V_i��W��Y��a>VdM���Ip��m��X�V�.��d�S�L��8�Q�͎�c{����V0�f>J���������\�>g��=+��<+,}�N��%#���L"e-��;���3��\����P$|��ç�9�Ls��=�.�������m�ޜu��׽I���z)?�/�m�/룩�ϧ���}_K���e�K}�+��o'�Z�WP�ʀ��noUg�t�>��sdǪ�J���>����><��-j3�M���䐀x�E�|Y��>��!P�tQE��gQ����E��R��>'P�c���h�yTr~@\�����k����e¨���ET�pއ��Hmo��)��}�z����}	�9�/�?�Q?���֗�h�-��l��������j��Z?�O�+t�Z�Z_��k��ܷ��4=�3�j��-'[�z�8���c�ۜJw���c����ֵ/��8�m��G�>�cu�VZo�*l�ؚʨ��BQ���r�N@nN��K��)l�`��yJ��1��Y��Ci��-�3'�z�%�d�|�I�ަӱ$:�C���T����n��Q떓���{݄8ђGM��V�TK�!��V%<&��X*ҝ#��H��q`���ҹ�˜Oy��M�B���~ё�>�]=���S3���H\�M�����P=�; �akP�E�g�g������T��Vm�[Z;�]K���;ŉ�&U�!Ig��p��h|���K��a��ɵ�_bu �^�v[�����΅H^l�]e���Kxy7��_�S.�{���1���:	���6�����~�~�(�|�Q1K�E��^�:.��67��0�n� y=-BS�\S����8OK��'��'"|ď���c�����
X��4�������~�'=(�<䴝�vV���0�=�#����k��(���������G��}�JY�
1Q�%f��n��$	��S'?�?C������a|"����?�?E�^@�l�T���DR��/�*���}��
�->@�X"b�$�C��bu��$Q�o�? �?䭕oD�p?�q0�[�5|؃ɵ�#��봳W��~�m����}����F�~%�׭���K����!4F�1b�^�<'/m���OX���:����������f۶����?��H��U6�$�
D��Zn���O��
K�,�3��97߿��u7p�G���m��}��ǻ���<���Y�V̪�7cr�Z��:-���,�؄[ؐ-�?��}}�yPū��:}j���A�;�)�.T��'�{��)m�<)�O'���*[���\�F�1�$�}%�H�� ������bc(Iu� HO	��ӆsۉ=}� �<�3�����_�R#A�� j��|`��nK��,c�A�P�l?�(���1�G�����2&�T��AD}:��Ӧ�i>��9b�`�'�����!$�n�r��j|�F��pC�2f�`՜���e��s���|h�ޝ�~[/�^�֠!���/�9_�2k/�?2�Zrs/��z�����?�-E�{�e,6��2T��h5Z�r���X�k��J���o'��|&��8ț]��h��2��uww�"y@d�o�9�}�Zn����$^��ّ��x��:hc�D���.��o#q%b]���dn��&]k''R�6��h�~�eb3�0m�el2Z��I�R~�XF���5����ؾͺ�f�6c[\k���Ɖ����?�2����o��>��q�q:�y�2��)F�pɀ�8�`6��}�ƹlפ�C����R�-�[[��o�7%�	:��gO����.�'�t�-�o��&}�ܙ:��`y>�a_�@%/��T\��nI!�%ŀܾSŸEmM/G�,moC�.a�@�KV�`t�S����6Zo	���"*��:N��C�*����6���d������Wא]����{�rh9��q]\�n\O�^ӎh�q#}�=ݸ	�lS�F��b�z�#��FǸ-�T��Ǒ'��@��Kn߭TQ��ow�c��nx��1J�{I����ϥ��óK��/uIFY�a��$��|��M�O7ez]Ajƾ��r��W&{HK3����w�=��Q��'����'��"��`�O���?;�K��"�Kв_����h5��J�x�>��n���[#��&�`�^�ܯ��ֻ.!��}�goP˓�0߬��/��G������'�7}����o�$����RM@�bZKR�E/�f�[$sQ�����q��x�ᘞw���m�o�0��s�E>���=	���N1�tL�V����Q���9��0�c���������S��#�n�ŕ��礫���U��KW���*��7�n|A:�����0��_$ȿ��ϥ�|Q$ظ_��%�fhcE�wn�)ә�M����o_�7-�(�
��qP�V#]���L����w�'�{}�^Sӌ���!��(�"M�)��Z�o��Z�Gc������F���-7�By��6�f�5g�(�u��25�6��C�9�6k6�(44�1BoD�p��У3tM��f�R]lI��^Id����9\�����%a	�˹�#�$�W46�i����[�h3'��1l���2�A��cHױ���aM�J4��%-m`<���%��R��ڊ鴋�S�''žo���B��Z�x.�K-�O�t��R�p�m��|ye{������4�y�O�3�%�c�ҞjK���`X���}�P�
�4��s�{_�@W��D�ɩ�r�<[y��3�ϗ���[ڹbNGW���o�X�L	�8F�g�.��F	h��h�/�$=s5���)\�1��;bv|��Z��s.��y���O,^[�<[v�E�O��eU�`���Ry��[���ьr�7w��K0a�m�]M��Ln��e�ͬ�e�)���2���(���6�l�-���#�'e�2�̥��e�<�����5�r����k�%s%��f6��"l^�*�N��&�ws%[�qt'�\C�;6���R�h�4ױؠ�s:�8G�9tu"U�<���3��j[S��j⯚-3�1��w`�pB��4s�%_"өJ&]�֐�M쭥�]��O��v��)$F�}l���$t�f~�u��#���j�i�+nv��t�4�hn�W��vvA�Mi�M�R���,�nJ�9�����;{6-1��CT�,&)ì�L���v�qT���_�&��~�3՗��Y�ׅ.�5ϡ�2��ӹ�9���<,�	C�T�M�-4O������i�nf�E�[y6������"�G+w�]��}B��ç��Ӵw]��=���*�JfՅN-lgƘW�9��8d^k����ռ��K� [Oض���]�8�b��ss���FC��Mü5	�Լ��w�����DBs��B��3�5�{�e���͛���p��X���D�A���@���+�#\��|)�_&Q�qΧ'�f��i�^���<W�.w�yu!;M]���տm��{��б��[[̽�27�e>E׋��Ө<���q����I������;���(7_0_�J�$v��%�Xj��M�6�z�|�|�(���8��c��Z������K�	\��G�(��6�S���U}������t�|#vfe���e�)d2^�N���j�?���`�?1I
}+pII����M��;qx�����tn��h������A�w_������B?��f�&�m��6[�U�U��t ���sX��R��T�������7���V��(�wc�!}e�����A���������,���$�_$��X��u7�a~>�\���7�j��{��BrRġڑ�1ĵf��/^�������5�ز,�+X�c~�ȃ���Xjjx(s;Sq�h��]�)ٝ�����1���S��id+$t��`��.���i���i&��|����F��R��c�b��}&R�	O����f�X��{3�낙rk�.X�wY�$>��UqG{jIG�
'2vF)��t��16҂������O����sd��C�؁�[$��R���ɓ'S!���������k�oN�[qH�\���+�՝�beRa\:-Vn�T�CJ��Q!qϠ���ꁱI���״va��X_Na��� 8��Y^��~�����lh\?����%G.\�h�A�L��D��\�d�f�����C��s�}���e�� GR�Յ�aQC�H,6;VM2�a��&Fl.��B�h]{W�g�uVl~�&���C�!t�D̹A���}��7yc��hfw��5%�����4&�iQ��؎DB~C+:	�)ě���0�� �WW|G���ꅳ<)���2����C�.�:�����dI�9F(Vy�z��R[:S���40���;�,,t�?�9�z�L%�	�܅�J�R�����`U"��\՚n�#x�%�4}0V��/���^*��L�;������ՙB��ur!����'�O�X���C/���0�٭/�N�X��h[��R��o� ta���?�O־��4�FV[�m}�U��ԏㆂ��V/�X�ApNY�p�.aek�lTa�e���Qi!�DJ�2 �⺟U��Fї:�+!��0f�@��3��s�$gF�E�*yh�%C�������U7f�u������Y����p|�N��XY��3�s�+��4,��9��T�,�����2gc���Ǿ�-���sE���H>�`�,
69�����r2������8^pST������A�n�^����0q���+�ԯ����PtH|-U)�M�^<������} �sz�"왽`Q�����SH؛A��C?�%1��PY�,k�W��̒x�χ}��G�cT�l�;�;n��0�Ej˔UT���-�P���J��"H��T?r1`b�X�J���6���s�4pN!�Tf�j�@/�����<}�n����,<�+Uh�����ꋘ�~��5x�S�C���rU��LQ�k".Y��HGG]����.����T�)"rϏd��#�~��/�.Αb��!��q�Q�������k^D4�?K;u��O��T�q�Y�W��Ы�¯7���(<��p�Ъ�����Be��ͭFy�.�杻O6��x�~3r��a��~)��(4�܈ۊ���he�=D_�~�S��1�ɺom�S��׆}��z]R�ޢI�EXqy� oZu����.��?���4�_������X�� S��!��aT~�Qx�y��~�UQ�}݋��Er��#��wߐ�[�����
W�ރqsQe��E��G\F4�K�VG]*��o*��Ҟ�T�kjO�y�dk_�W�7c*]z�QԕEU��Ee���qh@uq�׿��a��2�����m���F+>�3Ю��`ШQbu�5�َU����WvdWމ��{��}pht�C?��F�z.���@��#��d�����Q��l�;L�Zߌ�'��S��2�#.���C%�w���}��w4��\��k�M/�D}Њڑ2��wlRSCol�G�G
=�ֵ��Y�����1H5-o�!Ӈ'��a�<qb���hIj�6�H���G��+�:�C���#�lE�YX�Y�ݲɩ��P7sD���2���^�);V��f�Z����ZEU���GF\�b��F^�n瘘��'^�}���I����z��Y8��yVv:Dr��I���:���2�ڇzaٳ�q����؁��.6u6�A?���2�
9y���N���v�@evkV"��>vD�ՃF�"��9�{<w+���5:�J.'&���γ���N���@U_���ݾ��"v��;9|��#]_��Tھ���t��;9|F�#]_饑Wл҅λ����>k瑮������]�B'�\��N�j�H�Wzi�Eݮt�3�t}'�ϋx��+�4��� ��?M 
�nWȪĔ\v�r�z�A�����&v���L����F��,3m@�u����9�0�eWdjD��%�g:&L��L�(��A���	3h�e�E��/,�~)L�:x`���Ų�K+v�fF,�Y��H
{�#���>��Q����4�φ��q|����B��եY�ɑ�R���K㟠m�?"WX����p(�Ȉ�t�H��>B)_Ǿ'1h:�=%"Z}�_�q�M��}���.����W?;2黭�o��O��f̝fA��b�|o��1���m5ŝ���ԞݝM�E����U�ޞ�dUJ��� ����"(���A����߇�t|3`&�_����g{~W�0�����e���<��Щ�B�e�C`�����g,�����"�����#����H�w,A>6���{���Q�{9�p�7�	+a@����~����Z�cu�k(�`ᛣ*���������㐬(V���b�qHU����Ɗ����ZQ��8���]u���k
;�@�3�a�.T�N^�N�3��A�J��]�" 8��)�=}�*�'��ʞ��:{"E񲤺{"e��H	P�s�5��BT�k��鐋�~��?E
�<�U�9��H�o0�U��h�"��B���;˜;P��,�Ac��
e�)8�R��.y�多Z<.�� w��h�!���
�r4�M�� %@e'R9���*�B�%0��uBʋP/�Ӊ�����9�wA��Y�{���p}�\7��*慅�4(c*�<�L�*g�����Rдe׎�A�r8@[	��UP���o��E�w�Ȱ�/���_��ϯ�f��b=�P�|z��.P���*�o�;>TwP#��N�C�� �6��W����0V�D.$ZZTm�Z3��z\���M�{�5V��%z�~W�z1G�<�ġ�I�1G�e��Y0^���{�:1~	uǿ5�����4�j�)f?��
��b=�?RW�9��v���b}���+���G�x�P�=��
{zZ4�V0��'�S��>5�>�G�[�ԶA�v*L�N��*�k�y=�	]���֠���5T�=�R|�z�+0g6H�����`�u�A7�Snm�k�a�+�`�+Fyg�����(�a����/��-��׽�[��������c|�O��r��#�,�ܬ!�<�Fs�Q ���gkl9���G����ćR�(E��M������9E�)��_>p�E�I14���W��xd\�!�eh�G�1!�.�2L.��.�(ք��k�m��W�r8�@#��4��i\ ��J�O�G�iѸ]�^t�k��d�:�$��$�a:U:^�*���t��&�p�s�N�%�.�s��+�O��])�R��G��������#Y%�(C�K(�A�����Z�J���!��_�I%z�t�����w#䲧&����,#w@c�F0_��������0�&ZiG3o{�Q����`ϫ��\"�eM}
�&�Cx�=���c~�@���S��݅�y7�����)h�j�AX�=-�ðS�-ڈ6o�M�E�R?~	)�f��_�QO�T�b�����;��t�h}�)m�)���Xs[F���h[Y��F��U*1Bv���K�I��֤��oH����QLa�ǯ.��������{�?|FjOA���=�i�C��]��$�J��y�ͨ"j=sIE�\?"�����jU���S���Jqt��t�:����^t��@1)C{+�h?�B�G0F���W�V�&$M¿��$�N�Uc�7u�� o�t����=Ҍg����%Ԏ殞w�#�i�Li>�O� ���#t�p�[(�ې���گQ���8�=[l�����ȅxB,,-��Z{�%AH�8� ii Re@ʇ�.s�r��ɦ��^�u���I�m���#C���i5�M@��B��0\4\i�f@�`h_A�.�P]��F�o�[���r�a,*<���%�D������Fwc�t�`����=R��#i�3��t� .�a��aA���ur�\�����&�U���(E+OU��p�1X�LÌ*�'uLt~�D?�J�5U�=��Y�`i�`��)�5�`�=�9���{��J0���5|Y���HW��^C)�{�����3V�ԏK��S�K�����a)��Q+%���g��al�N�Y��ʡ0WzHz�*�G��脧@����k7OI�K{��=%�J�a�{Jz�2{�+=�k���G��
P����O�|}�g�(�P�ς�z5�K�9�R����I��zt�`�~8��/�a;v+q�k���+tPi����J�9>馝c�ao�	���5�����_Z�W�+��#�J\oa@HO8LP��g�2�e�|��<�y|0�ھ~4��k�@_'YK��D�hC�Ds��1�.(�wK?�6�vK?���*�R�R$�WP�1��U� 	�	��)�i����7 l���G�pG	U�A��7�_�o����DHWP�h�Zz�f�T3syG+Վ����d��6��6!�� ��Q�!3�&u��Q��Z9���cTI$�s��S(�C�5�7ِ?���d���E�3���"�\)ϑ�%{⾐=��,�ҩ}��$��PrM�B��	"^3������#+�|�w���r��(��Y�u��t,�q:�8nM�I��8�����*�<�
Ĥ�MPw8��y��t��1M���������Ir��1|��>�*�0z���?\�|��0�w�;߁���������㱪�t�u�0\�BzV:�G�wеbƋe�~��XI��D�R#8�Wʣ���b|\�:
��0'H+�����e��h��#���3�#ܣht3��o��CltF�~�t�f�+��Q��K�a��
F��'��S���b�3���(����B՚�=��/��'��5�E�.��xN6wA^ų��#[w�$|��r*z�A���lȃ��G"���+i���YU�\�db�w�	.�Gz�h���EE�����P9!�
�ƊwK`0�eX��~�b;4�R�{�4F�4�;FC>Ц!�����`3�И	%ơ0ژ��s`�1���6������@�E�^�<AQ�J?F�
�5�ž�J�o��' #n�Ѧ�
�W��gp�38-�y0�	�DL4���:�Hg����Ay����(Wy�,j��b�P�|�;��[g.���<�یc��=D�.��aGc���^��$c�����l��4K�-f.���o�9�3&�8���+�vC��LPa���A	�6��g��?��PR&�fe�ς� O��i�C�NL����;2��r-�epft�n��Dݓ��FE��yq���6���g�m�5��u�=���&d^/��#ج�B��5�Y�W+�� xm=͋cE��
V�3/.:}dy)�;l^��-�v��y��' �erg=B v~E�`y9��=��۱�a;��5.'��*Ax�S+������=���	t{}��,$�F���7*�+oa���<9)V���C�V�w�|���A���Q��H:ih�����J�/Qo������ ��̜d7�v�o�׭�?*~���"o�����g�s�I�����']��ENe.�Tf�z`�	��=�ʸ���!h5�-ƣ��x�0���F/�g` %�alm�" ;�#wd v�����%\�D4a��EЭ���j��$�+��鍟�o�6[�,ȯ���ۍ��(o��\ǹr�Ε�Q�
F���)�΄_T1X�<#��@�PgE/v���Y$��C\>K>[0�,j5õy/ax�#53�"6X�F�|^i0n��U�C�u�4�|���Y�9�á�!D�@΅-�,�|Tv�/~�&����)�+9��E��^]�	�K�K�邦E4˗W��?Kz��=4dv8�Q�+�������Ό�N�X���=u�f�����3�(.J�s ל+T�1�y��Ҳ��1��p{p����j�H�?	�z'�?\���^�'N��s2�cNЍ�%��k�1�ۼ�=�u�м���</�͜�Eio�Җ�Dk������;����MB3�-%4e�P��aʜ�#n�*GN����/�S�=p�t�W|��*Z~��M֠\*�,��F�#�[�#i��0�6|�j��o�T�����MPl��p|mb�)}O����,�P�V�q�p!6�8���
����!y]t������6�XA��flpj��3�����V��;�<��&��b�p [�+��<c�^E��{:����݂t�XAɗF��F%�RL��4��_��X����ɚ�X�3X��AZꍪ�����P�fa�b��V~�4od�i�C>�W�]��}��v��԰*���RŢ"�7Q����Y�a�al��?r¦_TG�F~߸�r��B�nf@ݙ��[~l�{z��<+�U�#?��(�fL�w��=���G������>(2�b�x�a�ZL��r����ߘm��2��0��af��̒£��
��`�0$h�L���ۘ����Ю�䲭
se[��K�M�+o�p��:.�Uച�ϋW���U��{"������v2���q"���A仂���
�L�FU��Z�F�|$8�	��h������\u�\}��`#�§�S3���Y/�XL���dCQ�ؑ��7Y�cL�q<�Ǒ���B��ۦt�,�yk�)��=5�7ҁ^��r��㐹H*�\��������WϜ����p���s��b���UI��p��]0t/[SQJ��J��X��G~��04�w�?�kc�9{���#��,^��|YKr��?C�3��ܭ�1l��N�ғ�Yf'[Q�;{�Ng�Ng�Ng�N�9�퍳<��N�6%}�c�A����B^l�����X���CE��Ī`y� H�&Ckl
�����@��3���/�c����Kl��_�C�>5v��|&R������T4�Q�e�`K�q�����3��+�����q�����:s�$����^,Ȟ���kS]�ȿZ��fpSf�*A���~(��		��s���F'���ߗj�[��eմ�d>��C�����g�{Hځ��(��ٓ�Xh�aW_Ѕ֜���A�<F���g�ix���L�Tx���I�`=X?{������2�YkF3��j�'3Г���|]м i	5�'�3ʟM!*��'���Y�S&��^��A��H��'v��MF�^\���
���R�����q�Y�}l���h�Qо��L�PA{��X�vi��:W�� ��Ѥ�>�	>���1b�k����;�>��?�)����r	j���Z�1^��Η{9�/���+������ɸ������;;9�%�ݽ��M��D�h�Il�6R���^%6ø,�#O�_���'͈�b�qr��Xj�Vl)�ڏ�#6��;k��K�&�5����J�]4;1vM��G)��}VN�F���+�p\;+�$���M ���Py� э���GE��ǈq�=LY*]���D�{ெ�J!�J��㻇���)�1���� Tj!���`Ƈ@^�J�CaD� /��x)O@u|4���@}|<� ���pu|
��
ߎ,�r)�V�(E"�ڀ�*qA[Ah,�v���R�2lX0�ю`�����?>�y]�����࢈/+J�p�C��EӃ`_/�]�8|��yr��m�.z�ėa�$sh(M~='��qW-+��܏2ܞ����R���r8G+��[g.��Eݽu�Mh�V4#���6����B�+ ��PF��#{�D� �шခ�=�7@��[�Ř�{������
1@���`1�]#%&�g\R﨧ޑ�^�2;;����� '~>̎_ d�e��2�[��/3k>����g���J���?+z�I�s2�9�W9�~N�?��*��g5�Yݫ̣�5�gM���~.�?�*����M�ʃP!�&�ߏ]�,U�	#��|��oa�B/�	E�1_c��Be|L�_���CM���߈��&8:~3�6�o���mB!W���,��T�5�cޭ�w�)������ѻ��3?A��"�8J��d�\���Q6�]S=J��G*��5�j��:z�N�z2=�G����{�S�������|}v�r.{]�_��(���o�(��׋���=�������Տdh�2��G|-a8a�J(�L�2�{Q�]2�c)�߇F���Bq�!����C���x��ſ��O��D<[�Oö��pF�9�$�<\v�_�;�/�����������+�d�5�u���k�@�X���*�a��P9�6 d�~�Yl�� S��}�fW��QnA����F���_	��	*��Nl`�YCA�OSX�P�P*��Qn��?B�M�hk��76}�U�g�珡 �	�*��>N�C����@�P�`���P�>}��#v�*w-Q��E���`��"u�&cӎ�"u�2��;W������?����(�n�ڀ$Q�{�G��ʽѢb*����o1Ȫ��"{��/��m7����_�ؿ~�82-͑`
���c����U�Ќ��P�����P�Fb���*ӵ"+6�H�i��L7�����"��8~��f�Zd��jS����HVe��ֹ��b��E������C�re7>pT)����Ru3��1��u�^V	��R�q��	X�4��]�7J�@���䁚�zN��DN!����r��̜"��S+�y�O��]��2�b�y��va�;����b8cb�Q!/�u'�..�Jй�����hG`*��P��=��F�l��X��*{G��������Pԗo�;g�`p=1Pt���g��R_���f�ȲDW�S��ɏ���~�9?��8�L)D{?�<�;��3
s�9n@9�vv���a�C-Y5�GyauU��� �@��S�9ǂ�s��ءՍ�0��KQ�\ a^	G���@���ӎ�ׁη
rN�a9�B����ʫB�'��
C�7����t!�1�ˀ�Rbf��?`Mi�Ӕ���1�F��br��:��u8�r�F�9!�0��̱'znf������bR}B�O\���C���
;�
ǘ_2�y!c���p0f��1s�I�b~�s�����,s0fa���M�\�*�U�-Ę+c�B�ىs5��Ęka>��7�\/Tv��ga�\��!
݊�^Ø�Ø�v�t�0湯�1���m� ;�ync��1���(�ϕ_dF1o�(F�uh���Q�{�(&�]Ę�c�= w �LQ~�1o0�p��}�c>E��:�g�1�#��U�q'V}��l���D1�1d��	�|�lB�%�nɐg)Pl�Pji0�ΰ�i�o���y@Q�'YF1�a>؏Q̧��Q�_�c����EV$�b(���A�0�*���0X����}�)4vj�0�y;a����X��0�y;+��&:��0�y��!�5K0��d�0o�g��@��P�q����L���F��#̿�@��x�J�am�\�I��f���(��0��0����ǋ0V':_��
�nfmr<�U��*Y ��Fu��aT}`�>�9���¹�0;a�C�9�<D{��AVs �ƳDՋ0T���0jξ"�j��*��N��Ո0� �\���:D��an@���ZD��������0_� �ݢ��4��0_d�0��揰u����k"̓��nb��|���%D����������Q¨E��G#�:ԇ0�E��"���c�0��D �Z@��32a�a����7t��#�|��!���$S��޽af�!�haF2�٭�w1fǘ�f`L����(�֖�:mi��1�20ߨe^��UA��@��!/׀�\Jsc0���a*3J`LK�S�b�a~�)�a����2#8�����w3Q��A�Je&9(3�A��L�̱�f�vP�(ee��Q'zQ&�u4ut ��s�Ay�p8(w��	�sG�j|>�7�:ۃ�?)e��P&�B��B�!(�f�2����w�Nʨ�_er�O��PF-��(��
s�{Q���ə(3��̘uz8���efzQ&7Fn��n,�D��U�B�i�9,e��23�(���o:�v(�=��ڋJOa��U�f��D���xY�1�0�8f�c��*��U� 1�BĘo"�\S��\{{�Ӭ:��/�T���,�}�c�|s-jhj�:D��an@���&D��an�����'s�6Ϡ�ׇ!̴��_z�C�i�!L����	C�i_a��'�!̴��0� ¼*��.�q��� �=߫.e��{����
���U��@�����"L��2
a�fM8¬�a}�t�����߈0���I֩벘�U����E����U�À�{���g��=/yy9P�gAi^.Lſ3��D}^b�Id�Wmڧ�^�����U�a�{Քc򆡊���F@Q�HH䍂�R8(/�*����*|>�o�'T�2zK�,�Ę�I�����1a�4+�ɛ)�|��a�ү�1y5��+� ;�Y��1&�
�r��rlT7eF1'�c���U�!:���F1y�`� �y'
�������(�91�1�������bL�)�|���y�ð<�8�ױ�[�m�D1�D��tgŜ
�bN�A�7�
a.F��!�R���`
���w����:�(�9s�fc��cs�ks�an@݈�	�fD�[anE���vD�;`%>���ɼ���~�;'aNA��E�b��asbv��#��0'~M�yA0�11�aN���"��?a�)�Q�2�e��"��G=�:�.h�.:����s�5/��i��l��XE�r���W��v�Q�hſZ�]��C��n��Y1$s-?kz�$V�ŋ5�?�����D�Z�����P"�0D��|�@�e�7I�(K�]@9��HT��U�k`4�����$��~OFCA���� �n������B����g��1�����&��&��������	������y_��|����ձ���H-_ϵ|i�fW˷�Z~%L˷�j��L�wT�Oe���Y�/:Z�ǫ�|��\���!7� 
����B�?��`r~	L���#aA~�珆��Q�cQ�vL�&[S���{�� -?�j�aW��i��P-?δ�3P-�>K-��g-��h�ק�ɨ�)��i��Qˇ�����g��g��E-�Z��Z��Z^�Z^�Z>���lϬ�����B�K���;Z����\-?�hY�2����L����U9oG��t\��Z�x����i�\�>7��W��W���F�A�E�C�:>u�Do@��&,�oE=���۠)�>F��4���:>J��TG�/q�t�����\����nu��P5�����U��,�|*��GL�5�j^먹%\�*���r�?��y;��dT���Pͧ���@5��j>�|6�y��<T�0�bX�	�̿��_-�W5���������柑������˾�{�i�W��,���
�L0��i;�|��oF-߂Z�������Q�w���D-߃Z��� ���ȏ `<�����B˿�ѵR�����KZ����߻Z^�}��G������f��?�-�����P��E-��Z~��j�e���P��G-��Z~��#��OQ�o���Z�j��B�oaކw�a	-�O�*d��'��:���{��v��V�=?*�7���<�9���,Fg"��G��3ξ�8�<�O�OU��Ь~v�z�}8A=��"�����r���,��t������oA6��!տ�d��o�����o�8�UGGP�]i~��+�ɴ���@(��z���X�w�N&3�	;�ۙ�v��^f9�����"اx�S=GM�u���>��:z�+,ؾ����a7���V��Ġn�������?�mY0\�}�9�}��NqH�����?3�bU��� }�ڰ����ڢ���/�
F���ދA�9j�9�}�Sp c!�`���Q��J���J��xZ�`��2����ٯ�ٗ�W�1.;R�ۃ����h����B��c2x}b�#�&��H��pr�$Ms�hr�&=k�)A�#Ao���!A�#A^�s�*��@�hI�NH��2�a�������������ό|��h����
*ky=ڠy��z��A��&�ڐ ��E-Xf�Q>���1%�?t<����!������Ȩ�����8�:�WuE�m�����,Q	
�z������{�;=1P�.Q�!�}���L����EBĘ=ZI���
�q�aC�;}�s��O�C�����o�b|���ﴑO���6l��[)�Gb\W�!BE��I����;�(����k&���L�(&	�1@�>������"����*�J�UV�a1ꊆ�!^������x�(ފ��U]]�鞙�~�?>��鞩W��շ^���iG��Q�9�d�w?�H�h�a�3Rx����1�I�J�
�@!t�ړ�FKRع)Ʒ���Wj���o2��fC��}殕�c�:H�B�3X��GSR'�Jj�?@�h�ܙ+S�MiZE3�I�C%�$��:s�W�+���dE_H����w�RC�J(F��!�[C��=TT� �c��Ё�dX��<���x�;����O}V	4(���;7�Tۊ%}�y��[�GO���DߕP�
"����oTᵯ���{/��L*�X{t�Q�id��4����� �u��3��TNmM�I��+NIU9��UUh��B[�(��OIGJ���tL���lSw�����ǰ��=��G�
�׀a���Zܪ��j�*՘=��́k+�TtL�Td�ѱ���̪�kT�8�#{�d�2{z�Ά̚�8��Xv6�:+�m��9�ħ��gN�<�q��мě�ܙ�~��H�̣I'5��)�ϧ��1e�،��u�HۙJ'5��Z�l]�L�~��`��*6 A�|�`d�k��{���%����g���	*k4��r~j����˝��2��ZN˰ZN��V�I�r���m�G�HgZgO��A��[̉��ψHi�c0��]����q0U:�"Rp������~���9\'���g�L����$�Ϸ�M���y��� � ����$piV+�0C���w��c���:�/^��%�b�*-����9�+<�(�4�U�t����a���m��?��h?�\��X0v ����+��#��n�)��z�^�!p���Xl��ϭ�;̂G�?%]�@�����޾�l������"�Ukx����Q�����
�a�]�AuX��`���e,�Y,=��7�6WiJ��H/K��<�@�Ѣ�t@ۭ�������g���L��Dffy�q*��A����ք5���B/�B�l�g�6�}O�@���iN&֭w4���j�xK^�䮒C2z�A�������@F����L�#(�0��H�@�>�n��<�0t�eH�K+����X"O���E��QcW@�?:��Cw�V���Fr:/q�\L�d�5���m 7M�*�BҮN�3a[&yx�h"k1��7��7�ā��8s�$V*� ���۔�ܦ�on��5
q��e-��Վ%� Y�!%݇)%w$��gۿ�܎g�����#�w`��A�f�����7��t�SX��Y�(��8��8����|G�z��"�%=��`�f��j�!/c��ݝ˿�MK�(���w��Y������(����]\7��������wT�Y]Me��(XarS��K�r-]M��Y�r�a�+�ǘ��\^�{J�la���S��e~@�J3yNښ�M�l�Js���r�"Ju������ĸ\���$��bo�V<Z%��2�D��+�$��{XKim�D�_�6|Qsn��y#׊����Ѧ��5tA�����������M��;-}?�TK�R�3��2��[L_u����ۭ���K���Ю�3��H�1p��[L_��̾ꓐ�Wݞ���"��_��_Н|*�������W��j� �@!ȁ"#p/������L��i�c��0����z*��j	��}�@W��V�z]��|�-��UG[rtg&_u��Wa±,���W�u(|��(��L��C��s7�̾�.�U��m�U�0��2��o��.���V�|���� _`�g�|�]v_��6���sQ�L(���������W\��������@"0:.��x�
��F�5����7�U��k�X��"�����7�W}q��W}2��`s���)�L����W܎���,X��U�����C�V[$�'}��W}7��l�ꓹ=��k:�J�0�����:6Z?(_5�U����_��L��.���\�|��fP[� ���~���t_��ܾ곹}� ۟Ƌ��d�U?:D�j�i�������?��[���������^F�D�	솎�����o��4�UH�3�� },}�6���H�P�K���d�uS����gw����R����;!��/Y�����U
�`�ݷ���?��o�T����c���񻟜��5%�nV��,�����ɲ�w��dCd7���*�@����e�|����<o޻���
|hD�C#B��/r'��^�9&XI�$����>�����>���
|�>�%������"�%4��g�����J�[x+���A(�������o���h��HK����س��j���Q�կ!� ���zqk���[�����ܔ�sS�N�`-��-J�c���Q	�@/M����i�h
x�0�orc�����,""#�����N� ��X2��2��k�F�@тP�����*\'G�x��X^��S\'��Q9��n�޼�&����0V��!Z���C�RR��ş�}�C�t�"-�d��
Z�]h ]��(t��1�m�/���-9n~Sf��#H��A�:���B�v���պ@G-	=��Kc�-z= �	��^,԰)Ptg�"�0�[Vn�~D�U�x�Lɇ�������R�Q���*%w1�5�M��ƣ���)���h��hDJ��Vdز�j���!6`�p|�!6Xq"	hG�T���B��1�7���R�h������Am ��(m�ֆ�xm(L҆�i�p8S���0[��9�h�Z�;"��
>�)�:,�Ĥv

��!�>%Wq5/��>\�Ƌ�拾\�Ƌ*�� �x�E_��`�~��`��0�	Ƌ���Ծw��ɳb����A�i�A�d�NG����Sam��Dh��ݵS��v*f�i0R��ܘ
��a�v���	�h��2�,�B;h���\�M;��·5�,xHc;Qz�0{F��SՌ7+����tke�5`l�L����1�tgO���7�T�'h��'}�4���'����:�����L�v�l��
��T�V�k�C�sP�s��]�
��<��|4�+�L�
*���J��~�5p�v-�Ю��E0A�&j7��F8[�	���j���ڭ0O�3�'ʔ'ɧ��[�Fc�Ҋ�-:��J�_7����K� ����r�����iO>�`]9�f#���&|��Rr虙�!����S���t0�9�F��aީ��a�UB~i�ƣ�L��@ՖCR[���i���R���3�i,���7�g���i����]XKӏF�h�=H��e��E�f���ӢRh��Y�^�����߄���(j;j����?��ʨ����w�z'���2��� Y���Y)yvJ���M��uj��,�""w���>�X*b^�lVY��4�A�D����U]�F8����y����\�����V�S�t{�_���2�i�@Pۍ�g���7��N��&������\�����d���R���1�2'�6�H��yڨ�n0�k7��F�}�h{З��r� ���<��(#%;F�,WG�[f:�����B_n��7������I	ëEj�Q1%����c�h�K�p���ѥ�L{�h��"<F#F�[��g%j_�N�����\7�bإ��فU�˱T��m�&���&��A�<���0��օG��|5�p{,�lŴ�&���8#�~B�gt�@��جD��`#�� #y]�#�1�r� #i��yS\1W�R`����KOo�{���E�yR�e�8YMV����y�[=� ��`Y�@i�:�m�@֟���a9�����	�l�rr�E�(2�Y���Z��?(؇�~�<�r&�T#i3ײ
Sn�0;�2�05]Vho�3��V�d��_�H��t]�I�1�����Dky�ky�k�ȓ;�#ײy�*G+Qْ�Z{yp ��AP���a@p����`��23�6u%<��k���9�]��~2�X2�K�JI�ȞŎ���'c��K2N�]ަ����$h��$qK�mX���\��S~4>v�'��R��gi�G���b�L2��&�CP�Fl6�R]d�E���^
��gn.^],n��h�����ᚨ�FR���Cm�|�h�ػY��b��@y�
�
·~�?����F����qA0Q����@{�m���r޿2�k��YI���k-jz����X����vj�΍��-����^u�?���P��!�z�cv:y�ә�{���Ή�$GMP�}��5EI�Iج���l�x��x���;�:����9`�m�A�\��0(�0�&c�MP4����V5Y@�rM�4��4ج�A: ��gфn�C�鰹�m�y��ǌ���τ�ʙt��M�y5�������nf��MgM}jqZ�d<���7�q3��b7�17�������^�>����>�c��qܼ�~�{6����gD�h�O��Z�ldh%n�o��MH�<��N6��ɍ���-1�Ϥ����+�͆�=����ܸ	17ҫy��ҳ�잍�6[`��j�fo[<�P�P*B%�;��:���aP�'��zUoX�M�#��d���f3���Zl/��ل�1�-��L��klB�H���3��	6k�g�T�`�������g#�<ɉ����!�lB�0��<TU�:��CC's�|����&���/}mCM���d�]P�P�I�xI��}G4z���H:�o�f[č���A#:�S���lR��
�ZCo���,��J�	��4d��D��\,�8��@#�A#2�p��tPe(��PӡFL���PN������v5��E#Z�TY�T��nb�J A^�_�$)�-$yI6W��
�JL&%��Qy�UGT�F��,�_�ȑ��Ƒ�I��#,�Y��ȑ7�x	Es���"E���CM�GA���C�E��@�FѠ��;vn��)��͠��Qn���)�6cD� 7�#77y!jb�E1f���{6^��Ľ/�uj���%t�$�MZ;�I�s�t
�H<�D�@F"72�[@[��-A��dCF���(n0y�<1��\t| `jQY�FY��qJ���ɑrΑ�.�o�$�%��N˗��k^f�T�⩚e���q��bx)���̲�9I_B���B�/�8�%�O����w0!�=L� g�~��Bl�do��o�o)r���� ���>�X]J��N�����0���3QGɵ�G����$h��t������ x�.'���� O��TmJ> ����<��*0�6)�F'���DA]�����ٓt�Fɧ>�Rdg�d���܆&36Ea��M��N�����$D�2�w����{B�~$gU�؝���((>�oc�a (�4Cq��le3J앻��j(�����U�s�Jˤ��VB�Pկ���U�&��'�u+�f")��6�H��W7��Ӱ�L�
�譟�6F�g���'�lSgo)�T�ҎؚR��o&�ҁ~��A��`�,n�����W:eQ����������Y;���65��Q�7��R�C�A�t7�s�!oF�c�����2���~�r���9^�Qs�C�r�5�1�U�i��.)�wkQ3��ll(O��8PS�5[��G��.X�OR�dCM]kQ3��<��%�<��7� V�Y`3���$��;��gж����N��_�A�K�]0Fj�WY��Ъ)�)l�(C-�F?e� V�?�&�|���PFf�͘��f?	Z|'l��v+c��Q�?��QJ�o�A��`���w�EP�T�=�;���pL����\�,��r4�	J�7���i�^�V����ܽ6��-�&����(7l.�m�asx�+��ʩ�`sQkasqn؄�@���'^x�{m����-�6�>hD�hD�ш��0;T��M�t!@Yr��$K��O�^ez�zm�'b�g)32�df�H>�}���F���k��nS�M���4t�rΡ�Q.:�6���<<���-�[���~N`���ɔ{ZYJ�S��Men�9)�b� Ox�p�P�$���S���{�C�e��2W\�&��!d��ɜy12�i?�,!ӯ���d���,��9��!�	sӻ�Y�
8�X����t�;��c�����e��k��3�HgO�aϷ�Bڃ̺��c-'�yX�H��T8���i5D�s�\�D��"+Y��6����틻R₥�.�=�U]�Wo�C:_ϧ��{uuʒep4��hN�V�ED�d���ܪ�v1���-(:���B�OW�}�B���3,>{B
WaE���;EW��)�v�����V�0�Q6@�n�������)uy!9zÂg��u;�[���˅RX��	�P�*��]>̇��\U���3`���1n��ݏƖ���L����+@�Eᕠ�WAi�oX�����������5�:�ֆ�ö�x<�0�����&�2��eꑘ��+�r�|D���*r��w�}��̝8�;q����&c1�ąw ӞF�^�\�D�J�����;��%1SQ�s�>w[�%��m��a[G.M��jOԃ?ޗR��F=)e��b�2���8��up����b�"քT`0��K��YRD�"�w�~��E�~��wc����N�M(wg`��������z=����C%����s���{v���V����Lɐ������h5���
V���O�H�ga��f(7��'�( ?�2VI�-����&(7�������EE�j��w0V�d�^��ꕿ�W:X�2;�䬾Y}.1J��w���fV?}�Y}���:��Q�(�=��H�G
�2R">�$���HVG"�6�m�8<I��H1�i_F:�LE_�=Sy(#��k�#]H��3�z-g�ʙ��#�A���ܣ48Y��z����~3��zD�C�6�"�`td0�u�<��՗"\�Z`u�Q�k�M%l��ꋈ����X�17�#� ?2��hY���[�����{�Ց:�G&�	f=���1��37��'�( lqo/:���,��	���-��m��MEV������2V�Mc��߉�k�^��ՏsVoEV_D��d��{���{=�7�
V���>��,d������? �/FV_������Y=Y}%��*d������k��ױL탙z��DFVom�o&A�/���8���� ��X};��/��G��NV�=������������w#�W#����"��#3{�X}%��ܬ�1����:d�z*����G���Z`��-�z��:o�,�~����ֲ��	;8VoGV?F���������ܬΞX� �]��t��YXm���O����0�GS�l���0c�>'�7-�պ쥤�Z8���(]�)��F$��Y���y$�<b�&����VNhQ�:�\6��l�3��=�uBB��j��վ�P;���� �>�w!�_�R�
�U���#�C�țX�߂"���Ȼpgd/4D>��#��)���c��>�|���/f�|�匄~�m�&�b�/��
�t~��;3����t�@>��|��r;�"���!������%��\��g�4���9*�U� �B�h>���h����U'��2:X��lƑ�%;s�$c�Џ��Kfa�MPn���͒h&�?9���K��-�Xb̾*����2B�9Ѥ~J�.���FJ�ki�v���?��:��~F/�}�7y�@z��o�<ݓB��4C(/3����
����""��!_�?"�VDQ�7E�P�فO7'a%Ιh�Q8��r�����XFٓ��m�=�=b~ED�f6	�@	���&rg�G(��G�21��u�A�v��h�ht�����A�h�v�c��aB��=�G����*�?��E�aw�?�������� :��� :g����"4����}d��E)=<�㩄w2x�))�-xo��>�'A~��N�	g�>�0���V{����N�T2��<_�A�}d����ȞX�����m ��&Wd!�MPnb��1�)e���!-�_��7��C��r-1J�
/��+�T�w�[�o|K1:Yp!��Ȃ��4z1�G/���\d�epIt̏·�ѫam��E��ǣ��Bx=z=|��e�`t*g�C���.!A��3�?M�q�9��b�P�˰�����[��|���@���v5��}����`tt���eVߊp��Vg�5g�1���H%|���7))�m-���X�Y�(��ttV��X�S�Y=�W��Id�Sd�yJ���?���r�:{b����!���YXm�������ȡT�1-�����F`pV������������fV�zV�+X�Y���ב�o ��DV���~Y�.�z�z/��#d�'��O�՟!�?GV����e�0꟔_2������G��F'�U!m�!�Xs�sc��V��7�Q�߅�1/(�<(��C����08���X����,���Iee�]nU�i-F�M��-�%^h��d�@�E�e�5�F�L�'�`5�^l*�j�j�i\L�� ���)iQ��D��C!1�j(�Iٶ�ła���J�3�0&�D�	e-*)�O󊝉*�����SljX�X�푴��X!�:�Y���s�ۋͦa��'�9�����:�&wj;�$m�2��+�a{5fH@<l�X�v(b�=d}�*9$-��i��� RH��g��O!GO!�B����3��6k%������=xc��7��$�P�R��������x�|U������Y��䯑��$�:�s���dTL���9���Q C��=j�I���6�B����p՗��G-��J��n�}8ܬv�g�V�i�R�f0'C�1��n���[�!���G����3��m̉k�0vb�����P��n��v3���5�[��؟a^�6�:v;,����è]1fa��IQњu2f��I�)f�)U*��Y�ˣ{�����zd}��$�D��:M=����=$w���#W�^�ݠ~r�Ӌt?ҪsT�Ջ�V�-�>���3N/�_�F��y�������(_Kb�^R�yi��5/��!�NQ�
�Ć�!]3:D�y�'Լ����-1�dƘ�~��c10)��ֶ)4���i�3�� ׅ�Gd��$�w-�="�����I�ؐ�±��dЄQ���$��ƦB�\B{b���ԡ�'f���X IF{b&���1x�/`�+�Tt4V�aPM�R�F�3Jcu0ݐ{���E�\����r��
����*�����c0!v/L����w����؃�|�v�6�����X
>�5��MĶ�Ŷ
�c�
�cۅ�c��)�1���!��^c�i�Z�Vyl��i�C�����DZ� ���g�l�����}���˼�^�faj]�],�9!��Ա���֟�RO�뫦���{I�D;_���K�j��sv�L�G��qa����|�v�Æ�Ft��&%�P���i9�/kY���b��.I�SM�d|;-�-�mI���ƴ�;�n����Z�D�&���Mp�Ш�@�z�^�Ɠ�p�p�����­��Dh��kvj�
�RwV֡��^=�n���w9n�l��pa��pKG�&K�w6�Ш��ޱ`h�E���c����W������CC��G�Mx3�6�a��_�]A��'���/��N�}����0;��0'��p}�3aI��1���.�_��z�z_"k=H�-4��r,�� V�VߎE qsJ�p�_ �	�2�	�h�E�4�FkӲčׄy&���e��<S����X$F�S�N=�y,}��~V(�&�b���)uN#w����� kp~��f��8��c�WAw�D"3�Hp�-< �?|���Z���	B��
���)��j9*?���?I�(N�o�Մ$�ߠ��Duq#t#��,W�Ax���Q�m�~�������l	�RDەՈ�GI�l�H"?z��HM�W�_�{����*��Wѐ'�Lf?yꪼ���rW�Ѧ������w�y�S�	�T�35�Sa�!��zk�M�����~��Ph1Q�F�*R��H��Y�F�¿�u����J\]�5�A�g��P(I]�u�W�����v8ո��.�p@$;G�*\�^'���~V��]P�A��x�����/\5q2�uӇp�k�Y8]����g/�䗤.'�I(Ķ�u�a���o�=�w���p|�0��S���x),�K�aY<	�2x ^��
��
Oƻ�s���B�'�?މW�Q�Y�
����xoA�Wj�h�0�W��	�x�� �G|�P,�j�C���a©������Q�E�an|�0/>FX?VX?^�=>VX'</��'��Ov�'�������'o�O>�O���&|���S\��p�WI|�+��?�52>�U?�u|�|�ix���`����,x�e匓.+��]�0�v������5�>�ݤ��?�x�4�$щ҂g05����5
�S���ڍU�v?�#�\ۥ�M]��z'^�:���7��7�K�u�fq|%W�����=��;N�rͫ] 
��W�^#t��t����V��w��f0ֿ��?T�V�V`+�:��@�4��H���S�2߉
��s>�ף�-F�<���	J�K�[��0�#��XrkPs˳h�s�4�N��Fͭh��V2͵��[�]s�C���5�9Ms��֠�D�=��kD�=��ی�{5�N�������j��h�D=rғR�o���4٨�-����w`x��9uò���p�^�J�\�;�;1���|N;�K}(G'����䋛{�"P�������H���A9���}��~��=z<jc�X�kr�#om�����
Cߐ%6�-�gɁ���@�C�	�瀨N曵��vx�a��n�l-���Z;x͞VO��7�:4�M�3z�h�`�R I�O���a�"Lx@Ix�4Q�	F�t�[Y�z9�v�5�N4c����n�G��`/���rD0��@�Dz&�af=���|h	9AmXBڢ�7h����6��y:�a�����SҕщN %J!/q��OtA�[�I&��դ�ĝR��˲�s�������C>����߮>��_�V��q�$o�W��r3�I�@W��$̂ڇ�2%���ɡ�d�E"��c�x�j�5Q��R�}�w�F�_�y��sl,a�3�y�}����A�D#_�c�Y�I�Y�Wt5�q���i�w�����<Icy���H�;�?tpH��F��/����<<�H�XG�`�B21mn�M԰�{<��9.s���`��*���g��<f�k�-�M�c<������I8���!5�ԛ3�ѓn� w��*6���֌w����6���n"K�X��՗��Y�Jj��)axmo^MI��)�u{U���cC�TT��L�8�ˋ�n&j+ȣ����i��9�$��>�/�� ��{l$����Ǜ����𿔺�o��h����nP��A��&F3U�w�֣Kӡ0q3�O�l���Te�t<��Ϩ"�,�XLP�뚲G���S�>3w���J�'���p�/p����� >2����U#q��q��+0�2t�G�Y�^ų��~Ć����������|�Kf�B��\蔸��2q9K�	 ������k��S�W�\W���I��B>�������Y��.Y�Q�.�����Os;
�;����5�^��I���#B��4	G�SBY�Vl�T�m$���/�,��ɇ�p{������Ndŉ��X�������SK�㑝�h�x���5R`ҭ����z�1	���~L�'�$��B�"�4&r�aB��4����"+�0�1��4G�Hc�z���+G��zˉ�v�,oCl�n�Ş|r�;����
����-��Mb3�[E[��=
!����+(�cѸ�y#%�-^��eHÖO2'WG�;�V4G������N�'��%t������{
�A'�u�� &���ē�kq�)�H���#�0�Q)��w,V�@uL���/A��	��3>�����ѩ�b7�Q� ��5�(W�N�Fه�;�}��Xw=��@u�9��	#/��%��"�(S��(�ķ��HDgK:�4čSLّ��8�b\�c\�c\�َũtxx/C"�*tL�����AB7��iy뗕�)O;;}$}$;�q��41�'�wIY��c�<ɲ��Jy�����tr{:`}��Pqx�7���,pk��U����N�9c�ڤF��&�v{��1z�jxJ�A\�p�PGpwy� &8�W6������S�N*^/�o�tk��\
t�@z�\�����<�5Ou���g�zׁ͐����ޕ�A�;f����&B�fe(�; �c	�a7t��`���/6;c��z�z'�u�S�S��.(?^x�5�!���k�q�"G���Aj���pv-e���d�r��BWl���PK
    +Q�H�� �  �)    org/bridj/PointerIO.class  �)      �      �Y	x\�u�����lK��#dc@I�7l��$�AF^�dـI#y�ь��`��l�:I�8	I��	$�ؒc��'�@hM�4m�4�IӦMKC�sߝ7��'Y�+�;��=��s�/���',QP����zc��=M���H"��dA)Զt����h
"�M�z��ͫsY
3�y
�9��\�>�=:4�8
�̀`)̝����q�����5��4F�S�Obߕ�%��+L�b*4L�=���f�(W(�a+,����@"�/hg:�S�B��Ha�$�:"�m�p2ؿ6��p7[��]69��������<��\E
�D 6L�TavF�ła.�I$,��D�}{8�����Yԛ��k�nv�t�ne�������`d(I��<�*;]ڃ��n��\f���u�09�*[2
7�E#}�X����yU �{C`�fۦ����Djv��4��P�HvL��2Y���P$�X��X;�yG���m#�ںm>4a��X��EX�A��P��Z�Å6�2j0_�U
��!.j�+��n{��l�@��6��s�k�q1�s5����RO2K&2�pT��ia���j	0כ��~/��*+5��j;�v�F�a=��N*���rܦ�U��]Ի?�dp��F�Y�\{[r`@ܺ'9��H(�dk��%i�[#���p4��o�8ˢ����������J+��C���d(�/�֋,UX��D����X0��j�@5�H<��k�5�pP�=.�̔�b��B���HV��a��rX&2�z=n��Je�e���u���zY�}YS�4i��`�%���S�6ׄ���=�en����b;��-�To�KY��J�
j�
�Ba�6)w�l�s�����
�^���7�֘�ID�5�����RU��aK���F�x�U��z@�v)@
����E1���.�P��aA�;\�d��>�/�~� B��sL[�`�ͦg�O�v%uBɘ0
�H7��Y,�pa��́X`(H\W�x�����_�fy���-�|̇��aY۟��e+H�̴�B�$@����nR�>|%ʧxC�`o\�>|���gء	SD�6!%0#5q�!u�S�;��&���^��/����!�iĝ���b�֤Xv~��d�kS�����a�)�Y�|�"j=��K>'6�����wY8�9��i)�Q[v\dm�L3�"��-zND����ow &�Ӷ�"Zg�k�8���3��E����f�?��k�ߴ�������F��@D�ߵ���p�Py��ه�H��1���v�]�o����n���D��G������S��X��c�:�j�؋�oeи����/f��Y���D�@ko��.s	2Ű����?cAǂ�B�d\
J��j������h'�mj��tF���_���ty��i_"K�[c�I}J��8d�W������7�H�ʿ��l8����>���8'h�E�.�3*�ҷÇ������ɓ�<P�"�p*��I���w��A�&ѫ�q�R�`�*t�)[�,/*T�eg~qYʫg�Dȴ�U��%��1�3�Rӽ��%�d�T��D�8H}������G�JO��dt��p8�|]zh�Sj�Y1��.#b��:=VYk�����h3s`�m�x���ɧj��P�2W�j�;��j�j���j�;�jm�:޼����Xh(${�6��͹�N4��E&�ֵT#�u�/+I	�X;�@�9%Y�i"�N	�e
$�)����t�S���E9{R���&�T������ܸ�[����L���9�|�J=uT+�?��d,�>���m���zG-�~�L�?s\��.��ټ֧��'?�2-�g�n��M"ȸ��Z��ڒe"9�T�GmAEF�2��>�'�=��,�:����Q;E��+;���ޣnQ�2LI[�Fﳔy�d�%�1S)),�����h��Bg�/���d�u�;z<��k�;C����Po0f8����,���Y�r��?����p��
��&�p�r]�Ҷ*��VO楻�y�8��E�fKܯ�.{��ɗlU�%���Т�_�m�]�}oW�I�&�0�6�{���c���a֜;Y�݋S��l�Z�s��a�����ݥݭo�����ݛ�����1gj��s��(Ժ�s���8U�20��?��3C��D�U�\ne{�N5f�N�$����>�&��'�)�֧�Vn����u	I���+���ׅ�t�uD"�o�x�|^�X����fȟF�T�<,���X���T��_�������T�{�3��?����� 9�+�s���y�p���V������ch~��|5�_�������Ҕ@�Ӕ��W�����3�5��v���"�.����`�a9*p)fc�T�l5�HW{�~%Z����܆v��(�u�J�kF�QY0�����8�K��5�\�-f	�����%p�����Hۭ2 �|��V�^��c��3���Q�(�n7�G�?���E��,\��jW���:W���:���!�E�,����8��n⿫
�W�)<�ª,��G�����9��EKG��Hz���}��EYʝNHʹwIR�8t�7:��؇��D/���0c��"3Q��w%-ZY-m,�Vp�YT����V��~z��N���X��t�Rɾ�8���3Iט2ҹ�D���N�e"�e\�z�P�ö�7]i�#�$õ'��z�z�o��~�m)�".�����[��(���>��k5�
Y�e�+�qW��N����q��7�^�X�P��T�����9n���!|�$�ո-��ɜ
�m&�7�-�^g�i�+�/n{�5���u���i<r��Sx�0�1�����q��auX�I�Z�?���Q�׳}n�t�ލ���+�8h".5�������l��b����F<h�ĵ�G�^����cY��c\'({O�;��1������ɴ�[d;��!|��ݿ�##`IN�!0�u~_0_19d�>��&<�ɣB�h�c�<)�)M� ��5���/k���䫇�������zv��L�a�Co�V�?�ɘ��&q>u�S��S��kg�J����v6��;٦w������}��'�s����5�[D�w���Y�����?�~����gP��Y��*��Y�sb��׀_��u������[�;�������g���-k٘~<lpݬq��T�ѳZ��_�<g�~���4��7����O���W�_z��y*�}��� �7����㪀�d�*2�1T�4�*��*T�í��4r;*���`w�e166�Ƥ���F6�*�IU���M|c�'�gv֟A�@7	���6�	�+w9���P��|�5����wBUa�N��vW��f���f[kS&i��<��b�N��Z�_��n��L�KX�o��2��7y����Y�ŷYD��=�.7��y����C�����x����&�H��(��ٶ[�Q��#k�.^�@څ��;�O��~Z�v�8�m�3cq+-�Y�ȶ�����s�,Nf[�m,n��yn/d[��X�A�yn/e[��X�I���,�f[��X�E�j7�W�-~o,��.jA��;��Z\�fqq�Ż��^=�]P��e���}�q�[��e,�E�j0��~��Z-r��Z�Lc�ԙ�j�3��
g�˜i�V�i,7�Q��|��ݪZT�X͉UK�P�JQ���JM��j�2Ԫr4�
,S3��m���Ɔ�`�oPs�b@�Z�%�}!o�}L��3���xm?"�+��[�+����j�N�B��8/�;��*n��r�j2��i�zC�%�ӒM�<aK�Ғ-�<iK��%[��-�IK�5�K�亴d�!�ڒ]i��|Ֆ��%M>����[y��R�Q���C=�P�9���ŽLQ���W��{y���G8(�L�(�яaG�5�[Y�7�dڋO3�<e?ë�c��85��g�$ዼt���9<�Q�4��a"x?���c�0�w0����`���5'a�����H=��*����U��R>��9��2>+���g������\>��y>��PK
    +Q�H�
�r  ,    org/bridj/PointerLRUCache.class  ,            uT�O[U~N{�[�:~�Е	
8(UJ�!?����C��.�G������`�#��LLLL�	f1�I6u,�8?��G9�soaft��9�}��y�����`+�1�n[��؝�Uv���{o�(nJB�e�x`���������,::�/��*/����#k��(wvZ���q&9Û�U6宀�
49����rQ
������R��[5c�$Mz�1W�*[�C�١U���j�����"x�	>�t��a�m��+��h1�|a��%�z����+�n�ٴXb�l)'j��`I�7�M�W��
�YӴe��ÃKgc�+�C5�oH'�&�_o��0��t�ܑ�vK_�`Ca$��$�ɲ���0�)��Q��$hʢ-�%�̬��e#��q�hBU,���W5��!q�2w�:d(,T]�b�-��pawQ�����L�T����+qbt̒�)k�-�Ӟ��٩���E0��0���䭍2�l�6W1�j�U�Fiհ-5r�0K�*���u��;��)�s/!�3��)�guٻp��O�'��_�l�j�Wv�\�JR�e5~��� C�w>��p�h��/ h�R��>��Lϛ�l����O>E�/��Gs�w8�b����d�ē�?�x���]�,�^/��p�^������D;��J��0����aT�Ԥ�2�ŵ�{��#�
��(�R�?�q�Y*D���E�����F��%{F�q�~Z���Gq��=��cAYc#?"U�p�5^M��Z4t����:�ZCy�oRX{��s�{�)m/ ���J��\<������c��B'�!E��p	o�$Dy>�;<�y��x@�te�rO�<BӮ�G�`��A�=�_��P�Յ�rM��0�^仌��'�ڱ�(׫ĻƨIF�0��OqM��Ƭ3n�:v1��1�=,��r����-�6~�r�����R�"w>����=�<��r;���$�i ���4�<׺��iR�/����i�28��ЁǇ�_��^�!W2���w��}��!4���PC�A]���n��PK
    +Q�H�_k  	    org/bridj/SignalConstants.class  	      k      u�YS�H ��p�A w��퐽�%�-�FA�]@.G��u�]c���V�!?`�V�5ck�Uy��7��i������ ��X�r�wPl����b�t������N�h�������N:E�y���O���%z��LV�T�C���Ր�׉'�#�Q@*�IcӮ�]'$.�X��iB�ꙤI���#	)˶I�2��T]�5)��0FʦΪ)7��l�S��%�Utm[��n�&V$_FV�{D20k1qZ1t�"O�ł�����Д}�S�KY�bf\P-�xz@7"���#�F���Q�/��xI�2r^�$l[��I^��;���>�X^�p���_����+��f�Ҡ���Ȭ�$�ս!�+�:O�&PǼ��'�)��F�+V��r4�q5�o9���#r��P��2��(�*A��`�����7��z�'G�{
��a߬a��@5�n�[<�����r��`�F����-l��F�0�R��'7���(�[^8 ~&���i'�?0r�f<��GF�-`��1=�b�u�A��'��>dt��`w��v��Ҥ�n��!`�N;-��S��S#��{��kU�v.�	\��0���?��&�S��i�3�Y�'�s��ѧ4/�5/�Ok>�>��zY�yԊ�U��їX��5_A_�|}�����5�o�oj��������{����u��?i����_ѿi~�~��w����'����i~�.i.�ʹ���*���g���b�y�����m����9�?.;{�%��Y��=��"V_���6;�;̻,���5����-������}ϞO�|�������Z��l����Ȝ~/���1���wE���ح��?YH����A�@�G��I6����,j�+PK
    +Q�H�A���  �    org/bridj/SignalError.class  �      �      �W�oW��>��zI����z�tܖ�v��I��a�M'ԩ�4}0�;^�3;�����B	������B�B�JS4��!*����								���w�ή���ʺwΜ��ιw��߯��-������,��9U�r��B\'��BgَEI��u����eK���Y�(�*�[�תT�� �58��O�P,��^���붼��U�٠��(���U�����Y|
[3H`�+l���gч2HAfу�-�ݞ�Ѣ�؂��nb��üg6�B`s��KJFYT/9S����ڥQ����jZn�+��%�N�>J5��$ 7
	]�Vc����5���U����-�i_(ף+�Q�eP��,n�NE�غ�8�{�^��X�^���wd�Y|Nm4�� 7&��[��Ca7���/�ܒ�籟�v�'��[Q�Ј�Nݟ�A<@�z��*{7k�V�?�I�bJ a"���H4C���+l:IEQ�G����}}ob=��h�����_��WT�Y�����0=?4k�������j`NජǦ9�n5��p|�\���r[�N͜]��^�s�t����M�ҡ�>�k�3q����
����cg��)�g���g�w!f}q��-��k�I��Z#��Q��΂S6�2mu��g'��֫N�,pK�^0��e��3/Х�P�J~F�";��Yq���m�Vͧ��7����e��,���G`��ӷW5��t��qĺT��k��K��*m��ѻC\�rho�)���BW�R7� ��\��(N��&ׂ�7��&�+H�@~�b��jS�F��XeSj����*'�D��UK�m����Y��l��n�Y�G'׽�g��v�����"6�uv��ki}��̉����F1V����5c��U|�`��񸨲j��ۼN�9
쪚0�2#L��VƜ��������������x�0h�[@���ۓ�R�/��e)g|�6o�Ur�jc	3��l�V������Aٞf�0yZR��%ѯ>���'B?���s�9�O*@���X~x����Ʊ�e�������������>�=�/hJE�R1�RQ����y��b�a;Ƒ���ӊ�q�q>����G�q�*�bơ��͹���M�?�� ���P�8�1�}��Ƈ����N*Hv��w�N^��;$��"�p��R"9�.zS�!�\K�lYv`í��~��O���Q��a=JH�Q:K��;���׈�y{�`�
٢.�����+��B7.#J�c �����=|N%�k�w*�zr�h(�_ӹt.uok��8x�*T�/�in���s�����.=
S�H*ʈGgJL���r��92�I�u����)�OC}��,5c��'i}�3�E�W��}���{����N
}����)�sw��}��[�4tQ�n)�'�0���z/�_��.ם\������<���cz�<��6��4A#ď���u�[c��>[`�Y�|"�_�d�cZ��T.������Ї��z�kR�5x"��\��R$�Hz��G2�d��H���ӑ���u5�bzX~%�_��sq��u��A�W���گ� �j����#�B$_��K�|%��F�H��7�GwM,��F*�����Ń,1��q�8�u��n��������W�^ǳx��\��<���gj�/�x������7�O�������v�H��b?;�S1������x�GpQ��%q�O ~%*�HTq�y�PW��?PK
    +Q�H� 1�  �    org/bridj/SizeT.class  �      �      �S�NQ]�PJ�!\���-Ң�\
(�%��5�B��P�3q:%^��}�� <4����W�Ÿϙ���M�sv��k��/����O ��˲���ĳ�� c�:W�%��
N�tx�֌ Z�;Ў4��lz{�����^{�a�٨!M0�d6)���m]3r�.��,�J�u�[�����Cۢn��21��#9]�VЊr8�z���e�О�p�M��HZEA�p�! S2{}DR'EE;�"��
ŵF:�v��:�n4�!ʋ�Y��^�^���*��k�����U�c@8��|���$�?|������l��@X�F|��z�:v�r��9�P�nU�b�����T�)��x[g��e��uwqO�fI�n�0��r.�㔟#E�v=14gϲ�h���֎�T<;��Τe�����U�Dfh��J��چn���a�۞G�Ze��S���
i}��0����"�at@C�l:�B�*y��B�-:VA�7��F� ����!�>ɒ"[�������r]��Lh9��3&��yL)�%<3�{�Թ��!XGC��8��qHq����^�*;�!��\����	\�]�^��=���\�%��)� ��Yu��7j�k�����-�� ZE׷y7�6Wy�dk]�3�_�A{ޠ�;_�����s���7�]����
/b����i���)�2iN1"LE�!���3BTQ�<����PK
    +Q�H/�=��  �  #  org/bridj/SolidRanges$Builder.class  �      �      �T�SU�N.l��-�`S,���`C�\
M�@-5��m�,a���t�wǿ�/��}ҩN)�t�}�?�~g��&s�����;������� L��aǭ�K�Y�Mo8�Y���U�va�nZ�U �v�{zڢ �^�5ʞ� �m�RC`�H,]J����]3�4��VZ3k^V`�kVk��9v5;G%�2쪷C���׼uO@�ɰ����S�� '�5kڦ7'�'
*N�d!��l=8�����SQ�F���pV�ڠ��l�TG�d�S�۠��������7�"�W*��vEϭ��eӰ*KF��_y�cg����1���hD�"!}�#�dk~�T�7������@Og�Lѿ�L�@<���?��".u�=����)�D,Rݪ~��*>��(f���_սW�sW��r��y��!�F1�y���X�f�����VP��%�z�~���;{��+�.����0��b7����ٖ}��2�ǜf�u5T��U_�l<qtcȮ�o��������)�b_G6̪�{u�-:'4��[�5��eܖ�@�f��Z�n�p���Sw�Ʋ)/jζw�SS3j���!~�\ltI��]=tg�C�z�'��{���D�;����c�}$p���3{l�C�~�!���a�g|��7�۸��S�z��M`iңx�񌸈.������MdB���~��!��P���3O1{*�+2��L2��!��#�H��Hᷘj����f��|0�3VؔMt�Z��_�a2�q�h�zү�A3tI�a����7������T�O�4+�_�(�F?2��\�}����x�+���#����9hs�:�D,���E��8V�sÒ��$��b�9.YC������?�S��(<��m�Gdך�)���G����~LoQ\�L�
�0�r�`K�A��|�0>�)�2@�c8�7PK
    +Q�H%�n @  �    org/bridj/SolidRanges.class  �      @      mP]KA=��m�Zf�Ѓ�n��s�CB�HA�>ͺ��L�0���z���~@?*���Ѓ�{��8�2?�_� �p�P����f^?R2x��D�Ce�߹�(�=�31J,d)����t0��h�ͥ
���g�V�X4�"�2�.I%�I2%����Ln)�v����!�jl�(���c��RTml.�6C.�J�n��qM�(�^4�j���/������z�)����{i���Bw�c����� s	����"�gc��A�:���l��{���G:�Gx�,��] eƎ��f�O��.;%lQ��2\��.8�hf,R� PK
    +Q�H�8M  *    org/bridj/StringList.class  *            }S]O�`~޵]a�o�L� ~�0D�ʗ�~$�&B��bB7�Q2:�:��x㵉Lc"?�?��?E}�"�8���yO�s������/� ���Xӫ�*����[�=ǭ���B�Z�V�a����ʮ]eT<A� ��Vi��Z���b��:͜�ʷ��q�Z�e�Ǹ�\���a�e�u�U��t�x"!�]26����!-����bP`���a���hV-�~�x�C`"]0���0��F��Y�c]���^g0$$5���1����<��hG�S�Mb*�����G���$�S��@nK@NeS�\M�2�i�C��d�l���$��ܙ@�@s(' >*����8�/v[�N=Z΢��X�P*�~�\69�h)X�As���9�Ʀ�9V�ao�;Wt\{��W���Hb�����c�ac�M�\���;�7��orM�h�y0��_�d>a {������LJ����� %�e)��J���G�tE�;�.��due��ty�P����o�����.3� �?y�D.,ƙ�I�;�-���|)L��!�B��"'1ÿp�ª\�d%�4�Q*n�zy�f#*�q�_c��w�	)XXbL�*�&�h�2Dg��A�Dͱr�����fl��99�d�#�>ϯY_�^�S�PK
    +Q�H��ܭ  #     org/bridj/StructCustomizer.class  #            �VmSW~.�!
D�b�M�KC#V�K�A*m�*E���\��d7�K�~�Lg����3:���N�L�';���sw�l )b���w�{�y�s������ax�,��+�Fi57�ڞ�Nx�kU�o���^վ�r�,�W��ƱK��V�SJM���Oʚ-u͕��@WɫV�"}�ÅF�A�^�r2�_�5*9�2u϶���&�ӫ��2��h��CՑ��q�����#�i�c�2I$�7��	���${�rٲ�x�l˲��)p:��uR:�m��z��k�p������ pd[C�Ĳ!+�I�W}v���&�ښ�S�#�ފ/��(hk��RC��%�ë`ElV���J��߄�u�3*%���IRI�,Kw�t\�ԥ@.Ӵyۗ��H~Ŷ�jŊ�#��$��o��Y��q�@:�h���h%q�$p�ވ�f�!�8�<!["���^⌛���t�U��D���"+�B.�!�f���#�?3��.�3x��8ˤ��n���L����y��[I�z�3]�*��ӥ��q\8�3n�,�ۯ��H�� �Ҍ�,�]+�ےE��覭崮(�;�>�V�I��3Ԙ��列l�"�q\Vhq&wV�6�:I�
�Th
��<i�߭:�i�A�'oaѢ�Y�(��,&���u�l��
-J84���O"�U���<wzy��p.�`����K�to	��+l�-Y�z���눝oki�����4U��pԭ���p����D����6,$��D(�@{mǈ^�{{��ۧ�e1�3ʦ�z6$6a��J,]�,h��WC/����Ei����jk���t쨉����m���홦f�2��F���<[�S��7��Ma�pf#jP�b�c�#iCB�0g	՘!��K;)����5%9���٧�z�T8&!�}U>�}�0���������G<�'�0BC5ۏ^ߔ��44��������ů��-LL?m�aj�z����� sG��e!L��@�����x3`*����>x���u<C[a�|�M�c�gN>���_pN`v�9
C���05���J�g�/�6�_����S��>X�$����C6�8���qm7�cOq�w����P�6�)�����I�ﰋ�� {c$���3|N�����k�����`�SCgh*�P�*X��c�2��V�&����%Ò�̄7h1�.���Mfy���d��#_�-r��;��������z�+��!^�~&��� l���Yy����x�������K���}��l�Q;��wn7�7PK
    +Q�H�#��U  A  !  org/bridj/StructDescription.class  A      U      �WxT�>���f	a!�@"�$��T��%�@�\�����$7���q�.��J�֪m��X�H�Vl�B�ЂH��~[��a��b�}h[k�����Gv������;s�?��ϙs�x�~":A���G;�F���v+��ꉮ��o1�MBP�m����H���5z��&���<��,'���У�	Aǝ΅^�KY[Zyr�ݸH$�&�G��٧�� ��i�j	��g�S �;7;87�}��~`�%�{�p��W W֫%�i�l��*l�J&�X���s�5�
�r-������J]�2��a#aAjf���#Ǉ��%bQ��Lحw\������q�_7���X�Y��~� Wg҈vr�կ����R������&
�=�n��c���$t�O��x/M�)~*!C%��M>�wj��<����hTd��k��<���]��=�֟�lL���J+�����aFZ��8M�t��i&��oMCH�V�t��_�Ԣ�W�����~��fQ��>K�A�s�����t�=�͈���jz� w�a���P.�6�z�]*���5&Yk�M����-�P�Z���X܈�M�-�m��5WЩuy�S(/F�<si1s�Ia�'��������#?���S���Y~
���f�e6,�O�Mgã��ii��`VhqC댲��
��a_E�x��>/h|F�̤i}�)v�6��/r�u��w��^�(�1jm	u!j�c��æ��)
<ҩ��"9;SDq��;��R�
EmҌ�(���Z��[��ˤ�
*�b
����I1F��!n�y�q/�G���H�0�x.�*�Ƹ� rD�N׭�����s�9����"/]H�?s�i6ښ�t	
t! 7]&���f���,QL��m��%_�/y�r���l)l4(7�KH1�Ӟ}/����T�S���!R9�P ��Օ��5&��}-g�u𱾄�1$�J��o���X_���|X[K�\̮�
�2�@���f�6�-,��H���uEՎ����C7{�&��̈.��b7݆���;�?�A�=t;mAntK�N�O[9	�軸�'V PM���^��^���|@�H�f5)cPg��uc�r� �b,Up!���vR$��$�;�*H��i�%wr�Z�AK��x!
E�7,K�ҏ�${QfU��-Z݈|c#j�~ܔ	�D��<��=Έ��A.{��a4`�C葴ԉI�G@�I�ۣlԵl��PX�SOb��SBOC�<�2�YV�6���Y��]����H��c&��2ss2���^��1\��R���-��X�-��:-��9�~�ߨ���7%-x�!գI���ר�3��;x�4�TC��<����g��_�\�C������g�>�,�֧$��$��f�K�3w?�GI��C{I	}�g���X��H��n�;��aj;@5+Gj:[cݲ��ui�T�p��V�S_������L�P1��^8-�Z�O���E���;A}�4�օ��`Ȧ��p����X2ޥ/2�:MBmp��C�C #'w���ϱ�����"*�;�8�^N������5��\%~Qz�[N8:�F�J.�efp����%��79M�
W�sUL�p͘U\U<q�>��%�}r8ر��N�v���,J�;��࿎���Z
��)DҶ*����u�tj��ΤOCZ�k<���!�X+�5�h����NH[|0x��cL%��rZɨ,%er�j(9�� <
$�8 `�A�4�<�n�,O�g�����Ux�PG���7c��ʿ��C�4g���x^��V>�fW��҅�U8oB�ȓ�ZsihS+K7�L%��ۈ����}�]ғJ�2���Zo�
��ҽ�V��
%Գ�P��V��" �t<����4tyB0�|yB^H��'䣛�X[n>����t�-w-B���t��)�r��<����H'��S1���ݰ�CnyK$O;!��=�1�^|����@z-����e�$)�F1;-���b� �X�^�4x�,9TΣ��n:=8��p\��`h�v���]��a�����y�H��M���A�m���>��d�:dP�
8�z�JH9�T,�#NB��b�Z������8K0��#9/A�\�p�9v�J]��N�:��� ��(�������9��5�[h|�f�,g�3p� m|�\����ێ�i>���q0��8Y�+��̕0χ��-�˧�iR.J�+��M�}%v]����\��W�W�7�]u�i���*�]Y`�r�:�?^�*C�,?2���eV��m��g'�N� �c��:�\؉y�7�B�`o ,��3�j
v�T�I��+�Ѝ�@ݸ�~�s�|ݵ���2th��:� �!�3�#����3ۄ�,=nAN܊=�����݁�y�q'��]�˻�[��v��f�s�]ǧޛ�����+9z(� �9�� �d�~@?�Y��R�y�#�6�,�Ӧؾ�2)�3�v�(�A��n�&H��^d�*���#�L�M�S��`e��I��~�}d� v��J{l�����rf.gz�} �~i��R�	��vVq�!	gS�h ��Z���P� ػ28�8=u�~xXM�\M��)�=&'�`�?��9l����5[���ը��3
�9<����/��ʹ�^�+���ux�7�^���M�-��{3��A�ٶ���e�'{�5=�o�y6иP���{CV�G�V��������W�~d�~8d�c^�0�w���"���BcI�������#!P㜴X�E�:.e¡��Xke��N᲏rz�GQ[�U�8r�	�든�S(�O��y����{���(�/����[�%���A�Wh�
���|p����όRz]LE��'�[�_g���\:,z�h��W�� PK
    +Q�H�LxM�    &  org/bridj/StructFieldDeclaration.class        �      �Xi`\U�nfy���6i�Nס����t�4��0I+--M�^f^�W&3�7-�"e_��"LUT�fH��ť(��n.hq���M�&3i���;�l���{n�y�� N����U�a[���k;sVZf"�l��m8V*�AL�ll5�F��~u�f3�h��,,Q'��q3��B:f[����?m:�i̈�X���Mշ�Nw*N.�����	���L��,�[ ��Hd̦��NL9B�"Qp�X�Ҫ�$O�+��dWNֿ�JZ�rOE�zS
��4�eA��T�Z1�0��n�OG%�4K���at�n+}��G�~���&wRQy�^\*9�����X��ik��Irޤ�c
��u���b:_� ��f2.P[�Ϙo9g�*�Q#P�H�JSdY$�z�Y-G<M
.@ ����pf��E:��D�s:�^��Rc�t�y/�JE��� �O���������T�`OU�W�L�����t�0w=&����k�U�6��RǙXD3�"�U6&�)�p���	��L��V	����H&����@�9	O`aE��#c�֏HѣV�����٤����4ך�[��i�U��ұ�Jp.�c�qk�@@[��&ۃ�bUe���h�|l"{���Z�J��r�LHqψ+�Q
&���SN7�J�G�J}�#<g^&!�j�ZP���ml�����U5i�j�i^G��g�N����#�� .ERG#V�z���N��qya8*��cw6�R�#�ѱ6S�VYQ���1eG��(�-pF���Gp��6v9���Rg]Kbq������#N�e�*���;J�\�7��Y����i����4}�d$Y`Y�@�"�Ǐ�2�70�.{�M�NO�H�����ҷUGoA��t�������S�*b����n�#T�B���H_������8�.k�q��H��v"��ݙ�{�ď�x����v"��%c�f$��P�]k%���H���H�#N*���m��M#��1j3�j}��϶s]�%�E�$L#-%�wɤ��HK[����l���L�3�-���6e%�u��I��Hx�Y;�>�N�C���a��
�q7�(��~Y�@��v���j.t��m��lr��#S�LΗ���u�������&P�n97Cxe�a�c�br$��ߚ���¾j��9NsPM�@�%<*A���~�C�㣆�Q[�0�f�%n�����Tjr���`Y�e%���>��>|Ez��mV.{�(C��WqP�~J�Ų����<gG�;�t2vR*��M�E3���+ߒJ��m�R��n5�x��]��V����s�����������Ű�r=��6����?�j�۰��k��S�L��|�1�D#���%b�IES}���b�rMR�e��/�+�t���t~#��o��t�#��%�
u*r�����8z�Xa9<��H���7&���;��)oFQ���?��t�E�	Q�)�a���<������l��K�ޤ��5�]N���9��)��j��@����;2J��Zh������C���Q���Yi�.��DҴ<���)&T�=���ΐ#���0�|?Ӛ�@�:L^c�i�/О?������ù�pǆ*&��A1QLQ[V[�E���D��-�qlM�+ֵ�vs�.���a�q���s/b�������񓢝VB����l�L�����["[�8��z��|�*�\-^KN��/��)WW����u�#a��?<��V�l������fc��-��eJ�*�Ζ����kyv�̕V�D�M�������I�?�P�ɫ�z�'�7��O�[&�w�o)�K,)��m<�5s���Ԫ}(��� \530�}�}Lʊ
eCqӟ��'RPG�N��\��,��j���}8��O�ڃ�TeQ:�?����{��[|�=��ۏp�5��e�K�,�'E���p�Cg��G�8�����r:��s�6�@��X��wr�ќ��f����{?|�GHm	E�bM�V�{����A\p74/�<���
q!.R�o��s	M/dt�K:3�� K1�0g��6����B���1��G���/@Η���a��V����r�"o�w�.l�)�.h��}�Alى�o�Uؗ�e���t�'�߃�k��`��<�-���|�>���W��{qm6����w�=�h�������E�2_�wN�-�-h������a� n�:aRuXˉ�>jxn�}����2SY�"�vfeqg�.7e��oC��P=�3_��0�E�$T%�5l"�~|�o�h�̩sy	��Uہ�s9��~�_��|�o^�S��������[���%�v,V^\��K	�7>G ˒z����$�E��*��i��4��1%S{���6��,�z�+y�]�u�����z�i#���|)���_�"���݄���n��|	#� 6�%���+��n9w��Ѽ�A|9Z͢���������k�^=R!����n>}�a?���\EamF7��p��M�h6����t��3��,��6�n���i�
ڼ���k��`�qq�>Y߉V��'����@kM�Y�d'N�a�Ɵ�/��,^�Ѳ���V�f� �di���� ����k���|���s�7�kCo�>� 꽇0�:�݋�
\�֨�����V�:�T�<z+�B���+a�!���o/����+�ϥ���h�ʢj
.��D�@C0<��ĳH/��JvaZ8X��/�P(�`-��Yq����������g��z�}P�D�K�6B�qDrv`�Р��<7&�Mv��,��-�wY"%�f��q��lR2�^Mn:�?��V����Z;���"�vq�<A�c����D�UxF�'Ѻ��vZi^�C�+�k�k�'��ل}+�ߎ��F급�7s����w�q܉A��~ҳ�/�^�z�-�0�.w��|N�C��ô�/c�XŖ D�:}�PK
    +Q�H�y��  x   &  org/bridj/StructFieldDescription.class  x       �      �X|TՕ�ߙ�����@@p�tD���e�|I��%y	�������Z�c��Y��Z��%Z�E�LE���v�]��vխۺ+��жlw������ޛ�Lq~̻�s�9���9���ÿ>s�<q@ OvV�&#�;�[�d��Z1����T[2��"�B`�c�Q5b��M�;�6���ġg̑ctv&�N�2ەD��z�'mE������H`A��~�ڢFҐ�-ᴀ�tƺ̘% V[�XfSGGʴ��z3�im�dk�rr�ҋ�d�����i0R�pI�I�nI5��N�^����z]�'a6%�㑘e&��NӒ$����P%͎('UK}.�+(BD-R�k�M��*�R���!&4������Ō.
��0n�X�"��e��X��D��kJ������L-���֨I�|��X�Z"�W�� 4L�xv{TX��1=���� �W��#��$��Qd�f���Q���h�����|���:Fۣ�*k{���:2`�*}qg{�������~N.��v$Ɔ+��ϸ|��t$�n&��4�:�|e/�EWhq��h�H$�#7;<X�`c��E:V`��}��9t�cWIA�{TU(�h�@=�I��lEkti9r�:ƢT�t� 
��V�,��R��y��(?��WJ�6�X�K�h33��[�RI3��t�:<\*G�>w&�l�GmF�]J���3m�L3kF��$"��6�2&V]��6��T��L�BB�LWl�&:��©lh?":��� ��J��LӮ냊Ǆ���х����p�c�����Mf(�&B["Q���ٶH؏�rk�N"?�TI��?)?v3=hhY��@`ְ[����{�/�=�O`�1���E�4�bu��ee2�%�o���M:>��8��
��?ce��U��`i�(p^��F:j�����_�FLy�7A܂��[)��HFdx������ȸ��6<ݹ܉�p����-�܊�d�J�z-0#<T��Oc�pw_ėXJ����<Db����q���Jǽ��ݸ�h��פcV��\���t:�X��RX��*03�7S�X�
m7v����C�*�f�$�)*��Z�a�ڪ�=��!�X�����JsG<kEb��P���G<�p!�q.�e�|�&��1ˈ�R��V�a�-'���#2)����T�{ҮH&�<U��<UD��W�M�c˓�;4��AXe!,1�*\��~;l��q�9�ʟ��]�XBBg"��R��SN��g{m����*����)g�=�fI߂�M���L���)�Ξ�Y�W��Րu������S"��'�c�l��u�(7#��{Y<*m��&�W���,�.ذ��e��T\�Й���פ�������n�v#�h;��:�(�?�M�*����IU��[R� d��ǯl՗�]��/�^ o�_u��� ��ӞR=n���V3�����T�&���F�����ŻZ#1eD��M�&ꥪ����$�6e�6���X���������
ϛ[�N�]��N3��bN!�%0#��d�+"{v����-���}��{�ȕ��c���ࡖ�j����[VmZ���q<�3���ɶ��W-������3ێ�s��q��W��d�#������_�`c�uٛO��I�+V��+49����w�i�_�x�� ѕ/���/�=�L���\2���m�`��t1B�
]��5j�@n�qcĘ %�Y�>F�/�
���6���K��L��R1����3����=QG��H1i@��^��}E,����f9�d���T���_D_�����4j�$��t�X|W��P(��H��1��2��wU�J8I��,7�bN�I�stL�9r�\g��~1? Η���R����X�d}���ǜx���⢠X(.�Wi7�M�XD:�W붇�H�zi��C�]�V2Id�\���ES�eҹ��n��D��x23w�+��U��&Wbu�ܕѸ���{Ti��<����x�:/��u�T:��U�	�.�نF43̪n�;�/]~�����.������!PIFah�i�Aq��_F˶<ޕ��O�p+	ц�Mb��w�o�v�nu�7%�`X���j�E���� �ZU�V����ufc�u%$�-/�nO��!*�M)n��l^x�<^}Q�|{Q�~�a7��iu�r��e�x:A��}:b�GR��#�<;in��٦��-�|�(cm�$���W�eX�.Ҫ��4�y?��IFW[oWP�mF��2��:R����V��GQ��1�#�I;�O��t#�YK<�l3WF�&��0Ҹ9�,>ȏv�eJ��/�'��� �����<G:�Q�s��d�Q��9��Y�q
��;P�	�ɚ����<�	�/{k	��O!���x�,�<�i�����8fC�r,*���~̱s+�0�/��B{|ѓ*���W���b���}O�ҁ9�\.l����8X@����s��qh
�PT��(�k�zV}#I��^�3FB
*ޥ��B��(�(��Y�ُ:.ni��^|���{qyq�=�+�M�x�_a�p�G�K(,^׃rW���ҋM���/�[��ᑼH�9��)�
�c����<��2>���E+�Gk7
�ڻq����N�y�8���Q�y��>�5��k�̟Շh����ѻe�JBM�L�U�����]�>\ۋ�Qڏ���r_�v7��{P܏[2��K�#�wk7��6P㵍�{qg�V������ғ��l��u�,�Z�+�)o�T��ntC�4��*~X���q~.W��U�MW�[(��ŉ���_e��)<q/J��}x�E�8J-Ǟ+��]�]�%�+��8�H�#��,~���x��	���9��r����:I�\I|>Ǒ�f�Ƚ�s}x5C����Sx���m�.�GNn��)����@Tgfp�񒝸��#!.�_�+�;�����H�e*���,�,M���5\A��0�Z�5X�u�����F\�����Vz��Z��w�j�J��I?;���x�Qz��OIq9�D���!�M��^��E����Ð��a�	�����k=мK��"L�O=����	D"��I�[;%G�4�vMAy�Q�Ӌ��	�����:��u#!���Q��O�?nd!���p������yY�*}�#i�hU����ǲ\�<�O�X�z�w(j����vٌ��Z"
g�W�2�?8*��L�chɱ$�}b�QQ�4Q��^Q>�;��pΡK�E;&&�xΔ�P����TNtߘ�*����4n��q�fZH��4"U�Q��b�\B9�X"*d�������*��n�n�|�ݍ��UKe6o^6��x�*���%�����,p����e�9���9��e���zF�F�H�/�d=:��%������ucY��\1j�eYƧc�ø��c2�ȺCnȳ�?9��<x�_\��r��wz�zKĕN��F7��k���d�dS���9�]���������C8�.�+o�x��c��b��zqF�/=(ʺa�H-t��eN��Y���@v9���I�)�Y":%����H�|��߱b����n���hH�?��ʞ-{��{ޑ�}X(v���<Ymee�i�X�W�����&~��E�� �'P&�x���^1���vF��zF$T�V��V|�]��7E�'�7s>�R�v$jx& {���M�>L�~6Cע�'�z|��z��%�܄�����q3��I�c|���q_�p+U�&F�v^���*��q/F_[qHt�n��_������t�Wp��=�AO	�Ꙍ�<ux�ӌox��0����x��G=G�Mϳx��S<�yG<�Iχx���ޱ8Ꝋc����.�q�J�y���w��^�~�N|�{'����E<�}�����/2�/1�?�f�em>~�m�O���c�3�a�\{�k�xC{oj��/�W��>~�����tq-���4�wsodS��RA�~�p�����E�ډ7JY��\��	^O�A�~촢Ȏ�=�d��N`�.[�%�o��!<N��������f�Q��>��V��
�S����u��4���DN�9�oש�H��PK
    +Q�HLM�`�  9    org/bridj/StructIO.class  9      �      �Y	|T��?'�d�Ƀ�@�h�$+T�!BIB $�:I�dt�ę	�KѺ�WwT��խw�b���+��Tm]�mբui�����~���7����7w9���s�=w�����%�c�;���@�Ԧ���̩�@gs���I�4�L�Z�T���uj]ә�搓����L�n����9Ȕ�H�����.vw�f:��R�(b3�Y�ѩ��;<��b�=��;����'PS�4�2hi�cF�k//��O��)7�|�ގ��ߎa��PM{0�no�0M�O�� L��V�ѓ�t��4����ন��}�l���0e�p���1����`�vQ�dr)�d�Ж��F��Lǌ1P�&��r����1VX*<l�MMyt�cJ-��{Cs����r�&�D�?	�z��7�SC�m�c'e�)_�,`J��!p|�3���Y1@�UG'����~�7�~$�S����.r�qLc�i'�d=��3���	8i��X�bو����E��Zx�[L*�NpQ)��H�Au?ƶ�y�B{�"jS�����moň|+k�#FF�Utz}-�w��{�a�Ө�����0���ڋ]�0JN�Ebqq��8��ά��K�� ��5�����Ȕ�9���c��C^8z��br6��t��Ú_��ɴRb��mO����nb�d���y[�����ۂ(��Bg�԰:"ڨ�2��k:�z���Zh5��E�M=�$r?V|���+��D����4윀7��z|-�F�wȻv�$��s"���s�M>���\R�$&4:[�v)@j�;�W+��U��3�kc��<ᔘ���M�u�^&�˔w��N:xt�P2Ύ�'��OiC:]@"ڼ�y��{�F?��Ŷ�g��K]t��$��p��ED����N�/�C:���Y�����0[�FW�U.�9]m[�*���E���x °ت&��M�t݀��i}�S�zuPNC���&�,�ߌ� f���B7�1:;�� ��[�]��%B�����6���(f��I�ucn�;��(M�I�e���\�i�����mK�Q��]�%�܍3���g	ˌ�{�>�~���"O{k�M�+�tK��۷��LG������ր�'�k���ݡ�65��0?΂�	(�Eˎ��#�r���U�^��#�������7Ԭ��/����=��n�ըѓj�S��z���I�ge��U��~1><-w�:=���5p���"$2^w]"�%,�V�׭���Je���W\�2�
��%�^�<���72���=�]㙿��c��7�eNj��뀊��<O �����y�dg!�婬��:�_��]^�N���Rz;�nKX���ޕ�=T���HC*=����#����$��Y����I�F}�ޢ����*1���R���)9$�$i5���C�V�bz"�|���R+ʋ�숸pP�<n#�W��p6dޖ�>�O{(��7*�#�������b�ܿ�r�D�����7�UGa�������}� ���[�yexJ�&�h\��)	�ŚxJC���y�p���_;��ĩ�G,�:�^��;�Kw���ų����&�g]9���/ �8��B��!=�i�Ŏ)qeg��:��sOv򈨫���UwJ��l�;�T��#�:p��j<�ǈc�p�;Rg���~�1�G��b2�v:[=p�x٧r!��o�)�Y���8�e"��&���Y�҃�@�(�`\t��+��ir�
W;��	������*����e��HG��;���R8��ӱE��V�
��aT��L. ��fF]�\f+��}��O���8}%E�oI~M�W];���\����jA�g��%�ŖH4<^���4:H2x>W��`��#�k�&G�r��Q+z<�ꎜ�
�vmm���k���K���_���?��=5�7%�V���� �p�͉Y(2:5_���r^!�O���#�Y��w��éZw���-vς�x
�P��&��ސ�sh|�^�r�Ƨ����0��I�:��`���>"�FE��}��P���6�̳����v�Sj�YV�[��_�54��܉�C$j���]C8��!�6�����z�n����5���`�.��$-4h�3�X�^��Xo�����"�2e�{E|��
YP�P�[�z�b޾� ����V�^��W���F^F.�m�+�#��o�E6y�BnY�/�
�}A^��-,u)�R�N����G�T�!��6�����w�2��Jn���.��j1Q+	�j���{��}*�V�;Q�~���2'��W���w�Bہ�J�k���r �Zc��4���b��b���q�څU�Ԙa�aU|��e��Fۖ�ˁU�|�YI<X��S���}�H>R7F���H�������5,�er�%		�L~QM~IM�n���ʉ�*ˍ�;�W*�ב��P_��(���f+��5���n6�%����7�[��B�R�++���jگ��̨&'�����w�Z�y�"	����G��ܯ��.~�?�^��3~�Ɋ�l��l����/.>��zGU�u�7ԎJ�~#�7�}���ܓ�E~L��{�t�i�����l�0ԮFG�OR0$�M�����,�2g@7��}�v���`eb,��/x�"jYy�u��L�s���o2�
����V�J�q>��'��\�d�1�z[T0G�)h�Ϩiq!m�w���}GI�@]�Li��'1*U>9(�\��ʒ���\���������t�1��{i���֋����
��?�s��r�n �0p��j��r�Sx-�O��.r=B�h%-)�O��P��¢�t̒���UXT�K�+J���.s?��x8R��f��,*���<�6�r���񄅨����\����c�%�Q��K�hZO�1�����`o9>O�|vl��A����L+��m���\j�ZJ I���K�*�{
�&�D���v���م�iF�*]YT\�K�i��4o��eY%�*`��'Y��'Y/��0u��J����<7�o�Ԣ$�/1���V�CVCk{hI�.��Cˆ6็N��z�BbѺ��i�as�AZfaQq�����|m��C�t*��ʤ��d1���ɴ�0}bX��b���Z�22�1�G����0|xH�f�z謈�٪�4�L�+SA�Z9uSI���g�B��]t�VrlW��-.�;'y�c�#��_<�1�,%'e]��R��[/�"���V���,5'�I�b�I}���I�GW��5+�н�n�q[z��2�<ݱ�2#���.�~Q�S����I�0T�/���v���n!��缕��ǧ�Ш���6ʒ5��7��k���I�7V\����{譕� ��D��^�>� /��-aU�����v8�>�ϩà{5��b�L��B���	)�&lۿ"�� C/}�)��
}A�!P.�D_�^�G�oxr�g&����xRX><E�k�Qx=�χ� �����"$���:.��ˀ�r$����W ߕ@u�\M��5�M���t=�K7Ї��)�l7a��<������������WhtE�Ƶ6�S�54�q�ֈ�֩Ɯlձ����Aei]�a�C��'��4=��rҞ#-'M����+���V�1���0N�d�e� 8 ��ЁD�BJ �!Qm� �Z!�����y�z�Av8��Px��{�PxgE82�PȰ���4������`�FmC(܅P�8��{��>���Fz�n��������C���=@���G��v���N1���a��}�%%��D��/޶�v�G��������ӥ��<)怦I4nҏ�f�Z�\�'�@Iv�	:u�8����t�� =�'O:I�a��	�}$=�qO�4x������� l8z���h��2��񠇇���rǩ�&��&��bi;���L��r�8�-'��"Nȗl�a<�����6�&¶^�NM!8�����	�Q@'�@'�@'������H.P�I�a�
F�����_�1<� ��374:L�(r\��&�\^�	o��g�N������_c�b.1��ˋ���i( ����r��a��a���x�5]�rd���7ͦ�������o��8�a`��š������^��R��0�D�g�����x��@� ��J���8ņ�����=|bG}!����X�hDGҷ��ч�Jڏ�����3���6�3�S���$��e;z��R-ە��q}�+[��.ހ����0�%cVF`�#��^�#Zs�3�<���M�MҟēP=C������2Z��g`;o&��)��S�����'80?Ŋ��?CQ����p��t��Q�=Bi�E��|�(�}�V��7+�'����z��xr/�ͭ]�e��UK���`:�`��`�� ���-4T�\ϫ2�+�~�;�7ș߂Lq���U�N#�,<(P�YR7t�8��K�K�pi	<ـ���6F
c9&�g���4DͰ8����p����T��Y|&�e8��4]���)�٧�)�
�j&\�@�x�Y$��q=|v��������zd�T}�����Ӹ������A����#TY%�����Ԯ��RG��"�6����W���D_e��2�/3����ϰ�wa�h4�Qg�L��sx]�{`��|���{ 'p�� �pyDˁ�E�j�XXo��6Em�Kc6�&�.� MT�1]�1]�1U�k�0��>�������"ΣY<.\Ɨ��X��̢���5�y��L��,35X�W�T�h0	C�PdTp-�B8p_�8�)p]���(p�]} X���L]�+mC�)4��b�}0l�B}����*Yx�[�i�<T��DD��V��� 9
��$�U8� \�Ċ��:{[l��E9��@p��&�����T��JpP]|w8��c���#��.�jp����&��-���JA�8vZ8H� X���R ��[8HM��#�;F9:v�8���`<�{���8ԙ V��S���@����O<{�{X�Ng��f xάK����>6'��Vp��@p��+��+Jv<r#����X����m��E_Lো}X�~{�����~x��������׎�� <a���������a���'��u�x=<>��w>0u���{��������5�χ�PLӍ�'舉2��������4V��~I���%S��PK
    +Q�H�Ǳ�  �    org/bridj/StructObject.class  �      �      �T]SW~N�aM��|)"�(-���ۖ�X�AL����7�d��	�t�a�{�Do{ә�t��aJ������'m��YH /rr��x��}�{�������sܺQqem�(yn��+�V��!�
�'w�}_X�|w�ܦ�c
\X�$��m<kٞܲ���ѲF�"�:�t����"}Җ^N �H��8�x�h���ؓ���ԙĚf4L�n�Y��׻,A\�L���7����",�u����g�����7_y
4�:�AH&�t?u��Yn�XJ�eBn[�+0כ��>�9��!�xm��<��fi#�d������:����fZ�jV]Y�f��鞕l�8>�L� ��9M�+n�H����&�+�'�G�(B��N��9�L����]��o{ұ)�:nDa���	�:ns"7�V���z�_�a仸�|&p�C�:�)�6��ҡ~�[�Qd��0xԫ�KJ��k�JM��Wq<�R�X�U�zV��>Ǖ�\�#�����Nj�)��o|�]�qu��?N�bx�'W?��~�#�a����"�hKNͯߩ����J�Ұ���s�&m��ڪXn`;�v{?4Z�u��Z.��}.�I�W"VrZn�Z�
<x�ʲ)I�hێg�ʚ�'R��ZԀr�/-��u��BYS{8�+7!|�5�6��_�/F0�d�p> (!��˳{�@��� B�F1��글�>��q\"@�`<xE0�oE�N�'Hg�0��>������#��S��ۃJ��c�:D9��_�Kz��ZP�qВߑ�儖��G�k
� �'�P�]����.>�y���F��0��n�G�#�����GT��?��ď���'�L�����9�!�	Er�&�Sܣ�,f�5��AL�w�]
��S�3(x��@�8E$�op��!��y"�1�-���*N�PK
    +Q�H4��L  d    org/bridj/StructUtils$1.class  d      L      �T]SG==�2�뀈��p%Fv]0�|,YŬ��Zeކ�65;C��R����ʻ/��ʂ�X��9?!?���ޭea!<t��ۧo�s�������s��8٨�'*ج�eI�Ϟg*L��9�Ʀ��UC/ڨ>Yߔ~Vk{ZU��斗xY��7�F�+��j����BM`�h4����":$�����x,]�3q��\�
�/�0m�4�U^�8W`p^E*[(k�0��È���R<:ާ��Jp|CQ
�/�.�tDeU�t��9rG@<t�!��%����T��z)ɟ�)�q�\|�O4�S��G6��f�.��ڈ��P֓�ɚ���T~r1�ϊ��������L5�ʎ/��l��������Z*dy����d��=ʠ��%S��Ϧr�<�Y"okKF���^"�H�J���R�ㆎ_e1��'� �e���n�}qr-�h_2v�5����\|����oX���ö�gq�S�ϟ��`A��-~�dӧ�ELbI����G�Asi�Mv�8Y>�)�z*�..�bؗ���a���!{9Lb�_�u�<����"���\�I�SX�����)�ŭėue�+��)U>�٫�\��(���:�b�dr���k��ϕ_�iU�
���}�����'�ݶ�8���A�Ù�:���M�=��pȥ+�_^c��op�7��+��7��]�.uy��F����t���}�ɗ�Py���љ=�r��[|Kkt�����c��.�)� �[m�Êọ:-E���q��Z&��|��E�`	׈�E�m<��UZ��E�|���=��MM����=<��^_jov�⁆�~�hY�h�Gsr O͚�W�d���V�8����PK
    +Q�H����B  +    org/bridj/StructUtils.class  +      B      �Z|S����Ҥ7��m�%��By(%P*�-kAW�X��@�K۴�IMR:�(������T�΁C��Nqdn:�S�^�m�9�:����w�M�4���_?M�=�w~�����O�,�h&O4�V����X��u5'�O��q��i����@E8i�Xִ>؜�(�i`3�itNSfi��tb�a4jY|����]�pK0��3���F:�f�1��EB�3��ʦ�2��
u�S�=������\�0��P[dE�� ��lɒiK�����6A:���;�E�`�hK������>O�L[��&�=���p

E#`�A�մ����w::�@"�����N�RH�jў=���,�g�Â�k΀�#�e�u����M�鱘S^��5J5�P��hWSj�2m�AS�L'Mc*J14�K4��d(e�8 �F9�t��`*N�87H�Fc͂�C��P�k��/n�F�u:�NW�TΞJ��27�8��ώӤd�v(�s����Y2@��`�-ў��&�}�[��܅ͧ3\TK�
�T�{�4SZ�ͺH"�&~��+���h�M�%.:G�R+��7-uQÐ+�7'�۹.:OJ҈����	���E+�4����h8�h��E��[�@l��֪[i���"
cc�%�F���B��xV@e�b��>+Nq!�Wԭ]���L-.��`��)4�G�]��4ز�3h:��M��NYhԆXN�H"��f��N�%����K0I��°h��3ia*O��y�fZ֖��ƠEg'\�-�ht(�Ͼ��ED�Nqi$�(�ts0ᤍ��DԄ6h� ���C-ɑJa���N��4��gY+Ӹt�X�U2K�8_��gI���i�y���BLӇǐ�]E_��J���;4�$��5�k�	�m�d�"�D ������@�z�A���F�MK0ތz�w�c!��p3��/BO��m`��'ii�e�A���n�;�8R���%�BG��HB�ɘ�$�k�O�Y�o .)�b��[���
�� :x��|9ـ@��0�k��n�B����]��5L�l� �Nz�Enڅ3�!�>l�}�n�"9&^��L��%9��~"��F����/j��5w �8�����a��q<'��}H�NS
$謅*�Y�.�z��%9XT�(-�O�`���M7���W�S>�#wdd���%Uk�d�q\�:����CR{���K/C��6��]N�.S�'q��3��JqŹ���u��� ������G�cs��4�h�������#�|8(�~l������T�Ԗ��eoM��2�'��N/�O�ͩN	���7%<�_�ׄ��eT� �~��ćO��VN~I������ԣF�a:�l����Jq�����<�Io�����#r@,�4�YCa���zO��?�;:�?)�9����/��_3JBz����u�MO9]�}I�������	���P*�ev��F��>+��hް]MР�H��å3����VS��<��-Nv ��@�k�C����&���>G�IBhĤO�i�M ��4�8 ��elM���`Vsa6��a��T u+��J;b�G��EC��$�gʽƙNÄ	j,⮱	|5�T�5�l���G�C`0���<�bc��ǣ$X�N���`t|kh�j_c��p[�leti �ܞ�~�e�CΜ+ҬĔL�B����^�'���:��ve�B��x�\�\���ǜXy�jKW��[��l3����\�s9�S�C����sZ>�Off#ot&��&�Τv����䓞�}���D�nW"hzQ}`s�ʟ�]��}+�pAW<� v#����¼��d�����8��c��Ø����\�2Z<��\�g䣱(M���I�c�h
b�ֶ�łm�:�)� w�n`~?G�:�O�v�4�!ز8o_�ԸA�e20f���<�,A5�#͕��Vg�C������|$��s�W#|��঄�kh��/�Rd�1t�Hn�s�#i	n2���uA��Ʀ��wE��`j4��sz����`��}�
��F�p��"Ьu�d$Л�@P���"���+T�C�v�כT7dJ�s!���(Az�<*
���T╁��lI��2�B�#k�#�dj�ꓣ�H�ut�� 7�����͗J�-I�ת0S����[��y�Bs��^.�\��!��--Cf��E$�/���[3^~"���IC�k�W�u,'�=lH��� hE������p��^���&7o�Q0���_�Q��(!��d8w�]0���E�;ૹ 4���_��.�{��$`�m0-{�J���6+v?��|߫��&�x�L�3;��6���L��M�j��fV�	�wc�)�ZgO�1_�H�K� if�H^{X2{+��1	}M'��ވ@������u�@���������>����~�eS(�<�3w ư�4�`���������AV��>���bd(���)i�n�CPQ"�"}
�Mf3�[�mA�����?l�h���|�&�* ���ru�9�~��/��q�A��H��^�!<�n0+����oh�Г�6���PS�,�1}_�}��[�̺��bm�X%ݳc�.$GWk�$8h�~>��'��$�8����3����n�/o�E�E�,�H;L��^^����4ě������� &����	5�c�M�pfR����͝�.~K<�M����
�]���o����O�r��4����E6�1f4�5�-Z�v�1�uP�ߧQ:���0c�l��y�C�Jp������j�'�]=G���̠:g��n�w�������Nh��͜��8m0*W&�h �x�s�U�o4wut�Ug�Ƅ}A�E�f��@x�A�2�~\(B�l��h
Ƭo&J�u���>�蒷mUCS9.���xLV��P�y��y4m�'uL�����/��+�]��࢐o�E"��"�S)�Ȯ~�(P��67V���?@#��f3�i��4���%W��N99���!���{\���>�/����w�>��k��ge)�t=�U����X�Z!. %d�$?Ҝ�� }*ȟ��d1& F���0c���� �막�z^�(4�3v&[�ȫ0�y���V�8
'������{�������G�젒~�즂~���FQ��	{�z�	4��P"M�3��i��l�E�P!_�Vщt���H�0��,���+��>D����4{��v���$�F�$��i�F�H1�,�E&.�%�t��x�I�n9����s���]�?��y�x<�|\�G;W���[�����ӵ��:�Ҩ -���GMݤ����}�AZkn(�裋qԅ��K��G��-O�zg��;Ӥn��>OP5�	���
�Lj�jl;-���zZCQZG�عO1|�)���P]I�X�+��.�+,��L$f���_;]�S8��n�O���]{p�#������\>���X���^��gW��}�e�/��H�@��j{�ar��ϐ���r����ځ�G���*5���J�G�8�r�ãUT�|���.��|v����G+<���`���{1��.����_�.:���n��I{���h%=���΢}X9�_z�����P/V�Vh�t�O�Py��beG���_pv�<�U���w~`~��Jw3I���� 5]� ��o��t#8�	<��[`�(L���'蛦^mh�Яf9_C9t�-���c��j���d�#�2ߓ�q<@?��=��Vk�Ňq�����y���G}��I�>z���C���:\��j���4��#&���}�>z���o�ѻ@��V�P�@����#�ZPS+����{�4��<D���ծr���CaHp D/W7�S��Gu�O�}L�%l|����|Xُ�|��8�-������b�����ѩW�.z.�Nak�U*a��XU�w����3w!A���ugp�Dz�Gb�/��b�-�(n��t�0���Q/���q[���N��'�ht��{�υ�vz a� L�P�#���N�_������_ңt.�6��|�~��5E�CV`_l�*�3�Ag{�O�E������x�^X�����8���OL.&��D,�)�U<I">���s��B��8�v�d�b��;1O�rxC��@�a�^���~���'l{pKE��s�Mt��7��N�-���ǧ�Dn}�Y���;��l�g�+�'�U�4���U��O)yF�:������T�������Z� �9d���/""_��e��W`��`�����kJo��ȶ������~^�tF?�=�?����ek�3ݎ�� �c8�Y]�t�k�>�~nrm��N>�-ɢR­�8j7CV�
�����k���V�D�\��?ȑ5��؛��]xS�Q5���@ey�����s�-���5ծ�*�V�\>� _c��=ǚD����7�m�v�$�B������z/�f!�v��L��t�n�6CVJ���n�����/K9����Lb/�}�>~`��z���U�aw��~�\X�v��B��Wtzd%t������ϰ �����_4Y]�+��{�q_�~�E�T+��ESX`B��bK��{��\��>�Wh
�s�
��I?D|z�Q��y�jxz��c��;��s��w{��Oi�{��92�ωQ���Rm�Kh4/����x+U���Ǫ�N���hmCF�	�m��#�e��x*�"�9����+�s�Gt�:�y'��U��p[�[���u�����u��AzT�9ō�_H�N���g!���_f�����/L/r3��_!����������7�ҹ�~�GɭJ�b�WS���&Ǔ��Ia� �_���˿N��JW�-ѯ���Q4"�C��{h�Mз�.�=�	��?#Ӿ���W�������}@�������d�7���:ƕl�yl���%��+�ɍ���P3�E���ૈ�~Z{���(��w؃)x�����F��V�cm'�8�l>���=fk[(���o��v���n�ܛ*�ެ���K���E�n�ԐC�馱��:�j��k�ۺdUeϫtN�����o������������*���d�)'f�-����>ry���LL؏jK���֪���4��!��<��ρ�s�vy%:w���j}��-ѥ{$p�>�k�8�"���w0b͓F�a�K{my~�y&�p��i�ͮ:�]����� �Uʁu:��V��&�'�藘l<A�)��4+/�a/�mN��VGxK��u�M�>0գ+�V�{=�x��$��Le|\�d���i�'�x��Lj�
��,�§��ٴ�OG�͡�Py�����h/�IO��;\K��z����l:ʋ�-�������G���v�_Υ����G��#+rؼ�+����9I�ыA��PK
    +Q�H�c(��  �    org/bridj/TimeT$timeval.class  �      �      ���R�P�����`��!"X�V��7,"��):�i�`�H�r�o3:��/| �ħpܓ��;��ɞ=����??~�A�aв�3%�Wv2��o$]Z�4Cc8�\w�Z�]+��eWB�A�§w�=�G��i6��U�9�U�t�!Y8%��Q���$t2H�P���!�D���c��ܝgO��
��A/C�}����$�.i[w��;��oG/[f�Q0�!\����3(Un��P�`T�]b�4l��F�rD)UM
C�[}��%�kYW��$�U��u_�u�n��+X��f�l!�יUSy)�eL�̧ڴ��9�=��=�FF�o10jZW�%[I}��N��S�/�D�4v]�\5���M=}�Y�$�v�)�1jժP����T�=�o�P��_霐�D��U��H��f5�k%C��t���j�Z��g�U�ڊ���X4M��\n�4,�U���2��j���34���S��7d1_Z��+C�����#�^BxN��;q}dW���<���c�qx���O�1ԇ����g� ���`^�J�OQsa�+���Z:\�� An!���E��W1�!��%�.�B�cṳ�4�"�@�P�6��t~�K%�^�}Ӛ�wH�_�%)bi���;�cM|������C��� RGv���
|�!�=��u���:��`�'D~ k����S�=�����lsx�M���T�.U���D�l��ɔ��dϑ= j�ʈ�PK
    +Q�Hڞ^�r  �  (  org/bridj/TimeT$timeval_customizer.class  �      r      �RMOA}�,�"_�(�Y�Uď%Đ`&h�/�w���ΐ��bL�op���D"z0��Q��YX�I������W5��׷� JXb#�X���]�Ț�Lh�����J�5�'���	nCG��WN������6���M��1��gfh[���������,r9����EoI�0a_���`Uū06���f����r�DrG�0(�Fe1��/�R���&C��X�H�'��?�6ݸ���+>�nG�-\F_z��0�\lU
�=U1�A�������2�����J����U\�a#�R-.<�ZY�������̫u-lxz��=�0��Ya��N�ܗ^P��0�Hߢ�$�a�cb��	�k�&-���-��hn��l��gN�L	'\��i/&"�+�+h�v�p�G�W}Q1��Ζ�X�kUE���;���̈́�8"��_��O�}�m�q�Ui�YkA ��+%Ɛ�7O
̬<��*���l���S��K�jщ.:�mK"1�n��\��tBZ�M�@
?0�~����bl��>�`�#r���+>c� ��P:)4� 8*d��R%�V�B��m�!��?�Ln�rF�0I��� �P�o��;ʿ�����>L�V��4���A;��PK
    +Q�H�C��      org/bridj/TimeT.class        �      �TsU�n�t�p)%��Xu�Ҧ<D��SE�-j�$���.nn�7����3� ~�9۝��V�tz����w^���/ ��
���f��ۍ�b�n��!p����ڷ��j��-���@6P�ܵ�Z�"W4�O-g��ik�e��|��8.0�/�2F�!���6�DI`p�vm=G�YίK�TI�w�����@�X:����ZUȽ���/IH�� �7�[{K�����_��m;Eƈd�0b���eۋY\����ڶ��.H�TI�%��WSi��0���]���۸�Ly��x�i�U�o�M�!�±�fq%��(�б�wi2�u*�"�Q�A8f����X7�L֓'�mL�q��ː~Z�}�b��sy�K�6+��\�)\�H�Û��\��ZmW������)�i�i,J\�4V�����5����i���T�u,����Q�6%���UW�O��ĵN4�N�Q���G�]�x����!�Ѷ�Y���"Q����N�;���$���'�A�ڮ�G��~E�L�	�"ן����=�e`����-oU�x�$,��oQ;��t�P[Ӿj�m�|�m�$���ꖳn��E�U� �U�U�;���C$[�:~]���!K���E�j�U�~v6 0ʫG�I�i���k�����3�إ�u�	E��D�G6�I�o7��6�	�&�t'�c��&���L�.Fn�I��"F�.l� E3�[�C�8f���9nG��Cb�b��� ��WB���h�Ѕ���}����/�I��?�R2j�����.>�d���Ͳ���.rK$w��7c	���yKB�bX�T��R�©��8�ބ�wH;�ia��{}�x��c-�t���� ��A�_���|�˱�i����Y���Q;j�7�
�F����1�;ς�b��`&�n�����	�Shѝ#ɠ�4��ޜ@�oPK
    +Q�H7C|Z|      org/bridj/TypedPointer.class        |      �W	{U=Sڦ�-�@Y�H�
�Z[D۔jC�hjU1m�6�$5�"��/����
AT�p�����I�yɗ��W&�w�9��3/�n��}����K�7j�GG{w��c�h{�i�Kǜ��=�A#>!k��ꉸ�#�a����j��	�P<ۭaF�+���ܫk�k(]�Fk5���)]=�������r$����ni�q4j��1��}:tTU��T���fw�}���H,3��i��Q�!�!�hA���mQ$z0W��!#qv%j&��C�,_��Y�|�[�yX }�S�",��	���x��Jy�T�4M��u,���`��rT�������զ�tǢCf[�g�v�F|��]
E�s�����ծrY���.s�	v�D5	j����fu�M�� �c���h�˴ʝ��v�=5�ѴT�{���p�d�i�HgY�3@�ב�TP��7�e_�+H��&2�����n\%��J:b���F��q�$]��<�d�e��J��6&��b;ԅ����P���f����ي�MCet��L��:�藜egs,��.�!�M�B;�U#���IV3����@DĘ�i��3et�aJJ����b�dd'n��.��l0E�%��6A�N�r�g9���;q� �5��Nd=�v��>I���()�FF�Cy�֘	��vu�G���v[����� <�����Cñx���x�I����r,����$�������RW}�	�u����a��r ��[�x��R^N�2�B{�I�������Cy��#��L���ࠠ�
J��H>����	�C��f�ץ�3���<���=N�s	�$�̂R\���J@��f:l^_��o��~�/�tNk���\E����x�[�8�����@x�/�����ۯ��E��N`Zw$jl��oĝ�y��Y�J�T���XE(60:#£wE�F<06M��B�O�r4��q�ϟxW�J�x�9���\��U��fb*�r-��G�6��Z�O�13��,�*�F-y��^wVj��ݯ���h�4�pj�ƈ�9�J�6��r�	�-H⼣V���Z��T�r,b���M(�j�n���6�I�Z���GF�1�ӝش�)�j4XΤ��J�Sh���b��̾.qz���M�o��u,*�y��%�x$Ձm�'U�Cj�Ν���֊ߢlr(�r������)�)I��4�j�H(E[���$�EV�Jjn�TURu3��Zr�_��շ�Q���U�!�)��|A���y�dm��T�R�J&������Z�O�3Mco��&̙�m��$��Z��e!G�T_Ev��I����zW_��T��O�NP)�R�\����Ǩ�?%�C�?�Il.ԟ-.8f��Z��M����ꋣ�ʟ�C��s�b��i����ͽ�$1Z�?;\�p�s�EIܒߟ��8�������݅}�88*�_w��^�?-U߯{������O�?L�N�
)��J�(ԟ}.8֪�y&�?�\}q�U���d�ᜬ����ᴬ��B�����ʟw�����gn�?��?�����4����~?/L�p��Ժ��P�����������INv��/������ÿ����B�iv��?,T�����4��:��[~,�/����J�'`��[��PK
    +Q�HB���   �     org/bridj/ValuedEnum.class  �       �       e��
�@���̴���.I�OA����(���>\����V;u�>��y<ow k�	�J�N$�$w.��<	Jy5A��l�9k�S�2uZ��w�/z�r����\���o�0��M�����>a�9b�*�i	A_,+�Ғ�R(b��1�eWI����~��4��c���PK
    +Q�H%0  �    org/bridj/Version.class  �      0      eP�J�@=c��Ծ|�w*��U�C�Ś�f&�P��	�i�˕���ěXPp1g�9���~~� ��C#�gf����d�P�.�1��b%�P�9�r���c0֖v�e�>X�������C��9�M�$VzvI�N�{�]k���2�G��G����m�?��#˾�n���w�N[T_)��k��ɩg���
�1�g�`h��O#�v��Љ'¥$�Me�^4�'b%�P�S`�����%��Z��hOdO��N�A�@x�"�2hel�x�7�b�z�;��
go��f�]B�GDM���3�p?s�PK
    +Q�H�7���  *  &  org/bridj/WinExceptionsConstants.class  *      �      ��kWE�g	P��P,��V�m��z�����$�lv��I ���4�&5�Z��x�}���9���V����l��x|�l~��wf��L����?c��C��5[�k�����J���W�k�ƶ�O��hob��&�*�+�Jcs�[۪�����N��%6�Q�se�9��U!f��3�l���#�+L׆����Y4�a��u��n�g��v�7����\V���K���������m5<�I]O��A�mɃ�pM�#?�,�j�A�O��b+�1��jZꝨ$<�츶����E��(�];�l���d_`�D�����+3�L-B��Miʲϣ�MG�������,����L'�|�[�З;��DI�<ʖ��<��}��UӒQ�â#���Ԧ���cw����N�e^�9�[Q�o���5���YK�ZV��6� r��ߧ��/���f��p �g�p�G$�ʠh��w&�)�}@4~H��4ԅ���1�E�{��-s�`'�����#)7��q"�A��<l��vݸO̬�I#A9��G?%��P�"ns���*f��}vsA���Ĩ,�����=��ъ)dt5��e���V@�{��Z �����F�1�D�Mu`+ ��6�7ί�=�pݚ.|t�f�J>�[WP�K�G�s&~����/�}�L�#�5q�+�� �I��nA��L�>I�K���e6��!I(�����`Mk�d��i�wD�]����q�8h����|\T}ET�/(�j��e��ܵQ�(R#�x��C�kq������p����^����4�yUs�>9au���Ω?ٓ$-�8�n�dG�*z��2�e'J�A:�Ɠ0(Q?��l"�Y���R���a<-�H��[�_�p���I��Yk�ڷp�]�Tcm�3��}\��;�mF���{���{P��w�x�jn�1�4�+�R�U��իR}asN�Quw�U[��h��i�Ws�z�ͱ,�X�Ͱa�?&�c� &<
~�����q��c�'��>�"|<M�$x��,����3�ς��?F�<�q�O��	_ ?I�"����?~�����k��?G�y��_�D�e�+���o�	~��-�k��&a�_���s��%-�B���Z�,k�w�����Z�=-�>�7��,��������h�Y��S��s[�ϛZ~���󶖟w��D��W��׵�m���#�	��左�w����:���&���-�����i��'������9t�7���ɧ����#<?�g�32���;��PK
    +Q�HN�.?  �	    org/bridj/WindowsError.class  �	      ?      }U[WW����b4Q�`�DQ�XA��c�@A�J���&3qr؛���[����R�\��۵���j}���>'1!
kf6�r�}�����x�8�aZv�w�6ҋ�ӆ���Q۶lC�fK��X�S3����G�%��%e�9��h����.=��y���<c��8GB86:�5Ű5e��E���]�P�.e���z�����af}x[�h�6�*���kʇ-��E�>8���N��H)胷,��ĂA��7�|��-lk9���>	���[(�U���Ilԝ/�4��u24��y���~`����5ai6��ڼm�4��S)�2�\��Os� uN�繙f8Ҩ	��*�Ծ0�$h7�CX���lc�F������l�U�2�7�=����>��u�,ۆ�Rؤ��u|���Z��,�y�3�Ă.4�]��/D�ڒae������;Ĵ!7vԒ��3�.�a���&'cc���H$:11;�K�6@x�|�M�.C��K�&�/Fg���c���<�Vǜ�J��e&�=B7E���j�D�z��#�#Ϧ����j��,O�^e��^B̋��#U��q�_tbB�qrW0F\���U�֍�saB2Z�(Lba�[u݇�0��$��@�w���ulP�Q�3�.�o�r�c��I����M�$�dm;�<�Z"̈́�pp}6cs�Tr�+*RHKPJ�m�bJ���g12X�ҙ�r�5Sm1��{������H?�������I��4�M�6��qn��8[�Ѱ}=U���"e٥u��L7r���c^��mSRPuۦ�ڜ8��&�4�fop-�cD-l�J��)�6�~R���q��bn���w�*�)>bd94�(-�/��rے�*w��z�WZiy��K�y9���ݮ[���)vt��"Э�bWw�em���	_ѻ[Ew �v@I�)I�4)I���A8�}���~8A�'��Q� F'H�-��4���{��jT�L�\��$S��iV0N�9E6Z�cW�&�����_edV5����q�7=���?�o��pX{�^��p��+�ۍէjj���?���|P��v��R��:3�8K�!�c&"d����ط��%���� ���/�"�_B��īd�(�}��0�!���?Z��G��E����p���|�#��p��KH��K��#�򏛿c����Y	�/q���~O����䞋=����p8^!f	)T��-�K�%:��RI���OxH����-��&5�{����Q�#|L���	>�үa>#�70��$���"?��1kU��U����+}t:h�w`����1�IR�UB��u�t�!���:�k5T�PK
    +Q�H���-   �    org/bridj/ann/Alignment.class  �             ���N�0��K[B�b@T,D���HE���X��p��	J�J}5��B\�%�����쳿>� �qB8-�ԋK��y*Ͻ;��|��uA�A�V�3*O�y�q"��b�����B������n�8a8m�B���%tV�TL�}*�N�"���c�|�y��2e+���}�p=b�����I�O�	;3?z����B﹨ʄ'��lga%3,�U/ulx������o�M�b ��诺8�u(�+�.��=����q�~]PK
    +Q�H�<�i
  �    org/bridj/ann/Array.class  �      
      ���N�0��mSB�_�,�D3S$RQ��*�NN�"WnR�I���C!�;�%��g���{�������^nR/6�c�,�|cD�ݹXO�,�&�\&��&�b{�������.Z��&��J	��ZK(�Yz ��B����G:͵J*6���K4��zK$L*V^��Z.83��Ҿ?�G��8��&���	B�ss;{�^��$r�47z���B�����܎��p�Y���p��8�T=^��vYӖ�`�ghJ�Ж#[��PK
    +Q�Hc��   �    org/bridj/ann/Bits.class  �      �       ���N�0��M[B�_)�b�`�bf��H-E!�09���	J�J}5��B\3�%˽��s�����'�+Fe����o��E!n��}a�˕F�X$�J���t����J��B������\:%a<kuDʪ��5����Q��?����t�?z~��y@8i�Ĳʔe�Y�`Ԓk��w��O�`vGؚ����s~OeS�j��v5<�R��Z'Fm�']��/J]�C&���ǈ�i�5}�v������]8�PK
    +Q�H�V�  �    org/bridj/ann/CLong.class  �            �PMK�@}�c�W�^DD�P�b��)h��Ԗ�xڤKذ͖�ҿ����'=X��{x�v��ۙ����p���6��9)}^U�}���c�|�}ū�e�ȭ��b�%���J]��/��2tV.7���,��B��;7�)q�po4L�)�����W�u�SQ�t9k��h���0}i��$�K�0\nvH�%b���G2�J�Kz��S:��곮M."�h�Ӥ&�T�ʹ��ֿ2�3���i�x�z��`�b��78��k`��6y�.�~ PK
    +Q�H���  �    org/bridj/ann/Constructor.class  �            ��MO�@�ߡ`� ?��ы�gO0�5�x�ԑ�,]�nI�k��(uz$�a�������ϯ� 78%�L:�i�:�T�x]�d6�#kRDh��JyZ%3ϟ�9�.���V c��M���JA�Ժ. B�q+��P���J�	��OF��Z 7�����O8ێ�*�����|_�Bj��%�ig�����G�0�tC? 8�W�[��yg��T�-�66y�}�e�V�ˈ~��x�yc�:�ʐ.��T&Tѐ�H"g��$�E���Dζ�]IW5ԱW���8(��PK
    +Q�H����    $  org/bridj/ann/Convention$Style.class        �      ��kOA���ew�n/V�&"hB�#�`�BBl��ؤ�Ӷ�uɲM�[�O�D�F�g����F���M��3sΙ���|�����F�n#Ws�ã��8�R�91�j:����6e0���qb�l�i䶝�q�����f�!�##��9Ƿ��I���d�;,��0��he�hy�w��Ԭ�����A�T~�o)o��?�'+[��:������n�-��L�����H��Mi�S���ӗ�^j�~�Ȭ{�;�!&I���˙K���ZN#��r�rX�6Z��Uy��$�`TEw"�qLR��Q
�cy��W���V4L`�癢<5��]��AP8��(PUj˔�x�(�4h>��5�}XT�А�aEARC҇�
RR>��H�yH��e�1���5�=0j�(�I�_1\�s�ӭ�cxm���l�us��ڮ㘮h��*.P�(��8ĵd����l2�)nS���)2�n�Dw��O��#n]`��&���[#�����|���Cӟ0v���1����qʊ�!~4n�w��*��9ǽ�?�e��r��'}!�����P5=>��f�E�X�
X�,	X�&X�HPHI_	����H�z5���^�:Xիr�zU頠����W�FI6HV[�6��C�zF��=* ��n%<�b4W+�PK
    +Q�H9�	�_  n    org/bridj/ann/Convention.class  n      _      �R�N�@=#`Q��cэ�;76�h#��jb\���25m!��\�~��&�Aݜ��s�̝����7 ��(�Q_�D~o�{R�f(�$?��@q��==�d_ov�M4��Uք�����j��Vg�/pX��s(��]
d�^0"��?�V��	4���uK`o����>%�<�ݷ��;y!&��-��y-�v[l���V�S�e�w�W�-�1�e9�f��v�{�m:��g�g���zl���e��I@6x˯��{rZ��Ά�v8��T��"oKI�xqL�@�1yH~�w�>O\�C<.���P�(�2�4l���&g[We�p~���e�[�ȫ�	�%,+(((*XQ��`��'PK
    +Q�H�kq�   �  !  org/bridj/ann/DisableDirect.class  �      �       ��OK�@����h��ڛ�X<���ٓ�HkK��x��!l�&�?�~5~ ?Tq҃E���������^~�Ɛp���
�*�e�3��,{��rA�A��ZY�%j����b�,�te�L��J]��O�U�F�h�g��!t���L�c����+���1�����v$�E8/���d�����'3��	_��{��"�;c�S�A-�/�ŔFvۮ\�	:�q0�T'r�D��l�����q��� PK
    +Q�H���  �    org/bridj/ann/Field.class  �            ��MO�@�ߡ`���ă�x z���Ʉ���z�-#.YZS�$�5� �:� �&�a���3_��_� .qH�K��ez<�T�x=�f�ͩZ(Ϩd��)�օC8YyO��:M��?�Fh�V�(PB�_�2b�I����29:��w���R���m|�qyJ��	[!O�����o\��~�KX���P�sv�y"쓶�ηBk�g�_Tn��z��Y�=md��Q.���Q�udx��;�
����G�+� ^'��@� bۢ�%\g4���B>����vq�� PK
    +Q�H�[��   �    org/bridj/ann/Forwardable.class  �      �       ��?O�0ş%P���B ��X�LZ�$U0H�9�)r���MZ��1��P�e�������=�>��? ��T`�|.So��e)'ί����R !0(�JK��\�iAY`G�b�e�U�2����e�O�u\޵�	UT6�V��Ҷ&��?֙�&�0$���ޏ���}N;���cK�T�7bS?��X�jG��yƱ�W��&��I��/��,�]y9�`{hN��`���}�z8�Q#_ �8�PK
    +Q�H�i�r�   �    org/bridj/ann/JNIBound.class  �      �       ��MK�@�ߍ��j�z<��C�.�=)F��b��&��B���?J��K�=̾�>�0������G��eZ�Y!���~<�v����B-�4��r�����.�+���W1D[��;輦N�D�9�K��R��Κ��М�OVo���(J�&7��e	����<;�X��L��ي�0~'�O�<����V��8���ӳ^�������@�x+�'@阮8��i�߶_:ة�.�u����oPK
    +Q�H��Y  S    org/bridj/ann/Library.class  S      Y      �QKO�@�V��@����@�b�ٓ�&`M�&�ӶqIٚ�B�_���G��������5�ُϷw 8����F�Wj�Uh��8�K7���z�"� p2CِZiU�ݫ����@i�s��N�sM>Y�yw)�8�Ɉ��H��DE68��]p�i��~�_�(K1���Ki�d�?�Ϸ��`�J,*O�<n��
n���Zû��C#�|��Z�WH���l*��J:&)�xݵzo�lcL&˟'�%� �5[j���(���td"�V	����N���2&4�gU�9c���PX�6�u����h��012���88�ZG�L�V��C����a��QΏ�/PK
    +Q�H � �  �    org/bridj/ann/Name.class  �            ���N�@��`�� �Ѹ ��Ƶ+�%�@K�`b\x����LIx5>�e�u!.Hܜ9���ɝ�������,��i�_�JS/P	�͹Z*Ϩ4���f�Ŗ������*��Ի��.����$NR�1�;��R��.6s���R+Wo�p�cM�2�8������/C6�|�盫"��Ď�:� ���يA7��?����՟���:����"�QO��ITp<�'��SC�,:8�ay����Ů��u����3�8�:�얲W�>�GB��PK
    +Q�H��G@�   �    org/bridj/ann/Namespace.class  �      �       ��AK�0����uS�ADD�0�b�ٓ�	���UA<������h�����?J��a�P�	��|}|�pT���J�*m�뜫������k�i���(���� ��w�R8�La��*�hz�����p��Xu���!��:��p��F�l]���`/|����6`'T���?dRd&^��qx�(�^^�)M]il"�;-�2�;��-��Z�9���D�_-x l��G�`OR���Ǿ�'���t�@�.���\1v��PK
    +Q�H5���   �    org/bridj/ann/Optional.class  �      �       ��AK�@����h�Z=��GϞ#�)1
�i��a��4)��y�������p�������Z|��1᤬2�T�=W�(T8�MYh��\/����T���>�目e��n���.��t�܄�C+qͅSׄ�Rۆ	���Қt%�=?����p֎ĺʸ�E�<�<��x5g1mO�x�:��TB{OeS�|g�|�4j�����I,o�]�:�x�TGrE��l�����|�������oPK
    +Q�H_���&  �    org/bridj/ann/Ptr.class  �      &      ���J�@�ϴ�i�O[�@D]ĥ��	�$�Q2m���&2�V�j.| J��`���3s?�ܙ�Ϸw �8d�*uF*�LQN���Н��prQ�N4�ʱ�Qg8]�\j���p�_k�bhRƅ���R�
5�\^3�*�P��Է�"_H��j���L��^LX�È�<��g�{��b��7�a�z�6"ӊ�ĥ��0�UG'RS29
����e��W��}ȃ!]پ+j,�,�鏒q3���3z����}���`V��j���hRmQ��Kb[F�����g�]�}PK
    +Q�H�#M�  �    org/bridj/ann/Runtime.class  �            ���J�@������j�x� E/ϞD*�(1
�i�q�v#ɦ�W���P�T��P�;3�f`v?>����K�ˋ4�=�emV��	� B'SSe��.�8q>�޲*�SN�6��	}4�Ŝ�9&\�l�T��;'4��TL8Z��'l]4{e�^�4Wې�P�D��!���d&�n����S����x,�{|�]U�Rm��U��6���b�G]����q�>��5� �Mt$�a����+wu��i>�-l�=����6�PK
    +Q�H Ew �   �  !  org/bridj/ann/SetsLastError.class  �      �       ��OK�@����h�W{��]<{QhmI� �6q�Y�l
�j� ~(q��"���c����|~� ��@�Ժ\�N�R��\��&��sօ�B��4���,-(�!��7]ƬW^�R���]�����NZј<���讔�I`�un������Cr?��ڑD��<;/�瑡%g&�7b��4J�fc�N�<�����.�[m�S'q͏/�IW:5�Y�	�y4'@���8�{�j�g�������6��PK
    +Q�H�]�ߏ  �    org/bridj/ann/Struct.class  �      �      ���J�@��5�j��\O/Dz�+z�4
��6]��m"�F�G���ԉ+�j.&3���mv��o�/ ���0FM��F��A`�t��:�0���R<hZ�zK���P��5�2��4�A�\��zVK}g<5�>`|�*�}E%�"��� sήVj�{a{U�FO�b�a�\�Ϊ����y�a�?��H�h��y���Hƌ{Q���T'��ԢAf��w�ֶc��Ð��B5�0	4�c�D;��I��6�����7��xh���1�Ӵ�f�=�=�q�E�l\'���z����Z�D�8��y��X�ť�e]��z�&� LЩ�%2M�f�Z��p0G�|���+,"O���i�X�b�Sʠ@�]���k�Y��0���4�c"m
Lb
��PK
    +Q�H�9��  �    org/bridj/ann/Symbol.class  �            ���N�@���b�A���qAԅ�kWK$J��İ��2��$����2�j".Hܜ9���ɝ�����MB#�/���ԓi�E�Y�D�O�RzF���S5�.�g�[�3+��R��׺(j?57K8�m��'���Ki�p��󍚩Ԋիb���Gm��t��a��ǀ�#��>�|sU�,7���?�03z�b�G��sk��j�'�\�	�([��цq.8?SOz�c�֛��%8�iy��*8bW��h�y�n����B�Bv�+dţB�_PK
    +Q�Hb�_JC  "    org/bridj/ann/Template.class  "      C      ��KK�@���al��j����.�AlE�>h� ]M�5L�$%���\��Q�MA�Pp3sϝ�y}|��8Ǟ@5]{���-}�vțjiȂ(N�L�Z���Mhl,��]vF���Oi!+P�:Kh���JW��Iu!��I�@��h5����?v��vK�`�ő�K�ɣ��-Mg:�)1��n9wݦ@�y�qh��d��w�e1���Pz�Q$P��L�|���@��4q����ȹ<�b��|�&��X�q8�[�ٺߏ��=�H�4-�!�B|j��T�wD��n�Pf]��
��pѬ.F5��\��r���6�r����d��PK
    +Q�H��{�   �    org/bridj/ann/Union.class  �             ��OK�@������?՞<�"أ�gOR#
�)�FO�8���FҤЯ����g{���{�}���c������âLe\f�����f�� �^ii�Me�T���.�E�+��ݟ���mR�*p��h	�"�ԭ@w�MM��Ya�d�/���i��5[�.S���l����������W���@G��8�?�sFc�|ͼ�˄2�+��5����l�ņ��/G-t�ip���M�p���]��z�c��7�	8t�ȕ�/PK
    +Q�H��.n
  �    org/bridj/ann/Virtual.class  �      
      �PMK�@}Ӵ�֪�Q<��x�$4b�Z��O�:��D�M�̓?��NA�%�\�;f�����%��Y>Uqn^��T�M�
m}���VV�S5��8��C�3Y��������s�N�*M#v�����ж`B��Cf�d)�t���pTm�t>e'��j>�<��h��"Z��O���C�[��-���.�#��"����2�����f<6s[.����:$WMuB��u��Bt��X��]y��d����
>����PK
    +Q�HoL��)  O    org/bridj/cpp/CPPObject.class  O      )      }R�n�@=�w��A-)�Q^M]�B,��PE EJ!�U6]M�Q�ȱ��8{~�U$| ��c�IJS�{}��y�����װv|5�{J���v����
G�����3�BG_����WC>��Ԟwsϳ����#Qc�N�
���5�yӖ���Zt��#��3l��j�ڧ<���H=�u�7��.���I�b�-�Nh4W���'��a��֊�`�!��J�\��L3V�_z�o�NL�e��D�����Ō��5:G�Հ���3TЮ/��֍w��{�	�5Ԁa��a�5���ѵ���g`-�Q�`�L<�CE��i�}
[m��n�+�{�87s���QO�پ��-�l����{JK7�P<�C刏ҐV��ՕcI*��5ג���G�� `�VP����V�&�!OyC��d�)6~D-O�[�Al��g��T���1��G@�������ы)n�tD�(�
���ND��]Th��L�Զ)�Րû��A$��8>'fg�h��{s�V�����O*��I;������U#�,)��T�V�A�/PK
    +Q�H��	  ^     org/bridj/cpp/CPPRuntime$1.class  ^      	      �U�NQ��.�E��o�j�R
��"(�h� !�Z�X��n�[����h"`$Q��� �K��l���M��әof��fN��χ� ư��c9��uG�m'4�N�_LW��1	��y[�U�jn&��os͕`���Jj>����+����O﹎���#�������RI�gP4��.��ʰ͖9:|� �����`�?�&e�p��W��]Ո���@-��x�$�F	2��;�c�����#�T��E�tSw�QXE�����0ZP��$N]2��"N=�����/�Z�3�
:}�Z��_�F�
�ℐ��B�M�J�F�55ON7�J��I�u����M�.�۠��.w�-f��Uh5��Z�A�Bh����-)��Ӹ��)a����_r�ܜ-�F�Ӽ'B��,E�b�PT6���StS�ӞwUS�ʤR�q�j���1�֤���&g*훸%��>YE��Ȼ"�C�k�m���&1%�����ys5�0tT�	�T����}Fjإk�Z�U4>)+G�YKS��K�,���n���:wJ�ВUp4>�{V�X�sw�"��irǛ��Bw�� ��fq� ��y;]0�����zB�i/�,��}t������7v�Ko=t�V��"�2U ���,�h����\�)S��d���]����ǿ��F֎0�v�����b� Ӈx�)N����H�9)�S�J��#��P�F}�	%ht����4�?����������$!K{-�e��)L�?A�6�PK
    +Q�H���  �     org/bridj/cpp/CPPRuntime$2.class  �            ���n�@��uB�$�	-�6-�� �Sjhဂ�D�TɅ�TROgI9v�v*x+��x ����B�z������w�����7 �a1Tٷ���,g4�ڝ��؏ܡ�m�`�?������;N�#��D�u �Ӡw�~$��ty���"ɝ(�:�0���[1�aY��1ǰ�H�#q��Mݞ���G2�c[�2�[
(2�(��C�a������)wƽ�#�����-D�nX{D"��8����ú:�R
�q=7\�Bl�0d�g	�d�Ɛ�u2��_�M:u���fM;�ub�߬T�ٝA�5H�e���E�c�a��È�q�V�$j�aZf1y��.9�Ig^�!�.��`����Q<��c��x9v���^c�=7q������O{����}!�2���kt�Tuh�r\�V��4K�A�Y��9Ck�l�c��<G���[�@�f�ɍ۸Ck�F.��As���S4?��������5A��=�O E<@���؟��d�xHky��EV�<��T�����Q��PK
    +Q�H%�UD  �     org/bridj/cpp/CPPRuntime$3.class  �      D      �TQo�P�. ݰs���8��:�|��l		N�s��t)WVRZҖE��&���g��W�-�eRl�{O�~�;߽���_�� x������;�����p�7��#�7�XS�2}~�u��=�I�/_A�a/2��O���ۡ8��;�8x���W���9w[J3�Di)�c�4\�}1C��e�u���-��_��˭�1\W��U����g�*���aq�cX�`&��I�)�v��|@<�dH���Wܡ6D���#�6�}�M��j�|�"��<bXVqi���`QF���,a-����Z�m�Ȏ"��3N�NI�U���P�w�$ӗ�+�Cn�Q���l�	��.�R(����B
�s����6C>�=M� �-���i�.]On���m��f����3&�r��L[��N��3g���>؆�x���Amڶp��6�[	� ���F�S��ZL?��K�N,��� ��2��:F^[��}���{�V��2�U��
�N�&nO��;N{N��|�#J/�v�B{�Wj#�L�dTA5��>��%�S����O���
j�'S�GQ���'I�BR�PK
    +Q�H?+y�  �     org/bridj/cpp/CPPRuntime$4.class  �      �      �T]S�@=K+��|�g�i
��"�b�f*2�<0>��+�I�N�2�_���/�8#����G9�M3���L���={�ܳw����� n�)è��e߮�V����_��Ю�ܒƐ92�M�1��E��[���lkז�Ǽd�}�o�vղ�Y��ܗp���Ź(�F�Δ���s�â��_�B�gx��Z"��Fۄ��:$K�mԸQJ�el�ۖ��Y����k���
d\f�i!*�J܎M��͔�qm�0L�������3'���O՞v�A>6����0uF�m�]R�dk�+�%<���M��R���b�v�ʰ�&�.P��!���F�с	W1$�)��u��*0c�!#�CZhfO��[���9�]�9�g��&�-B���Gm��-��%�:�5�O+*�ǂ�[
���h$��]���$5ѣ3�o�L/u���j��!N���D��)�������r1�{u�?M��)zj���g���d��+z�%��[�j�����}�o���3�r������Ы0(�����f K��B*��P�N�"u}�:�?�qB�P�� ��	&��d��Lk�0�9B?�Q!4a0��h���xG��|����]-h_��
���w�� Yd��Sx��/�Ps_�/�e��:�=q?���PL��T�Q6�*~=Ƞ�V:1����?PK
    +Q�H<Qe:  �     org/bridj/cpp/CPPRuntime$5.class  �      :      �S]oA=�
n��jk��V��R����AM��d��m�з�e�%�.�H�O��XM|���2�]�@�%n�3w�9�̙���� �u�_�uK8��n��z������N���
C�kM�5�����r[*H2�MW��rñ�)F��Q���W������S�ZHưWS�u��6�G<�b`K_0�ec���AИ���K���Q�7�Y���M
��*����;��x���:�\L��`�as1TA�!=�3��T��7o��E��"��h<4ݒ$S"����H�d�	J�t	b�	Q�ϑ/j�x��ʹ��� �M�F[�r�)b'�0�B������mVÂ�iT.h�=S����z�6U.TT�e�C�J�����J�����+�o��)�r�Y���7�z���?6�D�מ�����Է��E���"�R UH
�� �d,���Eܣ�N�3'��k�K��.��}C�s<�V% ������Hi&��}�'4/g��l����ǉ	A=D��M�~���^��S�Q��9�L�4nb5�!��R��PK
    +Q�HM�~�  �     org/bridj/cpp/CPPRuntime$6.class  �      �      �UkWU�7I��i)��b��؆��>ؒ�m	��Z�$���a&kf������%��k��%.�����wh��~Ƚ'����>�����O� ��o��Y��fc�Po�
���ն��23��2v��e��ږ��qD��ZqLۗnfUZ���)��=�
@�bX�8gl��:�b<�Vz�]�a1ram�%�G�K��y�Jy���Y1k���'*�,�RxM�Zh�4�J�w�u�aR�N;ꃏcP ��"�cX���X>L^y5� g+�Ɗo�M���dGB�(��6�9�����Ђ�"��up1�.i8�ae���<F���@4�|Fq%���)����I>�v�)0���(�Rn��y��8����n
�'r�'1�I��,��k����i5T�n�PP����/u��|îK���K�����'p�55Z-i7��J��I酄�����*�{�=�mߴ
�xq�O��N��d�$�!���(���iz�h4\�y�,)Ͼ��3�/a��bz���{��RM�w�`�8��#�7M�],�0�E�g"�{,F6$����)�b�������/a9�?�`/�HQpe�aU���&H��%X�����)��#�K�����^t��N��l94=�<��&ӢL���ͱ#�N�����L��4��tũֺ�F͒kja*�-���5�vOF��Q݋d�lچ�vi��03���T�i�u�h�v�r<�sI����ݷm�?�҃����GtpP�7����|��D���j���p.�����.����p�����U�7}��[�����o\��:���V�L}�ٟQx|����1���1C+=�%��;�R�\?�'��}~�G�+�x�vG]���\��RQ�Tt�ѥ�����4(�g0HE>'����2"�c �nG��B�/,E��j�l�6��Xq��cHg+x%zgcɠ|
0��@�?PK
    +Q�HM�j        org/bridj/cpp/CPPRuntime$7.class               �S�k�@~����Y��p��sj���l�C��T%��f�}��g��&%I���"8?��G���n�w�{�{���~����C<bX���aN�o�á�::�0�"g �����cn���ﭾ�#Y��ٮC9ca:V���v<X��¶�0��k�gC�1���Tp��]�� q��[�`x\5g*��%��d(�f��f�"n0l�1 �!���T�`s�WC��S<�JJg��60̍��E����0d�?w�x�I�Q�	�}�3��z�xN���QM�]b��U�`��n���e��f�Veew��a�!'50l�RkR�Ơ��p����)��GvO��v�zY쩊�QB������ًN��;D�`�6w�<pd��_�t<q8X"HV���(��k'.��l�����z~�A}�y"���[�[�
�JE	P$k�=eh�a��{�=��,Ų^?Æ�w�M��~��hV	He��}�y���H�����%q����wԾ�#X���Ӷ�'R`�x�s�Q�݃Tf���+��y�䱈�|�/PK
    +Q�H�ڒ�h  s  ,  org/bridj/cpp/CPPRuntime$CPPDestructor.class  s      h      �PMK1}i���[������H���YeEP)*��۠�k"��B�'��?�%Nj��P1�y3�73/����	��}m���ݞ���A�u��T��=r/E��,J�q��cn��ãgy�ʸ�������\)?Ъ/���	C���L04�����A,�:��$;�a}�P%��Z��[�(Ot�丨��!�a�T*��1�mU,��`��IIC3���7n�Fz@�͛�6A��4���mn$����Zj(���^:2�{��H\Ix�J	�<I���f�e"�|��N��K��"G��ɁY�d�����p������Y�7�U�nҝ��ܮCC��<����	���0�)bX<�a��e�����,�?PK
    +Q�H����  �%  *  org/bridj/cpp/CPPRuntime$CPPTypeInfo.class  �%      �      �Z	x�~��f7�l BH Y B�A@$� W���]6X��������ֳ�K[���V�V�Dڪ���U��P{h�<���g&��ݙ`yff����{������� ���xbcÆD�ssC����e�ʶ�X*ҭ��c{��$��@̝�1�5�zņ�j8��lYi19�������$0*�.�� �7���Nq%�r��P"�UnK%B�T<�G`��F���wLs��LMm�w:�	��C Pb����\kxP&Pܒ���Ь�Gb)5QӦF�PR��r�!9�T�	J���P"������)��'J�*�%�׷J�7DC���_�Q��P�3X�қ�D��zH~�7�-<jW�L�̬�Kf�+��6����vv �n>Nt�|P��Z��Nm�$k�Ћ�<$��H,�j�^�L怳�n�c1�8Y���&����^�V`Xf�f�3yIz`0mTS�����̲���C=&y�d�I֢�����N#��֭�'d<�xшi>�@��}w��2G�S57y0���Z�-���"��*3��D$�q~o$�)k��R�[�ً98�����a�C==j�S`��J:�~��ǖ�`�d�P�C�,'f��6wI��b�9Sx�?:GM�ez�{L�c�X*���a��0�*�Piʬ��	�H!bS&9{ݦd�Ў/�r��)�s��K�(Obgjc_��pL�M�;�Y�p��J
#�����cN3pc�֖P2�$�L�ba�I�8uA�1����Mz��DXX��!���"!�h�R�SE���Pt^8�&����r�{��X�B��s-�$�%�w�t�e�9L�~z.'���pݲlĘ-��G�'+�gؽ�֮J$�����4X��i�D�Q��ٗl�V��F�%��<�蘱-c#���z`��3^|���3��g~lG6�B��U[k������y\ +��I5��3��]'��"|Q��gF^&�&�ɨ�K�Kp��p�vQ(U;����+��Hm8c$�%�
��)Qa
T�u�P3�w�X(��a4�GRF�)"�&󲄚�G��f�h�����F�sq���涳�
����,>��.�ײ���kN��::������E�6=�%D��a��[R�cx!3�t9C��ӏ���虼#����|��q��ͭ��KݼN�~	J��*cN�i�>��h�4��3���PrV�zq��<J���C��Xl���X)��_�}8�('T�p�T��!J�饔�6R�Q��8,�> 0��,=���'�rct��X`��v�(��!^<,��Pq.Lr�\ѥ�K}x������.�Me�ej}yF�M��V�σ'e�� �i�<2DBQ2���K�m�g������L����C������]�ژY��|�8>!��K�=�Ӏ9�.Ë���DC�g�ׯ�&K��ɝ�+�ٗ6�l����U9���}%��s�-!P����d�=�S�]1����|^�z�'r�$��C\��I��>���&�ӈ@uj��	����o�<��ѓ1f��g�1��gZ��xS��[ȶFR�2m4�l��Jf�Ŀ��k��o����5�-�>�O�z��H�9�S��+�H�?�_{T�m�ܬ3s�$�Vg�G?m70ۄ���Bӧ�\_w��}N۹JxD- �Y/BڨY3e
�ݫ�}g��l���
�*�ᓢJ9�e���YV�g3�%�H��$L���ēyJa2��9��U}()�̵K�P��5�y�N��R��h<F�i��+�$���-���{{z≔j9މQSuuNQ-N�ꎡB�*��o�)�"gQ��!�˳���\��5b�<�:��;Ǌq���6�6E����))'I�Fy�*]��w�><�u,q�L����t��-G'WK�����<�F�zgGH;�����[#4o���7^��ϵu��e�	䔑g&��?��du4�:�H'vX?��@^��'��C?h���Pp��}�`=��:���w��xo"�.����-��Ԅ����X��B��ɏ�|rɯT�8xC�S�T��xc��/+�Z�\�PÕ�����x��aB X�u�а<0)������=8�zL�?��vb�!4�=�9k�c���i,"�Rކ��Ɗ�h{  ����f/�*�4^�P���zi���d3%�,��7:�:�������_�x6�r1
�KP�\�2�2T)�c�r�*W�]��zp�$=����}[��(	�G���H��5���e�����
��1���5uV���*L�s����*t�qq��:�˹{��ʽ�"����VC|��uC605_L+����
ܨ�|_���ь���x4'���I�V��k�$��ŰUu�&-$4I;�ܮ"7�j�Iu6����\�"��i*���Wv�I���B�m|�F�Q�&��x:хM،�/b��[��'%]�)=�ԧq]� �S�=Y�����i�
��F|�<2�������&�%�r�!�������璻�H���ۂ�q�b�Mᥦ�R���(О$k���0J5��m�ә$;�ˀq+�H5�{Ơ�!�E�߽{���`��hY�����e�⾵�∂��-�d�n� � K�?ď�Y�Ʉ*��>���W�G�C���+w�F��)��s	7n���`?��7}�K��?��'���y����A¿���#��	�0�1��#?5�25���O�Ə�n��/u ���
�8�!^��k�5$�fV�gZ���6��՚��3�����J���y�
�<��@�5C��0�f����Q�j�`���R-�������]y�u�q��4�S(W��d%'C�]�O�o;P�yL�M�i��j�ǻ,Z���z^��)�so�'MO6
!���P)��Փ��'������?��<�+/`��"����ɋ�x��R�-"�w�;�_T��*ͤ�� ZaU�V�[T�5HrP^�_!�W8-�@~;0���,{D[�(��A��r���U�Z+xa�;��{B��=jRZx�A�`�r�(�/�w���ħ�&����/���1MTi�*L�쁲���z��z�	����*���x���Y4֫�kL���U�`Լ��ꔷ1Gyg(�S��U���5p'�_�c�h��tk(���E�^f�-��Z�����,����#<.��o\|?����Ϝ������W��*L�"G�0�
�P-�]^C�"R�s�Ы��ɝÂGE�N�I�oO���I����3%ӆa)3�,�����J��UV6�j��V�-iдd�Wl
)AQ�OHqN-���y�2l��|r���<㢲y�k��b�&���g3Z�M��T�Ҟ�8.S�8օ��i&�6"�Ѥ�x5��i15�BxM�^S�W4�B�㵕����"���2�;��"ٽ�r��k5��bF�7�&d7!��ۆ������-@��	͝��C?!(����5�r�����c��b��&�B��	��pT���PK
    +Q�HQ����   0  9  org/bridj/cpp/CPPRuntime$ClassTypeVariableExtractor.class  0      �       u�AK�@��Ę�1b��s��"s�@C[�o�$�I�lD�Z� ��i=H�0��{?��o ��!<5f/sS�U�h[�dٺ�m���D���~���L�r�ϟ֨�6F��J}(�U������
\nO��0;w�)��v-鿘�ߧ�"�w����Mӛ���fB�R�l�8�ك�a�'\!t���q_"r7����PK
    +Q�H��؎�  Q  .  org/bridj/cpp/CPPRuntime$MemoryOperators.class  Q      �      �V�wU�M�vi�@[�ޅb� ��/�Z��Jk���R�ɥlI7a�)*��~+>�x�ңD�G��G���蟢�ݍy��q�����;�3���}v��O�������G��x<��ٹ;iX����)�cfjW\��3
�P>��h��fv����E�����
�E��*(a���󢈈a�����y��e@���>���Sk+(#�fL�Go��
�8�9l���Lcٕ�ETJ�g�:���Z4��l�'����F�%f�p4z̨�RQ�X���|^B����P[�",	f�[S�6��ےFX46M~ڔs��K�M���f�*c𭦩�l�����O���OOL��Hs�,XI�n�V3���Q�5�������p��e����f�#"����j��!���}4,�N����X)XG�
˩6���W�\+i�Q�E4*�Ԫ�G�����0������Y��DK��CjO��:\_�M��P9�\�Me���Q�N�h,�f4q�[<�_��e�f�"��T�S�f&D�n�u�?Ӟd�mh���ٌ�8|�P����z���HHb��s���;p[) �,�����ċ����ê�N9�F"�H$��u�؍.y�nBńP��)�;��XƲ��Q7�a8�;��A/��J6S�4t����w�P̚v�E��{ػ����F.�͈�`a7����M1!T�M�?�b)����m(��*�99䜷ڭ�BwDC�����dYk��U�n��H<�?���G cY���(#X���ЕHj�%�= $�^��U�s�/��� x'�C�7c6��L!{��`/d�I��a�Z<e�Z_�j�G���q��`�q�:� ��tAV8E~��r�V���-�]�?ω�[r�~i�- ���H�_�����AC��&�w��"�Tca-ڣ��6��;'�"��|HK�[�	�*��1*l"���X��6]*��!̖��H��9X7��r����yW��_q�~eξ�����%,�K�`�&^��b�I\s�Vy�UG�Z�x=�_��N�M��l5� :�Y	\� kǱ�4n$�\w7�㇭�������=����1�����cX��;N��*{�_��>W�ޮq�?�8��1쟉^�L�N��f�|c����M�W��>�w�	�c5.�֦�
����i�ǻH��<]�$FXV��p�pa. ��2o��Τ|����nC9g���sT�Y��9�ӗ�L_���}�#tG�[|H��}���#.�E\���]b���>d1C\����@��}�3�۷�$�=q�g*\eǵ8�b<���q�����iʼŻ�}<�}����Y<����������Z	�+	�ʁ��@W�E�� og�+%/��9����{��;|�JA����`�f1[�S1��u#g���4���b6�sy-/)�*�A��TTm�bgn��?PK
    +Q�Hg����   E  :  org/bridj/cpp/CPPRuntime$MethodTypeVariableExtractor.class  E      �       }�Ok�@���o5F�Q��C{qz�Q*��J/�6qԄm6kѯ�C?�JL����9�<������@-�Kb��7�2�A���d2��6����&Y��)(*_������!R_Jj��q`ʄ���W��5��A�E�O�?=�����{���t����Y�5C��-����2��oJ���prUB�p����k�	PK
    +Q�H>��x  |  %  org/bridj/cpp/CPPRuntime$VTable.class  |      x      �Q�J�@=�Ʀ�ն���
>h��-)�BԢR�q���֘�����A?��'Q,���ffΜ�=g����`�P�mW����F#���ǁ��b�{�]_�`�!��σ�}���MdJc�^B`X�k��C�c"Cv�C��;��P�ݟh���j��]��ܻ�H�������>���w��m(q��D�A�k��B�)�[$z{�[D	e*���#h����YT�(b���=��m��g͉����m�h�=
3NH�\Ʉ󹽒#qߺB}"�E+Oʤ(�Pm�G���A2��:X`XN�I��ʯz�2$�(�P�B6E��G�ԟ1{���,ܧ���v��"�(�ѱ�W2��5e�)s���(7�G�PK
    +Q�H�g�P$  �  '  org/bridj/cpp/CPPRuntime$VirtMeth.class  �      $      �OMK1�ׯ���������zp�x)ªE���nڦ�fK6�y<��Q�K��$2�7�����z� p�=B�0�06*���l��ǹ�*�GCe이D�Lŋ3���C<���P%�W�sg ����C����Ih�|��\j+�*4� ZE9�8#t�"�$��)���ƕ;^�'�� 6|��"��D����ߙ�e�_��Ѝ�DdCa��3��犔���<��G񟊹I�rEp��4�L��,�C������[���;�.W!31����~]<�b�":�d���p
����U�.��j��PK
    +Q�H�I�^2  �x    org/bridj/cpp/CPPRuntime.class  �x      ^2      �}y`T������d�	$0l{��&;a1�d��L�� ��k�nժ����TBE\
jm�V[���u�V��_�V�}�}o޼If����̛��r�Y?�����}d/�q-�w,�zԪx���Q�--��.<�5��4�]$��V[����t����ֆ�5�\.Z���6�\�'(�vCБ9�-YZՄ�<��kAú�ef8����'cq�u˸%�$g����X|���p<��	b�n
���H<9?�\�"A��/A㺘1�&��\X�Gxm��%�!�v���]4tTn.4�����'�s<�9����y���w�|������8���Q.���.���1..(�~^JFֆg�i2N��ij�E#2�!�����̦�T�)��PS�5�HA���M��nEW7E��G�4.��!u�WŚ\4FЀ����(؉�>����B�W��Ǉ]T)�c�4� =gZ7g���$#����T��A�L�"�$8>�%��I�ztz�)��T��0�sS�N���zfo�j���5�:�v^dU<_o�yz=��$��+G[+� �C�pB���Xtm8�,R�\�N�����E�9uC�����[tJ��ںE�/�^��xA�F}������f����V�k�uZCM��%�c� |V�<�ΣZ���Q�C-�yg��	���ä�)m�j �����)�Z���%��;T���ÓDbњPrf,����׭�&ׄ���%����S]N���;v���Ʀp}r�Y��3�mTP;7��3ɽ(#�Y|��h*�`�hǱ�c�{C�x�	���6����Ps�~vk���Eϟ��M����`�gp�M��;�PGOߟ��֣�R��Lwbf$�#6@���YM�D#IX�*��G�i���SH�vl(�3��4/5Q�G�i��$E;��V���K�s�崂[%|t�Ѿ�G�Wg�(d\��Q�qu� GrM+퓓A����d���CI����qa���0��d�z�B[������8�>�ݭM�хt��6�Ő�d��s�����:8"��2ܜ����~�K�2��p;�Rϯ�k��&��%#:��j/]I�  v��	pѵx�+7�4��ᅡx�9��!��t毹�άZ1�#���'t��A�Ȓ\,�����M^��6c�K�s1:\�����M�����NvZ��~������fX�����bXI��-�.ږOw�ݐM�5��^X`���b���@N�%��6��Ɍ�h�ۼC�[�2��ACw~b�93�`�у��هp��Lw�@tm�.���
��]�;rp4O1�E{`�:��1H,��ƒ!��f��;!��t/P�8���^z�*��t6D�L;��..� �/���������ji	G�+�D�2���<G�䱞7�P-�^�t���0�/�������z^<y	Ɩ�|�
��O�E�lDi�������jE���<C�,^�?�ӣ�A6�'���vj�(HK����ӊ3=��@��LK̋$`4CK�9[��f �mz�K�w;�9�wf��̋�	l��NPl%����c�Adq�:��[1V���rm���͊,Z�}̜��2'gBц�%���N���է�C ,:ܤ�M�����k�؜��W�6�5(�[���}��y>=D��T#�t��gc�r}I_�Z}�05r0��t������s��W�~Q�рJ�@D��;�S�-,�,�;�&6�:����)�Q;�2Ύ>ЅOLw��6�ׁ;��1t�a�Ь��#}wњx�]�=0gZ��cMLc<�(�2$"�-&cQ/A�Ȯk��\�'���W!z�%-�`�ч3NF4��P��K:̣]���)@�\���˲h�}tڇC����*�hq�Dm�>8W|Iu�8��c�m\b���愣P���aX^�$%%��]���01<_%p��{X��f�]�4_�q�)F�
V���Vo9����7ք��ܢ�}Aڋ�p�Q��
�.1X�ĳv-��aX\�ĸ|1V��yd�^����a�,h��Ij|�Q�/�s����ެ��������ɂn1x(Xkl����T�j�t�b:\���6"���5���a��Q��tX�An ���؃!އ���1�ߐ,�;��D���D��Q�d<��Å�;���������1IW�ʥ7�.rݜC���H�	�Feq����5�Y��BP��Ė�̐n�^�Є�^tY>�aF#�K�R�FH��]q����`X����j���2�h4����0*=�O�Ar)V����0�%���ߋ�i��� ��hG4)\b�CS�1����,�i�ɚe�cMZ��(�d��n(R1p�A���@F�3��T!�^}r�u�����'=�+����	?3g���<AG��sĹ�S�h% �t������\yb����g�SMU�|�bq�W����<��������C�	V���'uQ�3wm4��w$��`bqr�!� Ҍ���b͎ǚ�s{�O\#~�*�5º֖p����p�d��>���(s@���4�-K7X��=@���7��y�[�I��F���0b�˖Ɖ-�6/�?5�Yf𰂵��>q;}Φyۚ��	q{�aC���<>q��y�XܛQq2�v��a��ӡp��g����s�9�X�6�L��:�@�5��U����9԰�v�Y;�R1� ��c]� �� q�6�8}xI�!b���^�j'���c�=���Ma��&��aqgc�:�$Cڧ8mh��Ԅ��${c^�/�~�� <��f�7���և<�o��n�m���6�*�4���"SM�΍��5/+G����~�v��h���d*Ʃ�J�"�(��)Ō������5'w];eڇ�0���W�O��FY0ř��8��J����]��io��.�N��k"�Q�#M��Xr6\^C��$�U`�k�4F�`)��w�x�'�oz�!�
OjiiZ�ؕkI�I��F���E�[���	���bG��M|��!���zCC<̡�h�O|$>��X�]�LB]�SD��ٱ��xC����Pǒ���)�����C�՝��Ŀ1	�C0���JPa2f�U�&���0��#hV*3-'��5�$��A?���t�U� �ĚֆR�F��7#��;�)��յ�>)����2
��MpI'G�D{�z^9�P�n�̓K�[q��-wpL�K��Je7P�^պ�'���Av��o��e�.�%�����X<��T���d�<r䢣#�I|�����`3��h��A�Wے�x5�Z��Ɛ���)7XnH��p�[��!�(�K0�8n�5k�К�n�,،��8j��4�(!.���<���q9��9}�\��x�ሶ-�R.�Y�0�dn�;R)��#d����2Ae��j�֥~��D�T�UCY�4.xF�`e#��s{S6:wO1�%[�`���U��[��26)�Z�D39Vs���`.�%3F�e6e�gG�l1IȴMc��af�ď46�&�um̌H=.a�~�rf(h(jZ� 5�7�`V�3e�tM8�0� �z��p� �KZ���Y�T>1�-y{3a頩�l�0��r
���*h"XjB���I�	�L��@�1�d�=J	ߑ�b�d�� f�$̸0�=>�t(�)���
7d7�^Xx,Χ	BM�O��=�޷[K�ҕe���2+�\s2�,sg.S1��Y��kU�|Ѡ�CD��쇓J= T7�P�.�(���j��dn�wp�HC`g��jcu��k�fi�!b׊3��N4*�y2!�����!¦e	p��N�j���I��*�ON�\�;�����Po��� /��]>D�H��¥F����ay����U�ml��	���؂��eeny:LM��ٴ*�V`.%�ɄLr�k�Jhnw�5	v�`Ji�)�V�<r&��S�l�niɬ�������v�R�N7�M�!m��dy�܀<Y^� kn�X^�a�c�ta�P^Ƹs���YО˘��(�<���J>��Y��h�[^E��-��ݓ�N��MMny-|
2�D8��D�]��?����7������&ػ��	:���	[R޿�� 2�E��	rW���Tk<�?�[y��9�4F��o�qdb��Fϻ�`v�K�6��pp�[�ulh��1M��M���!5H���X�p.�������� �";X�,�%��UK�k����2N���X�Ì��o�ԧUx��5�Z��3�G��`C�s�ǽ6��`E�K�k�_9n��O>I��rF�$�"^����ǌ�{���m��$)��ia��Ƙ���04����u��%�3vlx��5���_>#H �<�Ō$��K��ijB:���G��9����,h�r��cֵ�1O�8M4�6��7\ޜ�R��~�%X+r�R0�D�W�ޓޑbS{�G����%IA�u�3Ë|�uc�?�k-a����V1���D�f���G|�N���!�d}|��U���|�5#i^��TUc��bޕ�勣��Я��]��=Pgmx]�'�.����G,j��x�$�<�?�'��S���L|�F��/#��}.�w�)���7s��:`e�ò��&������o�U��QB��kR��b��'��O�(��a=3�	!�8��g�U�.l�`G^}J*��9`G��>��u@��i�u����+�O>/��|x�r����	W��OK�T!�~��\�D��Z�F�U1c(�$J�9���P~��P���y�
j�p��B���̔�gf�S�ƾ�p�!��s����㼗�\��^�8K3�K��#�<H�q��O���3P%�&t��rGgn���B��#�q;.�~���P#��q����(6�M�j��37�m���=Fq"��b��@@�2���U�QH��:�ko�VH�����Ցh�� �T�t��tY�W�ۓ��A*���V�O���.]��C�'Hӧ��̵�v,C�:4G���K�df�Y�6��j�����s&��.���rF�fy6�m�=����z0&b8_�Y}-m�Z�@�N�5�Ʋ����� d#"��j�,�� ��ت��'���R����)T�wU��NPˀ��I?,�ٜ1�ʑ]��[�-��d�f���J����q�*�w��.��Ua����z�1C�KzB��\kY�!+4�(�[��TD��Uk�i��ϚH�����u0�YE=4O�2��X����;-[8˧t�G�U�(%vP���� �2w�{0:{��c5����*-�u��eo�Rg�b���X;:	�:[��Ug�s9xBc�uI8�E�P}اΧ5^Q�.��,ֻ�쓍H�A��^|8�mQ�z�iu�1&W��TH#�:� V���'6�,���Z��f'K/\VpBMO7[��
uZ���_"�I�A��Xow�}��tޘn��?�;]��xI�Q8�sX�:l�RP݄Hk�c�7�8�w�[��	�-���U�C'� �Ï��V�r��mȉ�}�����T�Swzi���2ȥ&ِ�\��]��^�Aei�e�qN��oĺ�1�=A�� ��>�3��Qm⁷:����a��f�Ƀ^�B��[��׵�Ly�����ݥ&��َv�f���2C�2 o����y���_�Ayv�6�马���T�9R��w�cj/����g�S�����j�,K��>:O=�UO���HRǏ�I��s��t�ە�C��� �3�,C���C��S������U���O�J���^`����L���zɫ檗}��F��·"Y��hć�;[��2�J�v��4xV�S�g�~�+�C]�������T�&�U��R�BI�i˟��V9~M��p���9T�·>}�:�~�K{�}�Zk7׭�E���W�Z��#	���+��}��J�7��i:���Pj�s�S��,�����`}��o�f�O\�>����S�����������
�6��w��'��^�R]�X�	75$j��)/z���xH������݇��a�o��K.�M�����j���Y����ݪ�i�y�F,pD6�������K���dm�m0TG�@Φ�- �^�Ğ����ǴCb`���R}-rx1U�O"1d���Ҥ�g��V��(�h��v��8�c�`��\/�d<���QȤw�֍�1�U��qñ�٤�&�-���x��z���ܴ&|�^la{��/�Ĵ��aa��Gu�Aϋ�F�y�z�>׶��y�gf3�|0��_(b��M�U� 9^L�K��F�^�Af?���� ���~'��'-��1��C7�!F�Tf�^��N���>�^G�Y�^kN��������d��\'�R,ZM���﹓]�m����u�m��bSL/{����{���������T߅���ꬱ��,��U�r�x��2]j��V��~J	|��$���]����R�Wg����0A�����R�z�b���0��f��F�qMp8AI������t	G������{>���/�i|pHo&-����y�����<��{%>C�߫�Yo��н7����!$�/��I?���x�hN�.:�t5-�E�;)���q�I��ݵ��u��3ӗg������3��s�\"� \"�&�!zQ�J}�0*/���I��f�l��<t�o�6P�@�)��t�>���C����F|^J����#'�B4��	ڸ�<�e��G��������u�������v�q��)Me��bP��n�[0l��[�6��Hs-Ɲ-��i�F.j�n�����ϙ��`9�	+]6�IQ[�0ݾ�z�W�n�G�>�������U���ǵ� ��H�pd}yP���^M�0z�~�)F?}¢ϸ��dP�"Jb�V\��gP_Z���4���i��<9-}��<0���V����e���|���Rfh-z����G�V9�4r=�l��=�F���/����(7����]����nB�7�ػ���wL��S�O�[�0{��{m�A�������qH|��-�����6��U�/Щ2ϟ��V�T�[Uz@^�����m�rs\�glU~��@~}���\~�En��G;�.�m߽� }����n���#h�.!��Zv&����#!)����B�x��F���I��)Ɋy�)X�{��Zƒz�J�nh@1J낃J��A���h���(y�%�	�������s[�a���������yxzt{�\H��"*����.��&�C��.���#�]����,Wc�k0珱�k�@�N���qt���I�B�ݴ��R��ʖU9�,���²�v�{'ݾ�F��ݢ����(X�,cg�ww�#���<�xj�W��;�����7��pQ&̡��f.-�������+� ����2�:�l���62�A��V�B�sp�=��z�V�}��1�t4�I3�n��{LH�g��=0"�?,�-F ؗ�e�aO�E9{�Gk+P�M}����6�*���[�*����&I�t�J��̫���9��[�Nz��(�ٱUހ�h��_;�����;n#��]���<��m߽�ϻ�f�)S0m�&g���6Q],feP6��ӕa����-A�`�gё�X�ڋ�s��75�QZ�=�Q#~�o����O�V,�pz��Zס�5�h�5�8\9��k��%�N,&�"�Nc�-Zx<+��jZ�`k��m�wf܍��~��fC���}z<_�$F{
��4l� ]K���,<�X�����}z�� D�%b�i��J�}ʴ�����e�bٔ=T�����.qb�W�--U���A�MU-�|q2�k�jO����$�UJit�xw�^���m���&m_�6��m�˟����O9��--k��{hزҀc�o/�'V�V��S���J�����]��"��p��`���&ь��R@DE�F�9?uP%u��a���]m.��v%���Dj���c�fX����i�z}��E��@��4�>�@�O1�g&;��D�8�d�b��Ls"�=�'8-�".��I8E+����~���7���֊3̩�L�D���	����h�q��� x}�~x,^\�l������ic��C�ďĕ�ԉ����8Q!�W�����0ڣUx}�@��"��՟�"H�b���aP�sĹ�B�1ww�Q�
s�fr����E�� ��k�+{�&�l3�|���<oo%{+8*�V��<vT���]l���;��U����;�RS�߷[������[���⾪�@���l��_��&�o�c����|�.�D�*ŘwgUa�Pw�)�Õg�hǠ����Q�f]��6�){������*_���]����?����C8��	-�@7C.ڍ�e� ��[<P�ÒS��8�g�s0�fZ"~��np/��`��+�����]7D�6�k����x!>�^�Q�E��K�i���XzM�,^��&�+��EU��xU�[������|�;�܊����:��-^�N��>�cN���t�-V�+��l�����а��@��� .�b4��D�q4XTR�8��UX�D�a���YL���J�it��I7�Yt��M?sh'\�>@����Y��WE-��m��O�q�Mǀ�E" �z:z��x���:���S���K��h#;2(,��f�s���"��%�������<iM@�<@�8���U�O � �<��l(>i���~��אp�B�F|D�o9XJ2�x�tlN��~W����:1�,xP��D����z �`��P��&{�F	@m+�Fd��7K/�ҜsHv:�����Z�+���7�K��V�����ئ{���k��ɒ���|�Φr���}7���0�)3!�mqe����`]Z��!�U�o�1<���#Uv�<�ﻉ����-T���ьf|�fd_��I�U�+A������83�3�M��XC��6wE�h��-� �AJ�*oYW;�LY��BQ%ʐ��v�Eo������v��[9��kqʖecʖe������g��B�s����gqU'�K�ɕr��=�b�p�M�J.�'��-G�e�0�T�0���m�	��'V �8	�)��4D���� |�4�g�5t���*q*�� ��f��A�=��^B�|����S�n�^tg�1�6U�\�d�X-.��H�..[�%�6q��&6��rцx�G\��R�)�o�k�'�:9\\/��&9Vl�G�����[%�݁��'�_���@9��쐟.YL��o�r �ɓ*��Jd �)`�F��M6,U���U.�& jg����~�.��~>d�<�T�0��D�3�!CN��X�z����)r5�"�=���y����
h��h�ԃ*䩐Z⽡K.(��%��	���d�V��vh��ם��ݐ�=ȥ�Rq/d� ��L���@y�l2�,��}D�ò� �e�]��W���/+�%��-��;O��˳�r������2jֆM@�ρb
�<��\���z� f��+�`�x0�o�ߣ�}�!(#�3��D1��Xqj-C�i��c��J㌦��Z\�+����G��G[����lK�������� 5}J��V6R<c��J�Щ��*'4����筼�M^���V�.��|W���&��r�N��TX��j]�����|��.����w���ʣ{N>H��|׭��̗#���̳������6Q���6y�&�ֶ���"�Ty�)�Iv�.��n򁌑�K/�N�~�4��� *O�K�;�5�N�g��0��i�d;��GrD�b�#,r�qJ����d�k�1T)�"���X���Nr|�%�0����A>���X��psKȏ;�������%��++��	�?pq��jL��N�:C:i�t���MOJ�$�������������a�Y��.����cA7�d���.Rh��o"�{b���^c��]��:(]��~��'�^x���I3���/;@�b��6K���6��gSշ�2C��~ihV�th�eA��}M�xÂl�����tH�7\N>�c��[�Ɖ�2GLp�tx��D?�<�R�@KOG�|Y��Z�w&��kv�Y�+z�k���q��� �Y�/3+n�2 _��%q 8N�Q��t >�՛X�J{)9�+�B�j�,�Z9��Q�T�1�Z���9�Ty��C�B���ra��S�a�Q\}��e��;�6ӣfBX�W�E� ��|U�
���Nb��X�&�W�	�!!�zX�����LG�k���W��M�����-�<En	��FUMm��1��@���q�K�4c5ͥe��y�mʹ�ʙ���+72��s?�����S^�V�.D�
�F=v�"A��6��U��b?��
8��_ �;�
xg�:��^$N������ms2'�p�����U��ϧE���M�q�/T����?r�<�J���ѻ����TAV(�O(�P"�R(\i���z\���
�B6�ZK�P��jUR/9��ɣi�<���*�$'�T9�N���IN���Jq9�Z�`�j:_Τ�,�ZΦ�;o:xTG� �N��_�Rz(�# �c�
Q-O����ɕi��7�L�cl��F�?�e��@N��N��v5�5�M�ة|��UfV��J�T��V�nWJ.3�[�ߝ���m�a��l�n���R�H��͞������jW� �<h��қR��U���U����`�h#��U�y�>�x���3dƨ�k.x��d#���c(�]��s%��* /�F^ZG%8�߂�����4��)�m�v����b$���僾�|��Zݤ��o�s��j�@���&��@+^0�K��j@?�m�&��טU_�q�n�q��c��b��N��z�f,cP�:J�N�d^-Iay����b����g�m�m�˳�Ny6�%ϡ�����|!7�j4������y]��~����y�D.�Xf��L���F�����Z���XR���m>��.R��K�+/�>�Vъ�̩A�
�!���Q������]��*'|�:��a_��z�K�m��ʕ���*S.�x]Oc�mTR��X�;����
���-+��g������X�uRz c��eWac@ݥ��r��L�pf�����J��F�p�u��{��lr�hj]����x�����A��j䷩�\�x���<�'�>&��0�mS�;
�"kA]b��}�ɽ�k����lrB��$�NC�q
Lo���_'�oCUn�BBΩs*7�#�F�#���	�w�a\K��xD7Z����+��u%���T꯮RWօ�m��n�<�-�v+_iCe�~��FCI�������Ju��	L�Hq��^�@y�Q4]Q�/��_���-���9�uf�\��WZ\EGʫi���F��i�����[��Mt��ü	>�� ��M��t���^�w���> e��
�E�|Pth�#A�S��*w�Z��8Q���=�A��F�r�}�錂�ܨ6�y���28�>�܄-ݪ��@���p��ͬ�N��c�[��n4!##�k$�����IQ7�qm�6����
L��) f0���q�9�O='%4:'%4:�Z!E�O��\w�m]�V�� ���� T�y0�W��:Q�� ��ɜ� �vu���w�U��z���]m���b��w��#�ߎv�7� (g�����+�AV'���S5�Q�|����6�Z�d#�XK3z���z��k䔯�E����T,��˸ۨ�����D��b?yP�n���+��u?u�C �s�z���)���\��,�2��2+ʕY�e�R����-C"e6�����b�;�M�K=�{H��G���S!g]�v�v��@�Uz_��:�ɛ?b9�G3�h�[�cWvo���\��}<��/zz��ճP�_U9�w��6Д\���o�G]��pv���0���^\��O����+�+ٕ���. ����9 ��,�:�Nu~u��l6�}�pn�%��?�\�������z�L�R��Ш)����[��z���=��Ou��x\4����q��\\����ڠ�\>�A����cyM�l쳃�)��ѾR髷�Q����iac=���9���L�n�0�b# د�ߐG���w��NR��(<��V*�U�Xy�*՝�S=�VUDw�b n?��?��ЯU_����j ���[j0���Їj��Nc�1T3L\�ub��|��f�&�����:����S��v�,�����{v�����H��x+-mS�A���}ͪ7�0L{�	�ƸB��|=����8Ԯ>��Fnk��30��{�2�c!��)�>�t���p���>s�����˘�1��z��߶SF�T�q￨9T���{���j1�~9U�t�:�NQ��Si�j�Ģt��AZ�Au:�R	zJ�EV��j:�r�H"�E>�.$jՙ��E���=�#��E�v�Y���!�t��n�`�]������r�25�(>���5�|����e�	+טCtem껽�N8�~zw�G�^��Q��;�A��r��ݡ2��M1F��Շ�x��l����>A�OՎ<��od�����d��k�!8�>1����pg�U9�4Ց�'��n��\�d��3yJ�����Ցq�� O'ƥLq|w����f�q��D..9z�����Qd�r;��+p9��^������i��a;�Q$���fe�!��ݤ�R+��1ߏP/���k�s|���
� ���W��#�J^o�<���>��Gƿ�w��d~1����%�w)�㎂�F�R�8��	�>�U��z&�T���ΤY��C54�� ���PK
    +Q�HK]E:�
  �    org/bridj/cpp/CPPType.class  �      �
      �Wk|S���\�4M���B�J�R��ҖNDت-e��REN��L���\�_�6��.��m:����&-�����.��}���e_�m�2��s��6��Cs��s���>=������4������t�wGC4�jX�n��=)�MC�}�����=;�h���3
�i�/��uzZ0�F:v��k�;5x-YK�A�=���r�2�?8`$������YCirW�H�F��3����.�ȗ5Rq=k���9�5�~���%��e[5���I�L�E�-ޤ�^�x��a����6����dU���odE�ZRWLΌ���t<�2�7JE^�^S�|����V�Mg�����O*D�������+�i}O{,C(�E�um&�"�F����*\i�U�b
�0fzo/!XWĂ-^,AC�qe�,�6/q�/e�Ie���/��u��2\ ��P�AK5�����FIu��j	�6�B�'��2Sd[)�b
1��d��Ov{U\�d���(|'��=�ޅ5,]�M��P���9R�*�<�
.��鋥3Ye����d�����F��U'Ffe�W����e�!�-�i�/���Kٛ��#��P���mF^���F�/O�S�2z�ٴ����T�/����(u���dzJ�6dӤ/��n���K�laI���X6�$:l��F�,,p���F��u�ջ�FJ�]���:U�Ń�x��vA��>Ae\p��X��3�Ūp8����X"��DO��D��{���YZ�>��9@j<����j8��,@ۋ8<��)���tSRb�5ʂz6����Y�GX�Ե��sP8w�<�M��ͤd�&���u�y�t-���t�\�TW�уm��=`��d�~��Va�2H�dvu'�o>O���N3A)wQ�7���6Mw�zJ���v�<�-�o�����H4l�>����%�2A�t�K�7��1��.��^|ǃ}���N=>h�XvO���q_���DQ�;Uj����?�G��f�1��q-kыK&��'�q���Aџ��Ռ朔Ȝ�a<,����c��D&�'��3��#O��k��$#r�=.�5��y�s�	�'~O	Jv�a����=�$��<�%��~�͝jfKH��ۋ����C�<��b��7=�c"�{KR֢R�_lԪ��y��o�x2aL�����&<h�Q�h��,f��N���1X����2���u��8fy�(to�3�W%{��W��u/N�<���^��<�-��>f3�A�=�F��x�{�A�M�lJ�ͪSw�?I��3�#���|g��S/vK�HF��&=�{��F�a���������<�<��Q�.<��騱��_��0�2f�,�I�'Ӧ�z�/gN~+p��q����;'
�aN(|�P�qx�/�1G�AT�Bϡ���69�ϒچ����D���V�QS+�iS+�j�'\ϣ}�
r���/#��p&Vb1.V6-�l��v~�!-Ù�A�<�ѭ�hj%zlJ�Gi^�?\sF��In'���p�G�����]�cX�ao����Pmc�#�8��~�	8&>�smؼ׮�|�q$r�kxQN��0��hW�-�� �-t������bp��З�ыxƊ�r:���������Ŗ����Ք�Zԡ�z�Yu�q.���k:u����cs���6��Gx�.���*��P���Y�f�;����n��f�`�G��:|�R7`eh��O����
��a����0<�Ͳv�R&ɪ����fa6�*���J��+y��7Wq���r���R��<m<�m]G��5���E���H��\G�KF�˷���Fq�n~i�5�ݭ*�Vd%v�֔��~j�-��K{35���������b*���f4��h�d�,Eu5͈3�	~9К�ت�ֶ��)�;�4vD�b���-3ط6l�b�c[g��Q|o��Y�<�a�@C�3�4ˢ$�_V�/!��\�en��_2�Gs^�+~�8�#��G��[���Ҁ��nl�<�}�xh?�JG�)W`i*�%���ǆpNN�yOr�H8���Җ�nˡ����n��fqn��U?��#�u�\c8P��dI�YVg)�G�����~�dM�%�>ee�\��9rؘ�� ��N����c�/��8�牉�8�#�RB�L�Jq�ʮ�s��Ӥ?LzI��א2��a�gY�;I����z�%�u�}=���:��5����߂��1��+��ĝ�K�sܠ99�H��0{>��26��Q�l5-�^������_����K��"�S��Ә���E�|1��1�Ӎ�ů'��� 9X"�yigM,�7F�~�:��j�rk�}�Ho����Z�5��b����G��'=y��I��m�Z���h�e��y����b�|fx�����>ʧhg�1Ҍ�B<�sN��WS�<\��y����-���d蘔KhHv��Q�&�w��#��G��I-�iv�gh�8��?���d�6kv: /s2|��Qؔ��l���u(!����>�X�U��WFڗ9�v����;�Q#;����9��F��IHݬ��U�z�$�bx2��'ջʱ�u�U<0��懋V���2�c9��#��Q�(��ˌ���8�7�8��؈�a���|�ޢd��ge�S1}VKj73;l"&]����氉��f�����X�h��5�XP� ���������mj5H|�hU2�������-77��1��)���E����>Q��n�6�ߡ����]����!����s��m�j#�[�WN��O�^�PK
    +Q�HA2R6'  �    org/bridj/cpp/com/CLSID.class  �      '      �Q�NA���
�@�F��ōgO0� Kv�iX:�e�,	���𣌽��KMMwUuz�����NΒ4rG�O�p6s�d�6�A��@T'j��X���F
����妪�I��:1��uP(�Sn3��Uw��'K&c�ť�$P�G:Hb����þ����w���Ҙ��%R�Y�_o�c��X���
�e��vzm��*M�Hؔ�/P�i�
	l�MĦr�,Ґu�˝�^bJ�z�G1m�l^ȡ N�����p�F5>�c�5%B�qi?��"O8�a���PK
    +Q�H�@�z�  �	  *  org/bridj/cpp/com/COMCallableWrapper.class  �	      �      �V[S�V�c|�
�Ҥm
%��M[��s�f�x0C��<q0�B�Hrڴ��K2��C@~S�����.�ӌ�G�{v��v������/"��j��\�U>���Ӳ�ye�=+�vwj�m�6����1F�/z��V��y�!������S���V�йu��hT��;�2�wtF7{n�X�h������b�Q�r��pL�hl[P(ۆ�*��r3|�hp�r���h�xq�t�H+�
4L�yJ�'*Е�h�Q:<�T��Oߐ����`��n�qV�]��rB�%�t=�Xҵ����H��u�h<���[�o*��E��$S���7L�T��2ӑ�6Eެ���CL(�M��%���;�ݟq&��T���3��J`[8�$w��!�1L��>~��/���c�<Qi=9��Q�v�n	���m;dt�?���^����_M��α�(� ��0+뵫~k�Gg�0��/<�N�c��k?��x������bR�I�bQs�Z4�t[��g��̟��G򞻦a�����ba4�m9��ǯ,��vC6��kZ-��>�?�����HI-M�(���I7$aX���%��1w��'����[��GJx�n�7��%Ƣ�;�k�<���xs2|�J�: y�F�އ�������46��������X'���DR�~�<L�E`ߡ-�:E����C�S���xH�Jd��4�F�%-�>����tCk�%���f�;@cB��s%��,��A��L+��#h_ќ"�Z�<��"S��H�bj��FD�6��$$�HQYw e�T���t�U^��B+�|�G.ő���SU�T������g��狙W�:�|#J���5MR+��{ �u�|�R�B���W)uh��)?F'�<�n�eTĺ��
~ߪ��1�c�2(!�3�_�(�PK
    +Q�H|cޠ  �  &  org/bridj/cpp/com/COMRuntime$1$1.class  �      �      ���J1��ص[�Uk=��V�
��o��P<�o��M�&ew��[y!�>�O"�3�� (^��d'��I&����������^5����^�Z^���#��R�d�1d����{'�&)���0�w��H3�B�D��v8�hq���"�>�t�qa�NY��!���1,��^��ۇ1��z=�ar�.ʰ���\	���1�s��F�n�j�mL0�v�ؘb,���b��ч��,��j�UT�;	�=���"$?<��8��o'BI��s�:Q����� T���#�4T���PJ�C?�y�<�¢�e��5���`���m�ZG���d�1ro44����b��y����qä҄-M'��0�7����:�H��f�a�VK&��&f��@^�b6�Ș<_PK
    +Q�H��S�  �  $  org/bridj/cpp/com/COMRuntime$1.class  �      �      �R]KA=�O�n��ok[[6����CPX���8�Ʉ͌���W�O�������݉��ā;w8��3g.s����-�3�צ뷍��������o}KU"bm������܏����=#x��C�<���}&ۻ��/��(0L>H�Xˣ�/�̰2�`f��PڑJ&�y��r1�Ao
IOƤ�-C��LA�ţT0�x���c�h�`ȓ?��C�;ꁋi�8�,!�m�j/ȼ�c!+,2�z��z���2	4t���� [�Hގ�i��(�R���-�=R9�]œ���9ѩ	Ł��}F:��{$����S��iD<�E�M�hV��Q��@߂N>eF����l����$�(�P�,r����7�!o�j%��K,�����|"T}$�X�4�$��2��ds	��T�(j���1��PK
    +Q�H�n�&J    $  org/bridj/cpp/com/COMRuntime$2.class        J      ��mo�P������:67d8�9Q7��$�˔�d"���ܱ.�%���4�!��e<-T@m�{O�=�w��������;�'�6m��6�u��ݮ���T9۷\�#2y	DxY�t*U�����8�.���^�����Q�����ai���J{�6�i� �� ��n�TM�j���0Y��M��4���,ȈR��JP8ݘf��?����N�	#V̽4z�Cޗ�yAcE�2�#³���3ע�`k2BH��I�<��D:�(�"�t��\5�<K��S���U�4m]sE�u��{.:�sMȎK�چ�
�2���Qf,�= (���8�!�� ���F-���]����-�-AX)s��9��4E�k� �K��w���$'ݸ��\3ږ���ϊ��ck|;S�țRy�;^���.N_�kK7�a�υ{i�ʩe	�dj���a��@��Hx'��?I�a��c���l�3ֳ������{e}?�[�]l���slǘ z��a��<Z�{/B�~�z�|���J���������4y��~�Ǿ�N2��P�>�C�#�����<����nr|+��PK
    +Q�H�U��C  �  $  org/bridj/cpp/com/COMRuntime$3.class  �      C      ��mo�P������:67�pnsCe0��^i	163��a��;VRZR�q�J_��P��B�!��=�w�������9^0�8nWn�f�'��l8}Y��>�l����� �p�M���Hm^xվt�ͦRQ�9	H0�L��=��>s3� �a�˽ 4?P�t�+����'�����7�<%���i���2H�:M�����l���U��)+�]���	uZ[T,50U6mӫ0�,,v��-	���&�\����,ri$�!�f�[�#J�c����ۨ�e9��������{�P���1m�����'��X�{�p��4�����p�\��lt#2%�:NC�VKwM�m���+��6���ܝ�d�ݨ�Ɂ�0���\��˭W3=��{��Y�X^D��t��k��l�r��ݭq���0HU��j��!b����7�d��@V�>Y��!Y��7 K߰U,���������b�݀X";E�3$�������b�+�J���3}�Ϡ�(OP �Q�e���dM���,�rLI�Vr��pBk�&�L�[@�Nb��������ĿPK
    +Q�H���  O  $  org/bridj/cpp/com/COMRuntime$4.class  O      �      }RMo�@}�|81.mSHiiK��V� qK�KԢTFm���Y��:�h� �gqq���N����3�og޼����� |@�a/�C/�r0��ċ���	zS�ɱh|���F�+�b��^�D��(0l�W~I�ʄn\�X�Th%��{�w��a�^6*�<���g��'z�p�<�Zu�vkm�p��h^l�0T��1�����	C���Xú�"j��Z����{i3�z��Po.���/8�O}j�g6�1�t�+��ЬgZ��t���lBċ�Ǉ'�{cIC��I$���
�>ג���2���/��<�B�"���f����*�M5�[KF3�t�e2Ց8�9����$�j��u2`p�J	݉y���aтi���Yth�tۧ�#�ȗ�c�[����;�Oɿ�S6���l��e�������B^\����&��J}��.�(2Ďɶ�(Z�h���M�xK��*�5)�f�����_PK
    +Q�H׉k�V  T  $  org/bridj/cpp/com/COMRuntime$5.class  T      V      }�]O�VƟ!����h���躦��]�4����%&�c�f������r�� ��0i�v�������BW��4>@��&�����'#M�D�<����$&'��}�
�8�f8�zk�UϪn$�����n&R�\��ԭMS���1�7�m=a��Z���a�Z����|��������AU������ӷTV�a��UV+�R:��c�dگ��X�-�c���c��r�X��L���<׋@a���7w��C۶n7�=���J����
�莡=
��"�>�����\�\Lj��S�]'����!�zU��m�2
q��|�!F�-��异3b�Y�i�L2�)8'�y�Vҙq�0����\�5��PpQ���H},���Д�+��jJ���s�i�)�D�O���.�g���)�-z~R�����¥���������\���!� D}���Ea��]�\�*���\Q���K!Kt���t"��>3��[5z����ݳ�U�����w�r�|cs���&Vv�a�[��c�n�r�rf}ݭ2(�1����jf->D�&L?2�秈7�:(+@�W�P�~��W�Ş���7��� ���ak�Äm^ �8F��%�����#����Os�|�s,�Y��������cι+�/8��q��ȹ'�2�^�����}8�N�c(G0�i�$1G�FeJ� �b5�:����;�?R>�O���!�)�3��w�=��?)��Q�o�C�������Y��R��!6L��+l�L_�.}�~JKt�mF��l�lU�����@���=�mO�}�d{{�XX�>�T٦�;�j��ջD!��+�0"t]�W��8���PK
    +Q�H�W��  �  )  org/bridj/cpp/com/COMRuntime$COINIT.class  �            }��N�@�ϥ��ڪ�h�Nג>�I�4�M\���Ph���\� >�q��)+7w��ws�����0��(��L�S5�nըب�c�M^'��Aw̹�+ �$?B5���8�t���X ���@&��T���h��m6���i3dvxC�0=�د�o�y�@�>8���'���f����ӽcF�,���v�7�{��^�U��2̚�0������$�04�<.�,����%tE*n�ǀ���p�y����9OZ|����y�)����'�PK
    +Q�H�yÜ  7  4  org/bridj/cpp/com/COMRuntime$VARIANTTypeInfo$1.class  7            �TQoA����h)U�X��+R@��o6M�		-�ޏc�K�]�w��g�`l|�����W�*Մ������of����/_�񊡦��h1��t��j�6;'ݙ�Ą;�F��8��.��%�+�n�1d���<9r;�1�#	��5�;%dĵ���B�-�2�_��Cu��R��CX���_0��]n3�~�cX��E��i�e�!䡐":b������3�b#��eH��>���$�3$� ���8�:	��UW������E�N��1��ċ��m1О����!����d�$R�/�VO�c�1�2�r��&K-��386na��M	�?,���x�����I��|/���3��-$?�M\�#�?�h*���I/�i�n��H0����L��������P��	��Րfђ��f��!�C7��`٬�J��Vh�I�2y�io"v��	�ʟ��c�S!��:�
���Z3�K�!�)�0tigR�K�^�h��������{�}�~��DJ�U�:���`�"j��xbϢ� ��4ٗ�
t����k#�v�k�PK
    +Q�H*mՒ  K
  2  org/bridj/cpp/com/COMRuntime$VARIANTTypeInfo.class  K
      �      �U�SW���������hi�����M��RbZZ�T������k�]fY�ط�����m�D3�L���Q���, �d�{�{���w�������y	 �2Ìe�*[/�+Z��hVII�V׫���xt3��I�ml�y�ܱ$0�d�钮��&K�v@%��d��,���ߌ?��>T[|�9J���Q����+�� 3\h�ܳt��vt�\�p[B�a��\�;��C�=;	��t�Y�k�k,{z`*�PT�Л�[f�^Q/2�m�>gO�D�.w�z3]��[�M�Yf���n:��F�����͔p�A�ꠅdVtM1TsW����5Gٻ�pE���DN���~WF�0�✠x��'j@�~;4YDW�gΰЉL]���2��)!��0�3#��T�U+�m�>�z�j��e(H�ʵgr��[��%ø��}�j��:��Y�%�>`�Mut�n�%�qSF ��?��^Sv�(M�uKbIF?nS�TM�R�<���Tu�tMu�Vƌ@�Q��z0Q�����b�ڎ�ˮ���URE��z�V�	i�Цj�I��0�!M|we���t�u�⨦FJ��Eg4���]��ΈK�!��.	p��J��E���)�iPu`����$�7�	v�k�&ʹ [��|�\�l�Wi�,�)a#�u�E�7O܏�l��r �|ɳ��c�4�#���kC\`+��@\�o��O���i��+�͋�ۙwT�Zq��vEpv�_i�H�d����h�n�!gu�V�Tභ3�jF��;������kR8[䭪�񻺰
gL��.K^�%姿�^��xFĈ�u@Ld���G�"=��W>� Fc�g��GƏ0{��V��=õ't���ar!CLa��}�F�l~v���&1�&��(���d�a�1Ύ�����_ze��bO)�S|p�EZ�by�'�⣾��D<>{��"�ߨAy��[�����Y7�$V�F�qPf_�=ⵝ{�#�,�y6�8��	9�E������[�K`����՟�*�64��}��`�aл�����k�6��7����!�N��Al�A����J��=jB.���!�kv,V;j��<X���W�~pKv<T *� Ӯ=0	b�1$������Y��a/Jn�^�����IWaʉf*j�34���T����PK
    +Q�H���!  �L  "  org/bridj/cpp/com/COMRuntime.class  �L      !      �\	|[����g[��Ď�˹P��8vr`BBd[N�Ȗc�vG��XD�\I�A-Pzp(��R -���|i�@[Bi�Z��\���������{��lŁ����ޛ����ٹvߓ����'�X�m%1%۲�+�9gAw���h߂:oc�@$�Z���ݢ��9M�HgZ�?'�-@b�'�!�,���b����$��A\����E�[|�r��R�AOҡ.�1�qLb�/�3��-�DO] &1m�iW�l�I��M����l��w�ݑ�Q�(�2� I�8"�:����2���$[b��f�EL<^�E1�xmZ�'d���{m����4�s7�	kF'��XEg�q���ltu.��`�,�D���e31v�$N����lI�$a7cH�?ǡm��X=|�S��6�Q[��,�nc'��T�,Oo��"�`,b��^�XLb̰q2	[�\p8��`8�s�X�'�����:�M�-޺N�����B���˸l�gS����DI�� z�uN�їIy�U.�k�j͌��j��]����	9GԻ�RK�]U����_5�������/^���M��:o��������:�A����d��O4uk�����������'tW������!2�������bW��
�R�X��)N��]����$LC6�@�zW������M~������T�����nsb%/�u�����Q͒�FVn4~��0�u�&H_��Q���Y��h���/4/R�-5��5'&d�e�d�<_�w�NЗ��=��V��v��N�������#�R.P 5y��W����ML,a;�*������qot�3��.���&׆fW��q��I�m�y&��$�\��V�����ҡ�R�	=�Mm`V�lY͸vհ	)��jipֹ��T�u$#��˰z�U�	bUk�-~&õ
\�>�'1ĺ:��W�jr����I3�T�G��w4��d�g0g��������!b��4i�6�3R�5�Ζg���_�R�Q�
���P�jN1,�b<���5:�uk�	�3���]]��4b�ǥ�.�4��<�vF����i]�ɤZ��+ŭ��V۱���e|)�)���έfb�0lv�8������R䴂�24���u���6:���ֆW���.<�i�0i8�0� Ci�2����y�	%B�p�\�<\�-"[�{c�@�'�����MYaB{��	v'�����/�D�Uj"�Ċ���y9�RV�X��@	�\�>t��=�a�+B�{%	�rN�]��m�3��N��H���
����u�E�J<�t#�5Wz����9P��l��4��`,؍{0��hF��X�Z7�(R�6'bhn77�$+�r[0i��L��`,�1�=�<3�1q׎�`�^/�:h�w�c͂=��*~+��h����G�cPnc�/����{�h��t�؎��ͷ�'��,q�c{ ��p�b����ӭ�$f�YQ��AGO4W�B��`,�pl�E��a��U<�q��;�u���!t��gH�����P ��D �;G �t$z	�n[���AVs����`�6����	:���S�m�C��v�H���🡚��{�`z�&^b��b�9R�;��	:�9��W0�@0;��k!�����ůū<�o0�Ć�q�ב$Q���S9���^��m� O���nK0�vד�e���
����pO�����6�FpF��@B��Kr���MdzA𿊿��;���)
��)��}A�x�g���J.G��#L8pQ&`����Hwvao����l �ne�ι@�u`�<ʷ��-������C���V�s̰�B�PO�ڤG�����hB����.�b��<W`�&Cq�ξ�hثbD |�y����0,wAc0��Y>��p����1ۡ�)��G�-�.P��˙R,T�5Ü�ڤ�_�4���hM%Q	n��#�dZk�����vu�0�}S4���d�$M'�j8ߏ7��N�� *�4�S��Y��T�4�Con�96QCUv%�̽��ş���v�=q��N⠋���f*�ł[Bq0A�Ax�E�{�B}��rZ�\�x����C=�����lW�Y��TnVCː~�Xi��f����x��>]oll'�.o-�N�yt����y��`��8�M����`� ���!�ڮ��c;Bn$�������>�ᝰ�b�׉ж�n"�VF�sc���V��k���C�BkAb���VyF���f'52�&q��8�'�?���*����Q�J���Ѐ�>�%�J�W��`�z�I5L'_,i?x���-�*� ����vg"���p�"�T�hy������y��+G��T�B�$]�"c]s����Q�����D��l@���g�m��f����K���̩)�α�ɴ5�8�6НHI�g��N��	�-/��cq���XXA*����
P(�(���t;�~��v�|���,t|;��P�|��4G��(u
�,���t�F8ْ�U��N���p���Tq�rjAGG8����Qv�ZD�-��D� �٬�d��@W�(t�W�sTG��%���(�3TO��pi*�3�,��w�Yk���
]FW�j	x�3�ݼ9�a`�9��*�����:bX�.��h,��/w��t=��!�UF1��	du����f�����Z��ݱP��Zt ��M����\6o�ff�l���"}\V=1�.W����~��e����<�؜�ϬS[p7}�&*�;���%�u�촗9��X�Ӯ��F�o֩jC8���'a9��i��̫t���`2&��i����Ɓ���<��Ydhv���+���N��ڃ�>K<e,M#Kn[a�QQ�>��Z��(��h=D����}r[�K��cG�8��+r��֠R��c�C!�I!��գ�sO!rx�b>��k4;=I?eE���#���feM�U�FRk�=���+ٟ����i��r�_��>o���	��"i�w�v�����H��2�����+���@���3L�飢�x�~�c��DE�o{(���� �
Ÿ�+���`=����:��P����ӫB�����<�HՉ(�#Q��3�ӟ�/��-����g��;����_9g�����m��;�	��?������V�|WG�����1�{_�a�����)FcB
��<Ƅ�@�X���pB�
u��q=]z;������uT��*A 7U��(*��E�B���]���V���s-��NлN�];Q���$3 ̱=�Lm��T����P�Tت�K���=fd���-���'����'T��ZZ��,9�&g�JH0�릊��\Y�u���	���6�˪~���,�����"�jY�e��Yj�MÖ`�"OV����AR�N���:0t���23��pI�]_�.��p�+��Ƭi�렚���2�W}���N�3oWք�� &��'�`f����&�Hl�
t�P����#�]SV5\���"�y�^o�S��\/9��U��6,y��ߒ}.=��,�l��b�ܨ����ܢG��~��Yy�<���l�3��H|��k���c��+s�!7�X��*��| �Nd����;Q��'�F,5��dא�J#��x){l�%�s�DԱ���[l2�g�'K�K�e9"Vw��j�{!GP(~�¤MM�'��j�����s�5|8���HD�����f,%��6��N	�WR����χ͔L����mv�
��;�w̬�3�D��'�y�M~��e��l��8�,ֺc�Z��ܻvD�民�j>N���f�]~N%K�y��dZ��b>��%v��v�:7���/!�!a?���wG�n�?Y��K�e��2-��+u��
O#�B]�@�@wڅ��8F\������.��{� ׈sx6�ބ���?|�d�瓖�Ǟ�-��,խ�T��6]��1�.�C�=�^�?�dij�k�8�,�]�4-X�o��`�f���g/r���,N�M�:y��-_Q�
���I���<z�mt���G�ϖ�����X��_���
!��DV������6yHAv����.�u�}>��W���d��O�P>���~�������*ɬ�,���|���8k�7����+n��O<�s����n���q��M>&�D6��Y	?ӕ���_0��g�V���l!���B8�f��!�,4�~��v����/�,y�P����_�W
a�踞��p~��^c�M�����*�%���Vu�I�[e�?���h��@�)�Y��ql(��+���l�����s@=|Leq�9��ۼIc��O ��U+�C��#9�	����[��P<�h��T��7~�mY�]���{c��U����y�R�w~d!?�����Yz�A�$�t��=B�\]ih�`�|�8Γ�3�at�3�c�-��;	�c�k��&fq�-J��h�Ns>b�G~׊��wmj��i/�R$O�*'���f�r4�h����gv�d-m�6��m�G���i�x)&�V0�4���4��6UO���>���(�R����ۢ�@|+4�^����J��k3�m�t�"��@»YW�^i����@��Q`'1�����kG�g�*؟V���1��]�#[&�6Ϧ����6�C)����ueM���
��S/`C��E��6p��h�� ԣص��)d�Vc$��@$��n(�?ȏ"m��n���h=޳�܅q�	SNSFI]�~p׬�>�X��q�ٵӴ�ln���w��_IL?.3n�IeEw�x�h|O0�{ҵ�/H@m�=�xGî��$A8����Y47����"=��h�����0�q�E��Қz8kך��W[oS�.Fa��R%u���M%b��O]�'�񗟕� ����,��"����.����e�:"qg�ؐ�i�G���=���B��f��|�_n*7��-a*�w;�$3�i�(}����h|��� ���½l�	{�������r>봥�Ӑb��;�z�]�����͛��F<3{Ĭ}���ym��s�G{eF2���7�`������q������h��kW�-���eδ���\�5��c0˙�����ĺ�!�2�;	Ɣ}�b����8M���b� ��o�+x�	>�*�\k�� כ`��������1����L�p�	^��� �Mp+�6�x�	� ����L|�Mp'�M&8 ��w�1�A��M���&8��p�����(��!��)7�	�&x��&x��&�\��6��|�	>�gM�.������	��E&�b�_0�� ��	��/�� ��_�r|�+M�W_e��|�	��kM�u�w����`�o|�	��7��[ ��
�&�6����; �1���-|'�L�݀�m��#����V�+&�}�4}�D>V��dA��5(m�����_u@���j����H�]qHm�m���MM�B~uMhZ����m���W��d�1ę��k��~�a??4���@>q��4G�úXT�~n#đIw�W#nc>��	\c�;	\?ÿ���Ͽm��
�5��o7p��_b�z6�����,|��t���x���{2}������g�w?O��2}�B��x��x�������]R��IC4zD��E�5:_��^������!����Mµ�Ä��}��CQȯ�/����]U�VR��x�S}T,1�.a��|�_U�}���'�@����J��:c��M-��TD^;+=	��(U��q�{�~y�)� ���֣!�M���ʨ�%�b���+��D.�)�:C�"�
"��y�0�_@�E�x	�ꕴ�yTJe�kԠ'�yw�WQI�~�w4�ơ����x��v�
��mI���F&�@Xć�q90�Q�~�nUU�433G}�M3+0�LI@R���j4Ø�&5�t���t� ���F�3��z�,˛G%�����q���[�@4#�@e�X�	ը5Y��yIZ��ӌ�����Ҫ�I�[VP^pT��%.#�]yAu��Gh�2K�e���������:���:���|��-��]V��Px�)EV��_w�.���i�\�
 y��֓�8OL&?�Aɘ.�+����w�F��P��t&�4���]�R��ѹ������mHs+Ls;#��4���m�2(�'*B�}J�HL�ö́��S�8Fۅз&��G�T>l9��M�g]ox����Yw�A1��� u�~@��[,,�`��N�B�Ũ�brGU�
�-��]��ѽ����C�}m�����b��P?�;�L�r1�V��41���2r�zj4����Q�./��*8|�5�⃴Ã�pn}&I�[Ӻ��q�8���=����J+�&�+%%���K�����tmU��Ğ�^��}SU���$��6��z��[]b��颪��)������M�W&���%�����KQ
- N嬚��6Do$3q�����b(K�z�-�ǲ���)��n�:S삡|�o�&Cq������(�'@Mwy�H�4���[9�����̪U���tH%�R��H61���`S�{�AL*�G�SP�h3Vs�!@�}�~`�Y�~*�Y ���y��?"���I{UFO��|����b�FB�b%�f�e��QCc�P[!TB�a:C� �z��0"l=y�1YZy�i�P}�I�Þև%�IO�3Y��a�8�N@�X���>��"���A��� �������C��C�G��%����>z#��$�}��'�o��TJᢆ�xB(\��l|��~�3�Ϲj�υ�\�������0���׿��C|I�_��e�"��_c�L�%�x�-�)���U���{yC�F.J�e�4��g��م�%����
�o�s�8qP���ʅ|]2(O��Ay:_O�-,y{@e-��r_������}���K{�@:f�nċ��\&{��!C����g����^���L��0�@�mR��c��61�. �sh�y��t���.�ӗ�/��_	�F|����n*7�Ct�x1�Q�]<~���зi�Kkh?5�����&�c?=H;����/��t)="����p�ka����U��S�s�j)��W�;��Sw������g�;�%g�]rv�%g��T+�$��t��c�l�%�V�|����!O����视snF��K^�{��<�![�U��������{���d�n1	�/1����Iʯ\��W��%��e�i�ɫt*]��_K���{�mt��o4��Oʛ�� >�L�x�A����JʻA��5:���&)�%�~oq}֘r}R&�A?�!]�Ԙ����A���b
�?`*���l�aНH�5��)��i^R�dY^yޠ����|])O�Rě��e��vQT��O>w�(�r��G������*����7�P��g�_*�����C�y���_f�_V�_3~���W�Ɵ����7
�:�'�֔竚���ꠠ*?;��|��5��,����Ǝ�L��qܪL,�U�����_�W�ݚ��K�]���)}�?}�h��7黿����;;Y�߸"Ć��ߑ�\�+���1�-:�Gr�������F�`yE,��<y��9QF���b:=/�b)����K��^��LzEl�_��{U�l��o�������j�w�n�=���A����Q<Ao���O�5luߤb/�.Y�=��/H�>��4�>�J)i��h�̣f�Od�J�K+풅t���u��n�v�Q4(G�ò���%��C��RzK�ѻr�/' c���r�\)��<��|�H�s�s�e6KzR��C�A�'b+�{�/��u�\.cK(���<�U����ݾG��˴|�B;�.�t9��-G{5Ld/�!zM�#s��(��U+TQl��ZEb�fӊ�p>MŦ٢H�c�\��e�p�y�d�@jvm�!e�0�iUG��{�Y�ўjaăZ)6=�C+�i�/�E�fǝ>�xeA���%�@ֈ��1E.E�+��a�+�?���I��zP�2t�[�.����	Y�]�L3�J�
#<o�L�d�c(� ���
����5mP�Y;�����̃��ojs��iImn�6��Jm���������%�Vx�vJy��Bp��T;U	�^	�5��2�4Q�Tʻ�|�֫	�4Se/+�N$�:1J�#O��B�E���lM�kL��Ī-�V��2l�RU=7��ʜo9t��4th�j�:5�E��dh�ѷ\���}��KeR[s�Q��'wj��E���rPL�R|����n_?sh%(�ƫ��W���r�|�\c0�b�]bc�F�`�R�+(ԈV���&ש�1]�@�
(k6�5wU����<\��bѪr�[�Sp=�e����h��i�����v�0.� Vc��PK
    +Q�Hc��x�  �    org/bridj/cpp/com/CY.class  �      �      u�Qo�P����
]��t*��Ƹ��81K �K���ɔr����Y�}�%������C�m	8p���s���{�����/ O�a=��N?��㟜8~8v��:Cu^9��ď�#��:4�}�d�z����'��>���C��N
��h��+{B���ִz&J0�ʐ�?�	ɻ��3�2~���u6�-��CN���A:�-ױ^B�庎Ms�c7��ɰ�\eiu���n��[�f׺����f�rfWm�6
z��Ѭ�t�O;�m�DH���ASܧD;ж+n�{Aϋ���eʮ��]2��h��M�'&��R���P�捣0�|~ �m���2�2�HdҗC��/�?`~� �&Y3K�
���謤�gd˸F�T�.�4k��Q��sl�-�%��dW)^��wPI��)�-��G73d�����J^�3��ʸK�V*�j{�_.K��v�#�&%Q����c�l_��K�}��E�Ҟ�LHͦ�(�PK
    +Q�HH��  -
    org/bridj/cpp/com/DECIMAL.class  -
      �      ��[WU��Ʌ�0�����b�
D%�bE)m	�vb
�p�N'�,:f�Ʉ�/���]���k���C���$�&<d��?�����sf���� \E]`�qw�Uת��kO��k�~����?X*� ƎW<�U�֪{f�K!.�u'�������\ö��-۳�����h���X>z<p˲-�@|fvK� 2$0$��[M����z�ٺ�4���*�}F�Yf��'1b�s�HK_[���"�����)\�5��c�����ř�R'�}��aod�:&.�Tf#1��'�'OW�Ȕ.aJJ�) �<�a���ɱ��`2C�w�͚�0UB��V#K�'�<JAC��~�K�B4��<!AR�$y|(������TF)
��4�$�M�֮-����^��0ߙ�։���k�R��xH�H��g�/]�],I+	�GC5��F0�q���gd�i]�<DT�Q�e�����$	�}*;��J����T����tL8��$��-��$C���!CIv^Ŧd���e�γ6Zv��[�kՆ�!/#e�6W[�U��Vƻ_�-�i��dێgx�c���T��[�Ij��L�|��*�c~%x��<G�1����p��Z��a����o@U��:B��Z|qU����X.����>�L@aU^�x��/�cTINv%�t��;�m\ν쉎u�uE����zC���ns�l��۸�E�ˉrj:G�w�'����=�t@�H�V�1�A���gP��U�s�$��Zd�j[�L�q|l��׏�2�8:��)6Y�?%��2��o�%�A�o�>�;[d�ix��3���Ia�����@��3��o���,�f0@��#3X�~��S�n�E����Dg��F�YY�� ��Ƌ���7�PIn�2H"�� 5��W���`7��_�-����2���տߞz��3���F��yWSk��F�-UC�PK
    +Q�H ��  �    org/bridj/cpp/com/GUID.class  �            �SkS�@=�}b-򴢢hj#/� ���
�A���͔`I0M��?�g�:��?��nMC!3ٛܽ{�9gw������u�*���+������'�~��9�4es����� �!^�ݕd���Y��i�f�{J�� �
C�����tϼ����7�ފ"�p>D|�Zg.����ٔ'��"À�����*9/��G���Ĉ�(n�?�:�b�TS�L��V��eJNL�Q��f�H0$Rb�b���y�ыAE��m��wiYʷǕ��S�j�h�T<�m��l��|��^ ���U$HQd��7{�%H]$���a����O9.m�l�'"$�8�,��1��{��)^�l��d��i�S�)��U�T�\�X2�0�G�	rl:�1��^c��v1ǥQy���$#�W����\ےU.ՔM>P���)덽�bؙ�l�u�K���������V5�lT�t8_�O��ZUX>4��IKz�(++jM��䳤F�н�q�����?���`��1�J��(���X�c�NU|�4�V6�������[G�p��lqz"�,�Q�@,=|y2��X��t�5g����z�j��(.v���>�mɯ���3���S��<�v��IE�2I�\=�5��rD'���u��G,'�z��T�u��-��u�̓��=p�K�b�2�x࿒���,Hw��z0� ���vg�8^�{0��'|�TT(���Ń�&V�/���Z5E��}-r�_�ֈ�Mz���2���<PF�?PK
    +Q�HZ3��  2  %  org/bridj/cpp/com/IClassFactory.class  2      �      �T�NQ]�ޤT*� (b/��"(-5ZB2I#��N��:0�4�i��/�� ����G���Mk�I��龮������� +x�0m�U�b�G�V�)�u��E����\s,�4�0���ylZ�����#��c�.Q�V�!��FC0�-{�ʢ��(^ݼgu�!��M�)0R�r��F� C����f�jD%����Pͺ�M�j�S-Qo,�t���7UZmo���R�m���\�xC�$9PnV�-Q��F�	��j��s�n�}v)b�@�qn���+�{��B��F��8�dg����ۆ��'"�{�}U84��d�$��ǝ(�0C� #�H*�Rx�r$4��<�CYe����.w������P[�)�<�L)9�Ӛhg׍�����#-�1lw���D�-0܅P���<0Z�h�Ҏ��ݔ	�ާU����!!O��en�b�)���n���IEؾ&z�3��z��N�&×.[���nXz}�?8�??�������u��iZ��2�rnm��,�~syu�g�}�&�&Il�[[ۺ!0K��� I&?$��?�NFg(���t��ɘ��mҹN���Y��ў#��n�n�rt��6D^	��{#��u>S]Y>���N�e/0�p����'��]]"�=G��3��@2^�D�2X��a�`��˒�X�ov y�'I�ye���H���Bn3a?D�G	�6�&6��'xJQ��:�fV�Xp]B�&�F��[�PK
    +Q�H0��    ,  org/bridj/cpp/com/IDispatch$DISPPARAMS.class        �      �R�N1=γ	��hJ)�<���ʂiB)M����X���'�x�_]!u��GU��Uɾ�s��������� ����85�74*yb2�D:���M��G7A���}�kXcx���Ʌ�6Ia�(2����yħ�a��UT����K���b(�O�P���%���WC��>/H��Snb�V�dnW/U�JC��ʵ�n�L"��S��Hɀa��ɫ���2�M���Pn138�@'/H�F�:�$�z'<p��0�wnbhv���|<��	��*�������\p�������9���ڪ��L���uj�U�&����%y	ױS0N����V9[�@ki��e2�>
t#�+S<tA4o�ʣ�z���wvhn<�X�
Տ4*3�"lb�X�f�]�Q]r��X�A��s��ׄ�{�ؤū�{jl-j| ���X�T���x��PK
    +Q�HT�W  �  +  org/bridj/cpp/com/IDispatch$EXCEPINFO.class  �            ��]o�0�����Y��Aac|6֖���M�PڊH�6����I��U�D���B���B��N�UE���9�y}�:�~��	 �ap��k�� I� ;^K�	7����m_y�K��ў�Y`.���EwE'#>����Z� r'�`�L*i��~*`�P�5%3�)���uyʠ<u�P�B=��:��ӑ"
���(E� ���H����xN�O��řP�Vỏ\�R�O�,0�$�%�@���XQͨR�������]J��)E�뿚�A�Re�/��w��l%7�%n��"D��˕-l<�x�XEsfG�����\K�G�3�YW*q��}�o#�י2r,�2���Tl85��Vzr���4rǋ|֥[u"��;���9Z��oRʞyH&�'�RB�OS��>������-������od2�X�a6p��Iy����	𻁫5������!&-J��?�'������v�]<E`o�����߽_b��\��}`��ˀ7,�>D�}^S��[W`�*T� PK
    +Q�H2�G�c    !  org/bridj/cpp/com/IDispatch.class        c      �S]oA=S�"���V��Z�6��!Ah�$H	T��@�0-̒��'�O&>��M�x
�d l�sg�s��9s�����3��Nͪ8��Ҫ�ZV�nZ<�ܖ�� Ú�Y_i��"�0?������30x��a�#mɰ�L&�&��}�������g�s���/��ϟ�b�;�hY^*����RQ���a�Hi��D9�,�1���^]�������ŏ�;�nI�/����R��`+�I�0���$��UV���� ��ȝP+q΍q|4I4Gh�uO/�)�)SV�kL�)��;��%�&/M�d2W/+=��}N9c9�*e�(Qi�3`X�)-��fE:7�PIմ����U��7i5��Y�5J��
�Z$�TS���(TZk���5�_�x�G�]��׍�R}�Lc���g��U�[@�(��b����p�I?�ASc��~"�d�r��������U~�d���<Q���r���iו.61E=�3�v��4>��;�����@��xAc���<$�E�v�
rL��K����w�l���9V��� >X'�cl �a�<ų`w�� ��[3xE6F3���0Gv�l�2�S\��PK
    +Q�H����$  �    org/bridj/cpp/com/IID.class  �      $      �Q�NA������
F���	gO0n",Y�iX:�e�,	���𣌽��KMMwUuz����@�F�Fr���L�����tݮ!P�����2��&3
����Ŷ��I��:1��:(
�8�&
\>�4�d�d�V��V���H�I��<�~��t׼R�-MY|�[�4"�����^LslĢB�<�q{�^��u�o0
�q'�|��u�W�Ȧ�Dl���Uҽ�y�3�K��I/�$��-�9���)� P�	�N��A���(��L���}.d��	�8ʠ���PK
    +Q�H�=�  
  #  org/bridj/cpp/com/IRecordInfo.class  
            ��[S�@��R�PJA���xAm�D�����0X.}�-�kYLw;i���ğ�3>��Q�gbLk��}HrN�s���ɷ�_��C�$0%��rh��Ri4���+�����"
���d����=�B����`�X;��o�ب�U='�nQ3�X,�ɛsɹO�XZ&Лa���"�T9��A7�6�X��tX��t0`̕�I`,���&5VS��	k�+ef����F�N@`�q�өfH���D�@*�oh(i�E Z�f�bU)F��թ�q�}������i��/��^}�*0�W	d:��2�(���$�z��N[��ô�-7�zA������[jc����6�LBm�����5Y�Vk�@�q��5�f"<�L�В��g�<����Ӧi[9�7'��pdKT4��L;�鞼�b����!5�4����5�2�y2$�Lz�^��;7Y��Y��a�saj&���®���0���V��=혬���S�B�5^S6NM�֎�l��9����%w��N����N�B����k��-gw�li�,�����B��b��m�O�A;��������}������/kB �S٦�]aZ`:�[Ѕ-N�K�y���u%�D6��g��m�ȳ�Q� $��T�[��=j��zf����!��n�*� p�p�Q� 0�����z��>�y���u�"L!p�d��47�9�F�����\���=��� �D �H#0�+�� � �9���BPX�2(9��|!^�%���eT����\)�&�� PK
    +Q�H��tz  �  !  org/bridj/cpp/com/ITypeInfo.class  �            mNMK�@}�6����*����4�/� �<h�}�����-����<	��(q�XO�e�̼�����/ ml�L��B59�l�f���o3��O�"�.1<�6���"��o?�� l{K&z7k.&�$��{�v��	n�E�G�P�TZ�W��ѱoc�*J�J���-��u���g1�E��`"�)���.�d��TL�V���}�c5�����Z�X���(�i?>������������E�vNbu����b���,lr�1�*�+�PK
    +Q�H�?�  �     org/bridj/cpp/com/IUnknown.class  �            �UmSW~n^X��WA�ڢM��ZS1�]^�b_7��.���J�	���t�ig:����s7��/ݙܻ9��=�9��}�ϟ����e��J]���.U*钳�֟ۿ�Ξ�A\<��/--�e��8��m�$+���N�{Wڞ����aդ����W�}K��x�aYܾ�">}����y2�����{�	�n�5n��6mA�_�o ��SC���a4�2e(pΨyβ��Q�?�B�#kڦ�'�kqb(�.
D��fU`�Uށ�-����DA	��{+]�K&�~�xˤ��Fђ뤭HW���V�~�c1��*�p|�@3R�sӴ�����W_�Ξ�J��8p�!|ʒ�����q$���3!�{�[��8ƕb���~V��n{��4J$H&$XrL�ɴ0%���X3]�fX�0����W�O��\�Q��eT��%|_S ���b�7�SGǗ���>�=Ү�5<`����s�WjQ�<�w��8���2�1��j�9�J؂ᙻr1��D�P�d��bz��|�"O��ήꙜҪ�����>׬C����9���RW� �3���T] �b�y�,U��Z֚ᚪ�W�@e
�-j;E����_K��.��I�t��[���\����m��Ѿ'����j��'�̪�8gl�� ʡә�BA.��>ݖ���uLrd�+N�-�9SQ�uۖ���U\c�E�sQ7���Qw!�u�Ks���W���*���1�˜7���-���G	?Aط��"t�������ɮ�!���$ �F��8j�C�猍w�u�zD}�?�P�G�\'����������&a�����{AK����� r��ԍ��}��#��}F���.�P:�ƽ �.Q���C���OM�����+��C�>y��G�F�M`؏.U_D��
X qư�g$��X!�'�U�u��{�m�/�K�����|J�|����l��	?�s��\�ӑl�X㞆�6�"��=T����_UZ��d��[��@)��p�_PK
    +Q�H��GT�  �
  5  org/bridj/cpp/com/OLEAutomationLibrary$CALLCONV.class  �
      �      �TYs�T��ǲ�$�N�ҽ�N�&i˖��8Mp�R�&�Vv�TA��,'t(P�G�}{��f��	����3���+'�6C��{�{�w��H��۟ ��C�qgל�K�^M�rb2�NV=�lx�cĝk�����Ljr"cx/3g�	˰gi�Z��%�����+c��3�jif�\-k���гE�0z7�<�Y�?aD����T��hR��C�]���RS#�]�hyFOe�:�3Dȭ��VreK%W��Q����
��ץ��ɞ���=W�i��B�Rl�!|0�̜M���ȧQPU���w_�� ��a�$]E˱IWg,^7~���Rѣ���_�^ �"��e�t��=;�F'�yR�Q�nF�vI�!ܧ"�C�m�I{��kT�!�6��4�����huo��i�Gy���{��k�O��+&�<�S�+��縜ėX�L+1��$�kM9�E��2T�x��B�����b�^Ϩ�x�c*�6��
�q'�PN�_v�rNNZol��+�_*��½*��bh[=1j��2���^_�-ْxR�(NS]���_v*TN�Ƌ� �uF��f^�I-Z������*�s
������g5D%���6mҹ��]C�t

:j4A�U�YC4tJ�R�UCC�$����ڨ�[��
zjhXC�D_�qH93T�֌i�&��Bɝ2
�F�hX9�5��ݜ���Һ!&�olӹ��:�U��G��N�-�FM.]��+>�Re�����h��ȶ��շQ߶��ݷ���m�o�}��-ݢ����*^wD��R�W��O�?�"����;��y�򾉽w��!��'�U�}ˈ�A���5zkr}8B��!�ǖޜ�4��3���u���7W8��r�cB;_q�A��B��X�A��q�u�A���K��B}?c��u�B>���M߻/���(��_1̰1����2ޠ2%��4@Ry"��e�,cl=�"�R����&��)�[ �������3��mL,!+��T��
u���?߸��0-�z>,!��%�鶄���6��į܌�k������+<��]�W���I|A�/E�~M�ףM�NpY=߰]χ�����)�%=OA�z�k�B��2]2h��^ח����Pс�i~>����f�#��ǘ�'x�R�?�W�K��K�C���[�*x[���ZE�p�PK
    +Q�H���   �  5  org/bridj/cpp/com/OLEAutomationLibrary$CUSTDATA.class  �             �U]SQ~�|����i��)��VI �E#�5�,�C��.-�3^�7�^�LC3]��QM�YV@�L�.�Ǿ�=���9����� ����b8�+{��B�.h�p:��ZY2MM)y]�g�;�l"��9���MC��t~_.N�&{m_ؗ$���#sb��u�Ȱ|A�bv�no{�ap]Q#�`9/����K�ReXL]�(��.�kU#!�	+2L��H�N*ri�2�RM���`�)�x��G1��
��a�$��{݉)���l��a"3L]8��ы���4n2�b�����l��f���q���202c�i��Y�#9-��|��P���Ŗ�B��7����ѭ�����e�����ba.�CR�Џ;#�NU�U��$ϖ��e=dxٝ�~QQ��G�$m�	ns�q(�y^�a��8�ڞLW4��RN�)_���#���ʯk弬[���j(e9�T
�TU3L��ڹ3JQ���Ny�^����VN~�Qr�4�ܚ������d��^��
w�+����KR�*W1C���/�O�=�JO�42��0�&6D��6���Q�Q�7l�Fk>��3X������Z�^ǭ�O� ��(6h>D�qj"�&�� �6��9U���q��X�@�̇9����%�)Fq�U�%rW�Ѓ�SG�&��~��p"EB�O�w{�c��\҈�9�;�Λ�Kt��P���3���7�yd��r'g�w�4O@���:��KĻ��$nw����E��|{goRK�����g29i����$��PK
    +Q�HO�8��  �  9  org/bridj/cpp/com/OLEAutomationLibrary$CUSTDATAITEM.class  �      �      �R]kQ=��mҍ��VS�m��$���CDX�V��4�w7�xC�[6����(� >�����5�(>ܙ��q�Ι��Ǘ� ��)�������p��ן�̌B"B�{�r�;l]v{�fϴzgo4a�Wa7"7�8#����*�g#1��k��@��]	���S�+B�V��(�TB�\�VM	/������H;��
�ח�)�l�B��s%���gb�,�	BF��M{���Ա��"2�&T���r�P�m~�LΩLZ��jK��x�J�7]��vp��*�����L�f"��vWN�7/,��k��ҫ�����l���ؾ+�}(�e/�[y�M��T/"/T�WS����0Y��������*N�-ϓAk,�S9�����F�)�O��1ߎY�|�3�ldp�R�;Q��O��8�G�8���|�N@����;��'�~����r
�{����l��S�p��~��e�\�z�wTc�!ԓ�<��ߠa�kPK
    +Q�H�1
  �  1  org/bridj/cpp/com/OLEAutomationLibrary$DATE.class  �      
      �PMK�@������j�� �6�GE(��졥�M��$[6���I���G�/Q��Aw�ٙ�vxþ��8�6�D��06j���r&:'�xXY��t���=��=a��0��J�$Neb=���Y�x�����!��4B�R�^Z�G� ]�>\�r�>��p�#��Fz!	�H'"��D��Y�^�
yW�4��+��U��(�e�,e�=8�^ěs1�X�7h� xf�`�1�*b�|o��S�K�~󲍭�C�=���	PK
    +Q�H��'  �  7  org/bridj/cpp/com/OLEAutomationLibrary$DISPPARAMS.class  �            �OMK�@}Ӧ�M��*�GAD=J��P�B!�b���v�m�l6�?˓�����U�Ń�2oߛ��ُϷw �:�>D�Փ,��y$�,�W�ҙ�p��N�����d4���nD�]�%Ζ��LI�J����L<	��������LB�\��]�G��<4	�{����#g��7Eh�F��XX-ҩ�_ ��\ݖ�TٟH���Ju�"乲��(
U`^gać�cl��.5P;yE�¤�M��;�ul��pԄG!������e���XC�PK
    +Q�H���  �  6  org/bridj/cpp/com/OLEAutomationLibrary$EXCEPINFO.class  �            �OMK�@}Ӧ���j��GAD=?�� ��Bh�J�Iݐf�f#��<	��(qE/t�y���>f�����	6	����Q�4H�� ѳ 
�W��3a��Caw�����p4�\���[S&6�S�Xu��o��T<��ߦ�hZ�#	��+{I��L|��yp�Lp�*���q�ޞ�JB'ԉ�&�(g�f�v�r9*g�4_o�K�ȁZ����2Q��j��"�/��fuVi�q���Ik��g+X�{�������u��lTb�b	�PK
    +Q�Hj�k�  �  =  org/bridj/cpp/com/OLEAutomationLibrary$ICreateErrorInfo.class  �            �O�J�0}��m�Z�uģ �,�DA�
��.({O�QS�fIS���$x��(1�^b���{ɼ�����8��X�0�r��|��*�I2���*���Ld��~܉#-�c����[��ߋ��t�f���o>�{`�ݿu���?[�3YJsN��������b��5��"�$��թ���\F��,�1-Y����D��.R���Z՚�Kِ .K���U�����,�ag�8�,l9�;xF�d��O+X�y�n�U����zX���q�a	�PK
    +Q�H�dP  �  ;  org/bridj/cpp/com/OLEAutomationLibrary$ICreateTypeLib.class  �            �O�J�@}������*�GAD=<�E��P�`�}�.�!ɖM"��<	� ?J�D/��f�۝7��o� ΰC8��я���~�X����(���+��J�"T�fy0���.�%D�]-&�(NeR9��~s9Mų ����0XmL��T��kB��x��E�n��J�E��]�A��0
u"��0Ję�6@����uK��6��S��E!M����%�a�H�"��q��o9�;y�����޷�8o�[%��Q���m΍�k�PK
    +Q�H�z�H  �  <  org/bridj/cpp/com/OLEAutomationLibrary$ICreateTypeLib2.class  �            �OMK�0���[��� �`Y"(����.�,xL�ASڦ���?˓����_�Ń��y�I2o����
`�M6�^h�<��<�"�z���*u*J��@�F����7R�r��%K�6�����?���XF��6a�7��X<
��ߚڰ��	ֹ�TyAh��\��8�`��)TA8���3v��\��D2F�0��8H�2yS��4_�s�+�kUw�e���(
Y`-�T���̼���g�O�ia�����U�뼬F���As����M6��� PK
    +Q�H�Dy
  �  7  org/bridj/cpp/com/OLEAutomationLibrary$IErrorInfo.class  �      
      �OMK�@}�����jģ ��GE�P!lA�}���!ɖM"��<	��(q<�,�fߛ��}{y0�6a�͝�H�d�����hrQW:��E�b#��~81F�������,�ͦq*��A���[��T<����9�	��P�}�
U�:�Gs}�.�X%t�{U�ѿr�Ł^H�0҉���(g�� R����X�/ŽֵI�j��4A&�R�؃��4F|x;�3��@���_,l0z�"ְ�q��n�����U[�6���PK
    +Q�Hkv'5  �  :  org/bridj/cpp/com/OLEAutomationLibrary$INTERFACEDATA.class  �      5      �UOS�@}���"R����"���XDji%Z��N9:i��0mRӔn~?�qp��͋��ի^�#8�6�/����f���}o�|�}��$��5}3�֕�v(S(�2Z>���EJ���ESJZ���q%[�G���H2� c�UV�z)c��������cb[ڑFO��@;Cg-��)�.ǒK��e�.w噡}NQc�A�Rx��g�ƖRd�I�bI��U���VV2h�}�@�SMQY����QIUCqE�ei�mGʕd�R�M�z����a��6�3x�`�ڔ��Dg��7`��
��Tz0��n����@�u륅��֌�򺂫\��Rc��i�UDx���4��(�g#�s�IfT�b�M1��e9����y�D1�<����	H� ��|˓�~�e�;�ՔC�S���i��3Ld�n�l��o���$aۣZV�#��2R.%銔��I~���*���rkĵ�l��Qҩ��ً�j��k%�P�rJ)*�QU�0��|_���¡�MRmM@�Ѽ�/��L��V�3r\�&yDU��hN*�"�)u;�V���J���4E-��-�]��c�<�=�A�E7�����;؅���	0M-�u��BP���Wu(�*�v>"|��Y�Cj;h���>>z؂N�b�)C���Z��&��<g���i}􈘏�R�"���g�|���~h���Q�	�A���'v;���_�.|��c43�O��}��;ѿo��'L�)r��7��>�+�4�6��5b��K?)�1�{ֱY8r���6���ݩ��I^��^�\ӆG�zM<U���AĮ?PK
    +Q�H�@��  �  5  org/bridj/cpp/com/OLEAutomationLibrary$ITypeLib.class  �            �O�J�@}��I��*�GAD=zV	
�,�o�E7$ٰI�~�'���G������o���73����
`�=��ͽ�J��(�Xg�,�\ו�D�t���>�.օd��?M�|>�W:�����x��us`��-	���UuE蜜.=��b�ЭTI����[���Q�c�.�Q"J��0T����H�/Žӵ��j�7�si�T��,q��iq�l�Cf~ˁ��3�'>X�f�>Elb��o�U&|?j_��˹)c�A�PK
    +Q�HT�r2  6  7  org/bridj/cpp/com/OLEAutomationLibrary$METHODDATA.class  6      2      �W[wU�'I�4M-Z)ELSl�/-HmII[ljZo�i2�S�I��A����(��W_����k����O.�33I��Ʌ�x�\�9�����}g&��ǟ �{��%YR��J$��I��X���&䄴�ʥ�ScsgfN���E�`���%5���f�VĴ慛��	`hEX4G�E;����P�:�Eg�S�����-C�I�X4���L��0�Jw�,i'ܡ�T ���A��,�G�m���������� 8W�dMThAOŨ ˑqI�eh�mM�E7�.���=aMJ|f$��������x��;+j&���0�a	�;�`/����3�	9,hɛnժ+R[�+��I�b�W�&xUFr���ĖEH��N�6�\��d-�/0���N��)OS�WW3�&�QM8I��B���\�,��Aw��2��*e�����R,Q��#\�����@0��U�&x�sc��xh���v�Ռ�k3N�\�����`�FlF2<��D��|��C��e=�8���N
0.kM�`g9W��o-�N���Npq��q(�8m\��Rl��	L��h'r��;����2cr1�����h��I���&�P��׹�7Ά��Z�&�V�;�T_W��coB�ږ�5�J�=^�^gB�t���PNT���E�9�ƶtTɪ<Cm�c��h�#�y��8���^�I���h��rAi�v�(P�1��d�Y�X�z�<���D՛��4b(�o��*`�G�>�S״YQ+*2��K�P�7�X7~DO�
z3nM�B.%(�������	I���%Q1G:�RV��:�Lk��}�EY��bJR%�rAӽQ�z�d��ZR���עh-	��w���7�G�-@���͇A�`����3����۴֚÷���ş,��8.�^�eYTb9AUE�h���c�ѷ1}����;Jg������z���� �a;��ӏ�?p�����A/�:�1:���o�vo��_,(�
�v>����k>��tG�#�k�C:E�]ƀ�@(���:x�1g�����/��|d�������v��_�Ƀ�A���t��0��Z�}eb���g#�?on�I|�f"5��4�;h"}e��쟧���C\�N��$��N�g�����J��%����7if�M�j��60z�����nZ��M���'L��T��wm{6o&���0^�<LNw�	"F�F��"��1���k��t�J1B�����8zѾ��;���1�CN�}��������a�*���Ì�"�9�\��T)�>?���V�9��,��~�n�|�~:oV�7V���Ћ��䥺N����~Z@�J~��Y6ɿ����N�$��'+��F�'�d��ͬԨ!_S5t�*�mҹ�|khŒ�ur骝"��s��k�
���N#����M:u�[���V:m&ܰ*��c���c�	]&&�ls��,��}�J�-t�o�9�����\���V�ȅid��ަ\�ɪ�Y�oC�-2&��9���م��`��G.�JW��g���w�.xiu��q	��S}�PK
    +Q�H��m�c  �	  5  org/bridj/cpp/com/OLEAutomationLibrary$NUMPARSE.class  �	      c      ���S�P��M��U�
��O�R|��(�p2S�E7�i,aJI
�έnt�V7:�Bg�q����ݤs�>t����{�s������'�1�a�[v9_���Z^���k�z~�0?Su�u�5,�`m�~ѷ�����	0�νMˮ]�ܥ⚮�	D�¶���[*Ck��3$�vd�O��N3D�+i�A�E�!��X�1I[�9��9*�T��/z�D�ؖZ��bɰ�ģ+K�iEG$t2�'p�!U�]�t=g��l��G8�(i�@��.�0\�*�q����[o�n
z
�y�3�`$9�g}�&A�zq�qR���3���s����n�ߑF֗2ȥ�����U|�/eHh��CG/q%ݡTm���}�e�4o����j<w�2J�{_<ዯӭ1�m�c�\�[��/��E7鄳VI��V�4���چZ������`��bu��۵J��������T�1M��>]By٪ښ�`paZ1Mݞ����;8C�����#������Ez3/��/n�3�q �=K?�!D����͹�%D<����c��7��.�>�8�H=��q�����e�/\������[v����]�N�f�G�8G��B��,�[dЇ�c�"!�I���£��>�k��".Q%[�A�%�ŀ�e8�hSY!�41�l�A.��Pc��1���p��,�G<�p���������`����3���T�� ����g� ޔ��r�l[d(k(�+���[�`�*u$Zb�Rxճg�h�`B������Z8���D�7��-U��0H������g� ٔ���=1�l��t8�[�����'�{{bX�V��n�PK
    +Q�H����  �  6  org/bridj/cpp/com/OLEAutomationLibrary$PARAMDATA.class  �            �TKOQ���1+OE@EۂO_E�0M*���fZ&eH;�3�&��X@bjb�;]�[��ѿa<w:} ���s��{��O�޾0�e�I��KYS�ޕr{{R�(Jk��D�6���zZ˚��?���H<[Jl&�`}'Q�m�r�ZvW��~x���O�*e�a�����1�)|���H4B�/����f1L����8�Z�V�������_74�VM��{ʫ躴���m򷕕BI���`4��']/Hj-Bz�����x��e�p^�]B�a"ҀU7�j�eW0 ��O#M.D[�&lէ%��V3Rj�5\�y3�o̧�@HE�K��Tr<l�����B���ň��!r^�'�qU�ܦ>�mg|d�7�R^�1L�-p�/��!���f�a."��i�UK8t6�����4g�a`2kٮ�%z�'�I^�}r$�m⮴�S
�ԔlA���1���j��UM������%���������o�t[+���+���TK`_-��ޟ�7��Y-ɚi���rE�(�9uE�e�R���ɂbY��aR��?�ߐ��h}Ho3dٶ���h# Nk��D.������!����q`�,�+�^�R�S��a�x
��=�;<r�,�1�v�u�ӕB�}Յ�P���B�Up#��=x_���0F(~�{n��$���.y����0JG�|�,'Ĉ7�5VO8&4�?�'|q���I1��V?o����}�O}́�t!�jt�T0;iJ�nQ��$��T��Hщ�����:��`k���:��?H���K:1m�.�qh4�PK
    +Q�H5��	�  K  4  org/bridj/cpp/com/OLEAutomationLibrary$REGKIND.class  K      �      �TmSW~n�%ɲ&����v[V[-H��HBJ,i�:����lv��ƙ����:�P��ӏ�(�soV	f��{ν�9�yν���� ��ä�յ�gmmk������ʥ�B�w�o�Nɪz����Z��Jau)
��Oi�xdh��Ե��j̖�����:Qp��a�̭cB1$�Ӊ"�0vD�(ҽ '9
Õ/#E�!�`H�?�r����:õ~+a�B������O���j�Az�a`EJ>QY(m�t�����HM�j���
R8G�Q�$V5�u�Ո����Y�iogd��Y�,��0,�];u߳��L��*nv�,�F�9�w�� J��	_3D�A�S���F��c�st�z�-3��^+���	\��Q0�a.U�r�Y�xX�P�b�oz��z$���-[+q"pj/���6�I*4���MJe���0\R�ލ���S�.�n0�ط�M�ar��~ํJ皥�bwS�^����Le��yۨ�;Y�x���G���O2�0O����@v���ż�s�(8�żCBA��cHJ�|!�N�Lz/�[TE�d9�j�Q5�u�j�n�5î��� ׭�c�-��Utw�gc���Z9J�c�ɺ��jf��ĕ�㘞��fs~�j�@o�|���M6�-������wL>��x?�ԯ�]$�?�����O�cX�q@�=���p>�?MyTN�����!�?�F��B���v#�xWi���wP�^	5{�9�;�1F�r���;�q�a�� <#�����S�c������}���I���4�s�M�'J�Ҧ_����"�hTH���1@�NTy!�����A�X�)]8�8����X�٦U��� ��Z
�_"���+Dd��$�������6���H+����=�)�v>�6��OH���M�=&�a�.l��bFs���PK
    +Q�H��%�  9  4  org/bridj/cpp/com/OLEAutomationLibrary$SYSKIND.class  9      �      �T�SW�n�%ɲ�Ƣ֊��-k �J�JB�jlꃳ	k��f��l�}�C:��LE��c���Q���� aư��s|�;�9w���? Y��0�z5��Y�Z����ֵ���B�w�o�NѪx��h\/����(��⦱eh��Դ%�Y�-�237�q#��%�n���bH�E�a� Q�1��ANp��F �8C4`��ٽ;����K��о>5��w}!� mq��@�㥅��%�!{�w�>��`�R�=_W���8B��(��ڮC���tG�W6ͪOgS8!�8>#�"��}�E���{�S�I����N��m43�pwwQ:��2$|�q�:QO�F�Z���Q�ta�/�K#�v�%�8�#\P0�!.U�b��X�xXMS�b�oz��z$���-[��D�X{5��6�I*4�Ш?�6}�a8�Q7y���q	SGvmEqY�W���\%���[/��,�:��~37�c2�E,��'�m�& �eȨ��{�?���1�y�e�j��P�.�9kI��#\�bH(H��BZ_H�@ku��ι��@�r̵f�bz���-��V�dx��Ÿn��oz4����+]s�?��AR
M�ݦW5�-N\�;���7�Y�]�5H�)�@6�n1ě<��1������[7���,��m����;��<�i�{[t�$N�)"_����μC��A�Qi��Y��!^U9�
��T2�^B͜���1F�r���;�q�a�� �F������u�b�ˀ��2ϑy�������I#=���4y"Jm��f؟�^��%���	�&�*O$vj�;X؋k��� ��}�\��&��o�B��b8��ϰ"�|Dު���0��F�[ZocE/G�����m�Пa����&��!I�c����"�-a�$le�1������PK
    +Q�H�X�  N  7  org/bridj/cpp/com/OLEAutomationLibrary$SYSTEMTIME.class  N            ���s�DƟ�?��vS�6�
�8��$��P��P&����RGJ%9�8����p��vҙ2��p�\����w�&+����>����V�����4^a�vܫ��k5����B��(�*�Ŷ�l������	���R����E�ato���_���_A�a,��̺�e0����$��ד!�`ٖ�!��\�`��8�q��f+�y#���+���:ñ}�mJ��jrՖ�j�1B�!�a8Z��_��gpǆ1�Q�#�y�1d�����~��p<r$�˓z�c\��3����k�Y�`��;��x��<���p �	�:���i'U��i:��c�k=�qm9!z������/��5.b8�W�)!~�Z�).��(��`F����]���p| $sB���]���W�!�
ق�=�e��p�&�%�L�lQȖ	-o�,/���Xa�Œ�XR�M,9M����0Z��k����/#�6/�7�۩��ڶ}k�\�<�
�����iz���5̒Ņ��m��R��<��)��O$��]_��,�3���dns��5#����W��Â5�c��Fp����I������c;8qSrQ��$y�]�%�OӽF�#e�X��X.S�!�\X�����]�Q1�1�w#x���܄ʮ�[h��#�m_ !�I������7%�Ԯ}*dߦ�ߢJ���@ސN���}䤐o���-4�<ޛ�l�61x�*S]$b��L`� ї���=b�~���B4���d����T��� 9��䀳�e4�d_3Rȏ��'�e�dp�7��Sb�U�0Pb���2��җ���1�n���h���_��,ta���Wr�g�h������o�-4��fp�7��;b�=Uw��0H�G�������B(v d;����1���`̟���pK���)����_�R�F!�uS�MN�B�مB����BI��;Q�#�C��h
/�� ��I���Z�&�����B�� PK
    +Q�H�.��  H  2  org/bridj/cpp/com/OLEAutomationLibrary$UDATE.class  H      �      ��_OA����_[�**�X*�"�&c%iRh�VOf[F�����-��ă&��~}���l-���dwf���;w�L�����"lg/[q�n-[=8�V�F�T�皞�0=i[EYqL�h��z�����N��9ͪW��DՋ @��Sm�f�����"B�aq�����,6��A�|�O�%���@j~;�8:�"�}�2���`���a%5?h]�.�2-+�!E}��C��>���	c�^���8.�J&���Lr�𶸃C�:_������W�[�d�i\�1��l��u��zG��率����`9c�vNu���c�1��
8Ǉ�2�����{^l��b�:�y���]���^͊7|��i)�=�ρ5{W��E�jַMG���(�a�(-��lT�ӎL<oZ�l�m�J�,����]u�SR%��%�����e9�o������B��-�H*�����<�8N������Q͂�!H�ym��[!��&�p58��/����]����������/ ��n���m��S�'�s܃���?{��|d��\��k����<�B��g��ֆ���q���5��Aٶ��8Qa�i�/��<��G���>|aM���5!���E8;�Y��PK
    +Q�H�M3d  �  ,  org/bridj/cpp/com/OLEAutomationLibrary.class  �      d      ��y`U���춤i�&�N1-�!������&�v�fwӖ+l�i�4�-�Mi �8T<�EEETO<��[�E~^��}s���of2����3�7�}��f�3;�}��b�u��U؉��h�Jq���:��㝙T26Y-���r)U�S)T�������
�c��hgf�E�p����ƭ�F�Ua�R��B��i=Ca��&u�-(�����靵�R�8�C�)�����s0̃�t.�����D,kb��*5)�+���dn[&a�Y���+씀2bZ���Da��PB:����&��h��6�u0x����vw6��ϩ�0|-��pp���l�t�h��&�m�q�
���q
k�-���O���L{>�A`�h$�쀑�l;���N
*�H�:��33�1�8-ٷCM'���5YPCb�T<�lb�<�y7���m� x��d�R�����&v*��a��TF���:���mU�i���MС�������4*�Ժ�5�-
[,�ϕ*��"Y���+��ײC9-���t���m*�A��S|HaKc�_���T>�I�v�p6o�j,��g�C�T�7_	'�A���}Zr�_M�?��S $ϩ��L��d<7�3��-��]�t2���xh5s�0���Z�m3�e��X:����})�Y��h�I�q;�i�a^*3�'��X���å-3 f[
`�%Ӱ�W�`�/��`���c+l%�H��~�e��07�Y�!'	ށTވ�<�0��%�r���Xv�H��C��B��"��C8��]av�	W9�J$�j,��n�饦�� a\aB��3�~��s�l�A�^6�e�}
[Ng���aZэ�bFʊ<��e�]SIg*��D?�g�<+��qp��%��*�,��.����P����$\��2~
���ۆxn�Zn�@R�v��"YN��%we�9�=;qֺX�&[K�򥙀4��򩜚��~�g�)��EV~L�>�W>;]��,�t,5�-f
4�DV��4/���5Պ&�#2��.����ә��d_Rì�S%m"<fQ[)�73����/	*V����c|�d�=ٜ��>�ǲ;�r�!-�M����,��
;bs�T���1ܱn����ݸ��Mp1��+N(�#�	��řB�dqldP�L�C$x�8;5+g��biDb��b��W�X��)���LU���Wv���������y�o��]�m]�j+\�ۡ��K~��q��C���(A�"���⡮E�5��d�*�@��P���Iۦ]�۲��z�R)L���YWi钇'��m�p�S�(luGv�G�V���x�\��U�����∑��>1\)0���:d���N�y\�Z��@N�R�������>���
�px�,[(ϝ-�U�����q��1�e)��)O�F<&� @BʒІ�q8�Q'������B�
En��fTW ���Z��UK#�!i��L�=�Oˋ��N�q��h~:�Y�G�?+E�*M.WF̵�{���*��IQ2Z�s��R�K��o8��a���' ���j�n>���넱T����r�yƱ6�+X#����lڱ���\-�rU����I�R_,��*\���cQ|L/T��V&�|�-��J�F�7�WS6k,�i�����l
�F��.�?Y��z�]Q��=@Ǩ��1����;�Y<��o�={%��)��dG��A=#[��yD�#��g�jqM��<$q�O�|���w{y�t'�a9�ŉ�x�۴�˜�&rOE1i�1���$3G��E��d��2Fd�b4��H��p�!3�"�w{�#�b�E$�"Ļ�."y�����Ed�"�wɻ��]�x���J�E�LF%wQ�;G�a�s9�����Feg���QᏃ*���wd�pV�S�I��("Q��FR��TjR*59���JMN�&�R�R�ɩ�H*59���JMJ�EQL�u�Ѣ�;�;Mʝ&�N�s�ɹӢ�wQɻ���?�p�����>�
��ʬ��<�X���B@���6DhC�?s��a��)y��7��5>%��D;�E$�bҤc�6�Y�&�Mt�n	�-�1"c�ȫ�"�v�g������B֊:s�k�v%P��=Xߨ̚1�7�X�5	Ͼm���dm�H ��L>u�@wӆ(m0�v�m��|"o�(*<`mb�gn�3Қ��5/8B8*�F�k�����V)V��Em��@��׼�*<���r�|Y7��DQL�tL\�Q�(q.Ҥ�E%*ƈ��^Qt8#RlxgV�N��Ⱝ)�T��j�Q�,��Ud�~���E])�!,��K�<��~�kD�rՓ-;�Gd�#������;*LP�5"���&��_#���5J|�ʾEeߢ�oQٷ��[��5J���Fe_���(ɳ\�Qe���k8�kK�®K�[l�ncDƨ��|TT&&:�[�w��m�]Ķn�²9�F���.�g|� �n~Go������@��1�u'n�j��3��uuh6u��L8�##bt��s߼�w�@�Ńb��xH����'��~Z:,��#��=���)�@k����o��m�3|�I�ac0�Z��	G�
s׈��kb���'�����8���P#�f�P/�^�c���5Bn씬�x�j���;ɋa��_�F�&�G�����a���a'S1�y�w��]e됑r�cDΐW��;e+����i\k��u�jǐ�D�P�ť��BeBOO������O��qs�M��p���d��e��Z���\y�|��������j�1WF"�S{�����U����DU7Ŭr���>���F�S�R����~8��D�����N]�?R�J�Iky)>���r������v�UE�u
�-W���q}����:�|mJ�OV*zi���HD !Nf�D̼=z���2�W���z��&�\y�^���g�jOCX�R�o�y��k^��WI�,�¸תt��^��䩉��^+�y�Z�x(쒀�o������#7���d�٘����Bux��2��7S�ㅱ����k�>
�+�#�����q��sj[ab�3��?�'Z�˘ZK�������u����v-���m.��*F4}T����P���E|�܊�����I�25P�����J���D˒|iZ[��)�An�J"�t~��QVO/����''��ǥ6�Y���9�z���M�p�b	j	���R�4R.MT�Z2h��</^��Ty�0f\f���9�HMK�y��Z����R�:Y���]�ޜrޓ���0����pW�
��/���c��U�A}`�n/Ǹt䯠���́Foq�➁����9�d�
��]Sn��`��k�+����S�ޠ�����#�����&7�M�4-��'�O'�V��i{���9�#���L0X�(�
7j���P*����p1�1��`u���NM�N�I��H>n��q3�p�}r���{az}�s�6�5g�g��+�3�w X���9����L����k7�kJ^>g������Qq�u�9S�:oGY��x.#+�7�3g���U;��`W�Nw���K1S��^͗��ʗ���F��ڏD�6�T���ѳ鮀Xs��Y��j릀�Z��[�u�@�pͣ�ѢϹ�MF�ru�z�W&׹�#�Q��s{Mҳ�˫��}]��z�����HO\^���뺦\��j�U.v�[\?���+�����[%"�AKP�~�U�J_�(\�����rg�)+w�����`#'�l���;�Dw�7p�b�g�5q�����X�y���X�F���}7��=�3p��3p��3p���Ι��ɚ��gO-��[���s�[����������qo�S���)L��s:����ͥ�>'sԷ����BAr-x�F�Ht}�Jϵj83#�EE�X���+w���rg�y�;7�����	���:˭�N�]'`�sP'`�'�M�DyrϘ.z��G��gB��>gQ���FNIb�O��ރ����u�JI�9����C�R���W��'��S��S��S�S tqK���7Hйu��A�� /h�T����AUw]z��bD�5�F\LhD�U�F\b��T��r�t����Vr�����

s7�����_��峞��ߟ�M����j����D�~�c�-��[�����כd����"7�g��꘭F����r��Ν,_Uh��m𻱠�}�,hw�[���ނv��9���j佈,:V�]�,#�󌠷���W��d��Ոc�9,`IB��K谀�	�B��]8e��bhj�{]��YU����}�Q�Ȋ6�~���w��W=�}��BN��9�R�,�u�񭿑گ��X��E�������]L��]����W�SkEt���>J��k�0譗z���K?�w*ݾ���i�L�W7P��j�[���Y�_��7���	n�º��ׯ�z^|�������cM�o�[�*�	�$���\;�y�a\���}�}f[dLu����t�F������Xv�������Z��^�Y�t�̬�}����N��s���MSk���'5w�������;he;�^:�x�kq��2��z3�>��I��n_R�/'sSO��K/5&���L@��jXi3��4��ڿҨ	P��k$��'����a�����2XX����-��' j�������&.�������1S�S�en����ھ���Gfe�55\��ؔ;g�K맮����J�G�w�.6���˴��a�l6�բ��t���ؿ�e�_�+OV���"��-j��W�c��	��{�� � �<b�cQ��%X�)��;[���6`�v��S���qx ����,pqx�N�]D�nb�9��s����|�!��� A��E<
���+{/B�x�8p��/� ��B�O���'��x]B�"�Ny�������b��_
|%��UĞ��������+���"��&��!|-�w�W���{-��zį~=��"���oP.f
��(h9Z6��������7�û�4���ldoa7CS��Oc[ؼ�Ǖfv{+c�}��qy��������!x'�;ٻ�~7�C�n�;�{��^v��s��G���������D�/ ����!�{��{&_*�v���Ư�5���u�8�`�}�~����@� ?@���S�u�	?D���g�g�~���H�����(��~������e��"�GI���*��k�ǀ��x��K��D\~�� �6⋁�þ+��8�����#;'���U��~$x�	4�����'h�!������)�_�_
��W�I��?�~-&���Dl�i�8lw����w�_�{��W ���I�K��L����U��#�����U�� ��f��2�g��	~9�P8^�o4m_	���U��E�_=���!�W?�ܿ�0r�Z�Nv���+ȽW�d�J�����|Y�rr���M��� �_܌�=�B������7� }7 �"���{#p��&�v"o	ѷ�_��}3�r���-�+��7�B�����V�5H�ۀ�"����۴�+G!�o>��v�c��� >��N�㈺�s�'ǟ���.�P8n~r���'��/D����N�uH�{��#��>	����؀̹�d��oD�x?p'
Q�E�w#w> ��苠��|*r������|�t�����H�=�/B�?�b�����?�s/�f4;>
|&r�c�[�������x�ő�C�ő��'���'��� �E�? ܇�x��)`���t��#sށ�8�fç�����N��~ ��Y೉>���"��!�?�G�x���N$������Lw72��s��_>��e���lx�|�� _@��.$�(<_�C�F�x��u`]�+����>��.*	�3�o�g�o�`?t��<<���pI)�6�~�`�w�+D�1�J�O}�K��2%�q�KQ��|��_N��/!W�+f,�����r1�\E����b�����
b�+�9�"���D�5��-��_G.���k/�5r�v�RP�^.Ŕ�ɥ��z�T� �����M�����RP����\�)o�K?�f��Sn!�~+	��f���$�����N��v��w�쿓�1��$�w�w�쿇d��$�w!�? ~��C��#{~��'���nd��D��1��P8~�a���C�}��s/9�Q��c�����s����� ���^� ��3W��$�اHe� �"��Ie����ļ���ϑJ���9�ER	>B*�/!}��2��+�GQ8�����p<	�U�������k௣p��(��&Q�1�[������������?�������~�@��h�#���'�	��(��	zJ�����?S�������%��+�O��O��F~��7��o�����{�� ���G��?)6�!��J�od�ߕ�i��c+�i�`x��D�3����Q�o��3��!�_��#�,��2�a�p�p��<��	A�I~<Z@���B��	����ł�܆����Ȟ� /	-�_�e����"�R���B�^�,�0�;�ֱ/� ���,�p���1��:N�|���%^�xg��� ~~��M�/�(x���f�r|����/�:Y�"���N�-��8�
�w���^l,�s����nB�i��N�|Z�t�K���	^
�b�g�6^|fh����g��
^C�Z	܃���������	�N�z��#Ƿ���$3|$[�.>,8�
ʼ�C�Y��>��0�a��Q|�>���e���5�6ض�v)l��vlW�v5l���H��c`{,l�����ؾ �/�ml���$؞ۍ[װS`��M����4؞�_��v3lτ�Y��
���Ys��o9�o�`�����PK
    +Q�H=e��  �  "  org/bridj/cpp/com/OLELibrary.class  �      �      }SmSQ=��ZE�0�|K����%�(�aPu�~Y��ڲ�,���*?���Џjz��*�3���s?����9�ih5Ǩ�iz���vS;�|�5�;
��?�ɭ�vX;�� ̐�u����J�[�T�������)67nwu,�h
ꜭ��)U��b�hX�����OU܁�Dc���f����,0^�Ox�۾h�3dr�����mX�p�sj@aՕ�t���ÿ9a��&��y�zd�B2�˟2L�J+�2(�V�pFM�U��\�x�K!cf��D�dT˕�����S��>q-�Hpߧ�0��Es岔���RE� [~��ޭ��n�( -5?a�5FƋ��o����ֲ��TwD�h��y��ؤ��:����:7O�c�)N�B(��f���L��hX��8���zߗ��͝m��ܡˤ�e�.wۢז�o�e��\��4e�)9��F�F�L�G{�)�D^G ?q0�ߠ�%��(2���O�_�&�W��~)LP|Mߘ��a	L"M]o�޷xGQ�S �q��[�LQ�P^i��:��gx�:��/%x���|KRF���8��B�ؗy��؇��@�{&��s�r�XR�a	')��w���5mƃTZ�{�5B�	Po�9ȷ=҄��z�I,�"[�B���U\]�"�O���^G�%���v<��;M��ou��I�PK
    +Q�H"(��  E    org/bridj/cpp/com/RECT.class  E      �      �S]OA�C?Yk�OEm�P���H��D �ɘ�v-C�]\�<�o"��`�?�e<3ۀl��C���9sν�N�������i�Ѱ���U������A�������N�ع�m�l�Y�wl���^��۷�,F#�3�����+x�)0�Y���h�?D��8��].^1�d��z�0(J}��b�2-���h��$����PŲ����u�4j�z'F=�;_X���f��A�f4�y��QF�uG(��h"���U�ȖL�I�����L)۽�����iKҲ)�-y�1����|�q>��@7E�4rN	�@v��&�)Q&e�㇘���{Bz0\�	 ��1�U����`� ���A���0���g[���s��pv��(U��լ:~;3�~~ȑx㺞��\���Z���C� �ʱQ?&�w�u�<"C��~��]O/��A�k�K��U�)�]jQ�"*k�~�H.rB��!��a�^bM�F@.�A7�6�*��Gf@;uBwr�N��%}@,�Rt����<{����I��k��)��A����qH"y*��XE7k�d�x��ouEf�ދ�^dB��G��ˤ)�����^�%*�f��.^Į��]�s�V�E�R/fC�ڈ5�L��{��C7��.^į䅧+��{�ԋ�P�-�#�L5k�x~�a�/��+�
�NL��!{Lؔ�PK
    +Q�Hj[��    !  org/bridj/cpp/com/SAFEARRAY.class              ��_SUƟCBh-�J�V�����Sk 	���5��"*n6[�4��͆���Jo�ߡuƉ3���C9���6!��?̰gs�=��<�sv����+ �Qe�5��l�ҫGY��8�����/n����^�a�S �VS�w*G�jGb8�.]>RN��R�Z1�l�i�z]�1DN�ZSc�p�b��xtE7t{�!�^�M`�8�g�O��\��O.��zC,��<6��V��B�#��mÉ%��8�c�ä�y3��-?1-[h2\N��@9iAN�ތ�"f���!&��s��eN�-��ů00
=&\�~$jԌ�'1�8����EM�����h['�|E�Ni�!�V�jZ]3l���W�0�Sr�&��@rk�yniP���Y�>�%��ns�(�DG���uta`	7y~�Ԓ�>�C<���^u�֩�����t���g��3u��,qt�IB�N�f��`�I`E��s�适A����loA��.��J�n�+V2k��|�Rb�@r8���dހ�1��Z��b6���%�[�r����cy��sӬ�gc�vM��*��Tj�}~!%�ж���f�3��/ʮ��i"o��غi�Q��CCy��A��D���tz�����|ɠ-[b]��;���u��y�]��q�lZ�V�k�󰀙��}R�G��42N7����5�Lb�hܧ�Q1s��I�AU{�WH��3c:j��s�Bܧp��u���I!9�J��_�Hζp5�-:�<sE�]���}ъ?���u���57�:��X���8��#k��|�[��H3�=��bP�L�`��=&�4��),3X���+��R���>di��`^��B�f ����/�%|�eR��E��ߧAV�3��?�5�Y��`t(�����f0:�����O4��[��%	d����+�3���f6�I���-|�b �_���k� �%Wz��Et����Pء���|f���o4��6���<�{��݈r���.z���m�5���?s+��~~�����*UD��{�#��%hn�G4���H;)_U�PK
    +Q�HR�ė  �  &  org/bridj/cpp/com/SAFEARRAYBOUND.class  �      �      �SmO�P~�mN�E@^٪R����ti ����K���_�&f&~�������6>���s�}��<=����/ +x�0�5��jî���jzu�R(n���Ƿ;�7�`cݪ��h��N��2�8$����Ƒ�0�w����[�o׭<C��pZ�ȩ����5۵}b&es�)@�E�!�����e�	d��r����M��1���)ږS�Kd"�w�OG���Oa#�`�a��<�q���k�/��}8��ZNKa�d��$�bV�]EK�y~�����6f8�,#��ЇO��0+Hd0-��E���W��[6��m��=w_�DS�&�"q����>��K-]Ij�y��bK\�C���H,qOZ�I-qKP�����j4vC�gήѰ��c��CF�]k�U�Z� 3L�ݴ)Qp]�7|�si���j�V�v,�x�O�G��J�*��Ř��o���%��Ni\�����<�5�T�*�$����S�6��{�>�U�њ�� =qCr:��$�~�9�Ɯ�5��|��<�ϋV���������@�:�҄B�w�&�{�!|�~�T)���D�X>��]�PU�b@R�j�CR�Ct�����$>M�h�b��6�x�g��h�P�Ë�����m�Gj>�M��&PK
    +Q�H����w	      org/bridj/cpp/com/VARENUM.class        w	      ��}p�Eǿ{y��e�l�'�M���&9��o$�\����K.�]�E!IC�zI�5�����耎��#2"c��^�7�Tt@GtG`DGt@Q����Ӧ�-��}����߾�s�w���أ ���u˹���\f߁��������@*M�Lz��f���K����š���\SYZI�fW��/�ғ�"�����(d�w�ӑ�����&��i����ॆS3�(C�"���q��5GӺ�X0ҥ�D2�P�Hb:�7��㱸i�Qz�h�Hp*�����S�=S:�F&��,�
�'
�n�L(���q�z�qK�XdLg��3Ѥn9�LXP!���x��T�͔K�$�P|,�L���r��j�E�����Ñh(�t�"�m�A(8�O$c��.jRq�"4vIld"4J3���UjRj��z"�ф�*g�U:{�h3w�8����zz��P<2��FC��=�'��`b�S�N��CNLv.6A�H�3�C�޳>I���!�f��Z
b�����5�]^��,�oVl����
���A��*�2��M��J.����s۲��hv�С�ӥ8�KG��1�C"�K��4ˊ�v��e�2+;�z��E&:Sէ��L	L"�0-��:�Bh�����<'�?Ϭ,�fW�sN3�ՕL61�&Pu.g��s��C^\H�!*���������͘Xpv�"��!:	KN���)�)�%��_�[^L���?�v�OM��<��Ѳ�1��h���W)����O�=u�Ϙm���ڗ����vڨG���S�XKE�9�y��X�X�8D��# ��0G�k�J����Ե���~��̵e�~�C��P@j��r�zʵ�,G�k�@���pT���Q��8,��,mo�r-��J�opT�VTk�-�ז�h��Zז
�j{G�k�@��sԻ�\�^�G9\[!Р��9][)Ш�8�\k	4i�S�f�V	4k�G�k�Z��G�kkZ��-�:��
����m��h���h����m������mX��[\�$�A�sltm��Fm���E��,���t�@��E]�
ti[ʱɵ#�����v�@���=��Ѷ��׵!�^m�8����q�kw	��m7G�k������7V�7�_ۭ��m%�Y�A�c��h;̱��k�n�6ı��w�ت��6c��n�6Ʊ]`���rtyBe��������B.9;�U����l65��8��E����ٕ�����p�|�s��~�m=ӡ�~}�����B8�]�� t��o��9�h��KQ���J�r�
�JC˰ʰڰưְΰް��ѰɰٰŰ�p�a�a�a��z������]���{{����n60�b��p��v��{t���\��0��K��Z�c?IQ}:��gc��G�E���{���S�0v���:�W��z������]�݈R��<��E���ȃ�ԋ�M�₮u�#q�x�jj�dJ��;%g�y*[)�]���K���l��u!��3f~3������甩�k�v)�ӥo�6@�Z-���h�wq�f�g���m�ü��OSu��C8pj�?�5y.7y.��!��S�Zz���']��W� ���*���T�����U|��?Rh�*�Z��Z�F�ת�:n�*�^ş����Jܠč�zܤ��J|NR��+q�_�E���mJ|Y�,|E�;���,��u%�T�RX�K�����,�p�G�8*K-�Jܯ���JS�)-|W�ǔx\�[xB��������C%�V�Yi��J<��Ϥe��J<��/d��_*����~�ċJ�$k,�N���xE�ZxU�ה�����'%^W�/���_�xS���W�m%�)-�K�w���l��_G08��1�l1�2���y��iS,[-&�)�F�u+W�ҦJ�Y�Z�:m�e���i֦EvX�U�vm:�z��WƯM��`�.ez��-P�_���o�e�i�]vZl�2Cڜ'�,�S��6#r��F�	k�Kv[l\���De��&�����뚄|�\��+�|+�t��+�BW'�^�&������$u������l�F���B��;	��݄G�6�'��8F�6#��x�Pa�iB��g	���	U6^ T�x�Pc�eB���u6^'��x��`�mB��wM6��f����6+#���Eh�Y��f̈́�����O�`��F���6�F����fA�&��	�6�M��4��f�Ľ>z�x�."��UJW#]Z�ta�e���b�[��j:�n���v:C�҅�$]F��E�*]Boa+Ĺ���O��w�<6��l/�gY��d7b�}���~!����b����O-&<]��B�3�Iϥ����\�i�-��s�cHx~���%�x�@*σ=y.���\@�t��d�"�?PK
    +Q�H$!�'/  i
  g  org/bridj/cpp/com/VARIANT$__VARIANT_NAME_1_union$__tagVARIANT$__VARIANT_NAME_3_union$__tagBRECORD.class  i
      /      �VmO�P~���mT&��Dن2�_�1 Y2�2?.�V��h���_���`��?G?���
̵��;���9�9'�����w �Xg�uc'^6�j-^�ۋW��x1S�e6��J%{U�ȼX+͗���k�6�.1�����Zv��*�1��l�F�bn�kJ��e�l�ٚ�/3̝5#=�]O����Q��s�/���o�0l_��"��E$����f�YR5�L3x#Ѣ�!`�A0ߨ�J��b�����nT�#�6ʗ����A!�m^Y���R��߷/כ��fUg�wPn3%�n��-�羈	�Ўbڄ:�lā��T�-K	w0�$�2���D/E�P���x�:ܲ�A� ���$9#�bi�t�t��Ҕ�!r��څ1���q ���Z�m�a�%%s-b~0��R�ax*-�E��^Uh�zE�eC��ue��H���)�ݲb؞�����fӠu�m:[r�����*E��ҹ���lR{���L���>����.gPfO��O���埢ݘN<w9*�Ν��n�M������RN�#[���	N��c�� �����~%�2���W��O�-���5�O����'��1
��@��c_p;�=��O(�6��~#e�,a�l/�����=mC)c�iA�`&����Hk��0���1�ܧ�Q�>���ɟ9��1�8mq�YN������Nb���A�w�_��&~N;�.�	����g#e:KHZ���	'�p藠���"��m�'y?������u��c�߸M��g�Z��Fv���� �q�l�VW�?�!�*�PK
    +Q�H�a-�  �^  Z  org/bridj/cpp/com/VARIANT$__VARIANT_NAME_1_union$__tagVARIANT$__VARIANT_NAME_3_union.class  �^      �      ͜{|�ǟ7��	0\�n�\�p��H����$9�ᜐ� hE�mUZ�[/m��k/�����jKuKkm�U����twe�+�]�>�eΙy�ygF��q��$3��~��w���y�?9��`>y���d_wUG_�ksUgooUgrkU[uKc��ճ���o�+�/�o��>��'x8���,�1y@e�[S}���ͱ�T�D�U�o�n�ה��&Uk���>iry�G�X{UǼ�/%pΐP�A�Q�ZV�lP�15-���-uy0�JG!��4�������E`�͇0�#Nm��hk�FZx���l��0���n��z�h��B�2�@N<I`l�܆��D`*���F`�z>f`�ݱTS2�ͤ	L.S�xc\�X�"��4f�l��V�gB�ߑ�}N+��)�
�T%�̆3��b��na��u1��#�yx���ҕ��R�%�'>��H�6m�E���x��y�Ln|��R�,�fKѬ�M��*��a��L����@5�P�Z
�&��m9y�����<������h˰��I/�zZ��x n��J�q����}� ��F�Z��jZk��7՞��V
`-��Y�G � n�J�n�6
�R�D6��,A�#h�IF� h�@'tQ�EАU��<4P� N�ڌ��2-4�ˠ�B��)���ǂPG!#0!�%:z�<uH� ��N)�e�~)+u�N���u%b�!#�ja���o��ny�d�C#�K� 94&�4��|�@ݮ����ߞ��FJ`|���%$Ј׊-,�k�F��+�;�Ӵ�<�o�＿�����Zg���jv��r�:�t�d'���]��p���E�+�����WԳ����JD��h��BY7�<�6�M���8�;�|o �П�ハ#�U�x"�c����C"�Ӄ�l�D�ax���(�-e.Yk:#��ԫ���%��qx����JՈ�Mt\�MtW�k�2t�D�"�͛b����� �a�7�w �%����|�|T��k[��,�!���3\�ﱁ�v��{�v!����h�s�X"\�W����Ѿ��N�="�vkuC}uKK�z���%��a������v��G��ۑ6?�C^�!q����������oxo<��*�z�j�-�@�w�Y������zoQ0=��h�����Wq�w�ػ�y�a����-����Md������@���A������)!�x"p��;md�;��������ӏu�#����'��1��_��>��5�t'~��������Sx�n�±�X?N�&��Dk��ɮe�$�K��Ԭ�����C
�+Ш������:�Q����B�bR[�1�@C@Ͼ�;ڻ2�;��������;uK[C={�)�Sh{�t3S�bi�yx{�u>��Τ�ۣ�͛J`^0u1V	e���K�r96���}��T�ķ1Z�*x��٥\��V�d�S���Fg�q>{5"g���KNG��t�G��r���4$�4�%l2D��S4��ϐO�@��"��K(�W�\�W�� ���J�*�7��*EP��<�B�GŬ�f�u���V7Y�U,��k�O��;���L����ihe��Q���>˂,$�,(���u��=����6r]<���e�T�0;�8�ϻ�\��:�%x �BFI3'l1�i�_���Z����{b����Q��/�!d5��ݚ��ʁ��>q��e ��o�����x�:�H�pZ�L��j�w'���>���6�u��9�w�Z�W�MB!kצO��U�Bw">s�]��(k@���KВ��1��4;�UYC�q���:0,�L>(,�U�:,]2��.��2��|~+2kPV�B���k)�w�k}n�=:k�N1	��|��t��(�m~��W�.��>�WR�G�����<+*�+���|��y:4k�:�����`����@���R
>u�t�_�8<�fu�\w�Y�����'�[}2�:k�������4������Ak�Q�䛳����5���!���[���Р��_��p�R�o�>áA[tp��!�ؒ�&kH;��J�z}g ��\��#�S�h��/0p����j2�|��=����&�:cq�q2ҘH��j{����~�9����z t[ ��ZtY`X����1���r�n��x� @v��( �8�<��a"FR�3 �b�+����A�s@Rɷ��#O��t� �>	���S�d���Cc�x�%Kanţi�"�H���ߊ�4�&�����ja��P%�^�l�F��_[r@�7��"�#���(�@� <��gp�%8��6��L֝C3=ۓ�)�_��_�ۘ�ĝ�9�,d�7��ߠ�28וŰA�����w��Z�$��¼V.9i=9,��$?���W-L� ��rx���r��d�?b���ͰʕA� ��g��EL�͕A.f���A3\lO���=D�0����vo�|.�<����a��~�(9�&��� o� l�dp�8�,FU�BBa��kg>��@�/A�Pt��20��G|��	�3��}�1g>��`\�Hr2X�Z���V�T�f�G<��g"��P�Z�N$�H0(`	���a(P ���ӼQh֋�P(4��ޤP(L�Y����H�( M��	_�[ܞ�[��Y�"�Ђ�{u�QX'gx��P��WJ�R�Юz��Uw
�{S�廐BE��Q0QH���45_
wHi^�v�&��N��d����.�&�-2>SP�3>�?�yT1Bq���=�c_������6*�[d���4\�����ݍ�>�?��ޥz��]���{�ݍ,½E��r�P0��dU
�+X̕r���A�����
*a��ih<?�t?�v�G��(� �y\�_����$<%�EK����k+ec;'��P���ƴy>�#	D�y!u�\����`ė�3
�g�YG!/!����n�݄��	>�MP66�#�W��5sHG�0�7�Եr���5}	R������ש�&��N���ecC1��P������@�$�>/����!8�a��ax�Q�	$xR�Au7�ew�?�&(�qNrs�����`N������K��B���;�)����~�gH����MP66��Hp��|UGpT ����r�d���|	��|_��T!�y��F�݄_�|ݛ�ll(Ƌ��ba�c��4<WH}Q��M��!h�|C!��ra+�|$�(ܿ����[w�o{���x%l�7a�;:��\'�n�k�'��!8ڗ�;
�w�w�B�H�C�Yu7��	��MP66�n$�I�����6!���a��c|	��|>pr�R�ߪ���{w�z���x7�F�Ř�:�c�#�n�k�#���K�B�(��f+d/�M�Uu7���	~�MP66�;��]��ksLGp\ �������ik��%xL!x��(d?< ��P�M�Ow�{���� �^��K�q��@���3��,�%x\!x\*�Y$���������_o������_�<�#8>�#:�'����x_�'�'�B^C����D�q%H�7A��P��B�og��	�~ ��o $Ĵ5'��K%�$���|��	����&�N0ϓ�bl(�#����x��,B0D4#	δ5�}	
A�١�� T�I��$��#�ecC1�!33��B���NRߔk��5'�,T���Bf"�Y��n��$��	��&(�q9�����1:��\(��k˴5'��C�9
Y������&)r'8���ll(�5H�V��ND�IH�/�0�ikN�%X�,&���A�m��۪�I&���MP66㋑�%��;x�DGpJ �1!�O�a����K�D!XB�;
I ��p@u7�w���	�Ɔb�B����x�TGpj ���ԃr�����T_��
�R2�Q��H���=��$e�+�	�Ɔb|�Y?�g*uK�]H�k�˴5K|	V*+�c�I�^$x�p?����tw��	�Ɔb�	> ��3��]$��\v���s_�4��.�b�4׭.vr�{QBO"��T�,t��By.f*��"������V��t��.*��r��a�m���nv�SX�܍z)�B�0ə��]���d�א��xd�na{F��퐼�,e����~�x�c�9�!R8�z��ׅmr�7Y�#�p�,Oo��(�t��R8.gX�4��uz��f@;���j��H�/��Ij\7��:�p�|8�a��S�k����p��a�Դ�Y�m��y��EP�z��<�����d��Ha
Y��P��l9����B�/�R�UHa��a�&w
��EHa1i֍�����ak�9�UL[3���e��Q��\�(�|�c��(#�*���>ʮ�eecC1^�������9�Z+ �:&ic��s|	�Q�q.'��H�Z��1��$k�	��&(�q7�V@v�:�e�Z+ �:&��ik��ܠ��\N_��y�Mr�;�K�	�Ɔb�	Z+ {�L��`y ��
���\ƴ5�}	�+۝�0�{���";Ew�D�	vz����N$h���o�]:��Z+ �:&�TH��w����]����~$h�����n���7y���� �V@���D�i]�̴5+}	��q�)��_Ե��Hp�;���ecC1~		�lk�	����RG0ɴ5��L(R!o!��u�H�ם`�7A��P��E������n\=�m\5}7��?������`y�@|��p�d����a$�4��0�IP�\��PK
    +Q�HĔHHQ  �	  C  org/bridj/cpp/com/VARIANT$__VARIANT_NAME_1_union$__tagVARIANT.class  �	      Q      �UMS�P=�~њ�U�"~���*�
����u�2�]�SM�:�F�q�ݸх�t�3θp\���K"Ĥ�.���w޹�w������a�d�Ѝ�̢�VV2���3e}5S������R�y*峷fJå����Me�Y��1toPL�^6o/��A�Ar��+JCa��j�zZ��7�J��R�jՋ��
��
�
�㪦�W����]�C	�����&���4���0-�C�E�hZfV��
AB�Z�:q^���G��=&� z���A�=��3ė�YX���f8��1ه?�(H8����õTa��^��j]� �>����)F��f��? �I�K�?Fݞa�=��5n4xeX�D#�s##�H���n�� w��#6X���`Y�n�l�Gm0���;EwSm��bjǄ� �g^1���s��79V׊{'��Ud�����)��i����R-*��,V���1�S5���.r�����5S]�E��R"�i�I̺FH��׍2�UP�i7��J��k�#ׂb����>-�OӛL�Q��a�qD���d'�]g��%"�GkItӻ 8�������P:���<,1K��,�:�w��>����cQ�;��TD�l��5�ҟ�I��5�T<%1@�7Dju��8�}��ڙ&��wz?y�;��;}�&uQ��`�����W`Ƣl�ApK="S|�/��PsF6��K���xF���my��+�E�܃Ж��/(���H�|s.n�u�2�-<o˃7^��,�����`�#�-�w�	\n����x��S(3�+����qKpdS?��!��W�$m�am!G� �F���_7B�(�t��Y�PK
    +Q�H�;��  M  6  org/bridj/cpp/com/VARIANT$__VARIANT_NAME_1_union.class  M            �R�n�@=��i��6�� 
�p	mx0 Y����TJKԷh��Fκr�|H$�|b�X4$A(�vf|f��m�����1���~���ޠ�\\�oXo�-�l��v:��i�Ǉ��N���40��˨����;N�!͠'Q�|�6�˻\�����`(�3��2,���zق	x�w�*�Fr�����t���Q��<2Xe��a�^6%��6��g0+ե��*ޘ��n��옻�H�V���Æ=�#���q��p��4��p��"h�@��d�q
�����oX�mMGR�;���6�є{�is�a{��6�c�6���ב���6��z�Z�=��m�K�u�Y$Vm�D3v�� �V�9m9��Jy��)Zn��}G��n)%���G#1��)Mi*=����4#��}��'2R���' �Q"]��'`�;�]��G/cB�X��[����@��Qq�(#-�H�ޤ�e�:��x��5�>�?��,�.�<�òxJ�DV
W�B_�,�t-	��PK
    +Q�H=:]��  �    org/bridj/cpp/com/VARIANT.class  �      �      �T�N�@=��`�R�R�.��@�PB�i
U�$@�c�8Vj��qP?��*��P��U����(	F�/w�w�{������'�52L�VU.[z�\V�uY5/�b�$�)�	`c��m5U��|����0��mL�+�
�x�߫�|�4l�BK3D/�ZSc��w6��Wo%3_*y�R!stPZ+5�4���k�]���=��x�s�k�Q������bQ��2�44��r���t��uNKx�a!<d�؟��T�v��N|RJ��u���b�R�$�v<  � �0-b
3C��2l1�喈�h�9u�VI�Ʌ`�&�H��j�c"3��^R�9	ֹ.`�
��]Pl�Rset�R�@O���ܬ�v�H��c��Pmya�����`�;*$�@�ʮ2|�����9l�H�&U7����}H{6��ѷ&�*�0�f���}ڬ�M��*�U�n;����(��d͊Ɵ��*��b�J�����0��	�yQ�,/3����7tJdô�JoMl���f�R�C�WI9�ЬlMi4��R�wz�x�)���{ʇh�K|�Pb�
#��go(��K����q*��| ������t�M��h�rPNr��[�Mk�� � �1�%  �d��	��w��N�?�/�+,�������[爌�brxF�
�](��I):G�~�^�r,�t���8�8vC`g��&^v!��n�Cu���/���ݢ&�������o��w��(��g��Ȓ���5����PK
    +Q�H�3�e�  D  &  org/bridj/demangling/Demangler$1.class  D      �      �TMOQ=����(�"R��KJۦI���!Y�jھ�!�23EI\��O�u��&~�[��C���m��v1����}�{g���u~ �ÌaVS%S��*�HU]�ԣ�f$�c�'jJ���V鐗m��gB�jk��<p1��$C��0�m����b�K{+���Ɗ������ �:U�'�Q��\o5��iB�������c#^80����y >(2(��F�s�*H��P��mb��h����Zu����+�<�b�iֆ�lU�9C�������}?���&n10j�lZ�j�t.h`M�2C���n!��3�]U1�kV�w��6��?��#�ٚ���M��$�j��>^%� ��!Ű�U@�'��OY7*�䱢QV�=��Ԓ�we�wS�Z;*q����vz�7ջ�U�j�L\!��-�Us��1�kݻ��#��1jf�?��%<eݰ������Qa�o��:%��HA]"�@@��19�	`�V�-S��F_<���}���)�)�vp�뙐<�)N�eI�s�r?�	���Ot&�f�"�\U���;L%��Rƕ�t}��[�']go���OvV�#���1C������Fp��:��,�yʚ@w)u/O�E�����ʕ(!�7E��/^��K�>E��^a�^�ʎ#Ѭg��oB���Z&C�����K\����f�n����:� C�B�~d	�5�:�Ő��PK
    +Q�H[�Ċl  �  &  org/bridj/demangling/Demangler$2.class  �      l      �T�n�@=��qskӤ�{[B��@MC�P[U�J���5���I�ԕk#۩�/ ��� ���G!f��y�����9ggg����� Vq��d�]�e�C�#�4�k�fW�70�]�* B�P;�T�}��֡h�
r@n�4-Wsu�tLf�[+��� ӄ����[�4X���ή!���n��+�L"���Fy��5� �I��-���m��d�����l!d�\�1Gg�@g	��CT�8��/��6ʿch����=~-U?�a���\L�<.$p	�	�&�Nsm��6�nnL!�;>�[8�I����&a1@���鹺1�����r�	�q�I.�E`�J�$�(Ʊ�a}��@Y�Ȏ��.�ԭ�f�k����''�l]7ţ�QK؞'w2��������55�g�]۪ml���epw%�	w�w'9���x���mq_�a�l��m�P�V��|`���C
��D���N���0�4��{��5��7^�|F�����
�&�I����9�����=ox�F�(���CH�?![���>�i$Dn��AHkW8]�K�[>�[�-%��*��M�%V�"y�?p�+��O��D�1"驜 z�U�v�R����8g���w6`�sbHEc PK
    +Q�HfD�  (  &  org/bridj/demangling/Demangler$3.class  (      �      �RMo�@}�8q�քR�RJ S�
a!ĩ!�����T����W����Zۅ��B�?����r�S���{�~of�_�~:�[��6�`d�hDr&����q�s�J�?�Ao*NE��FSf6ʄŋk��s�Ɵ�lT	[1��0j f�F���Ax�_�Y8�'>�s!�R����t�#Ԟ�|'Ξ���a����d/�*�5Fs�K��P�L	A�s���·]\E�A�\,�����gG����L���ӻ�f��V	�6Q�5o���&��[<��N~��}�G����	���7�M��:�95�:�H�X��<,6�R?N� �����8C��P�����$T:���e6���%�4]%�T�^�������,�Qd��
9��ʜ�X>���ʻ�[������sx�ae߲^�<M��&���
�&ǻ�.�M^�£�W��PA�����s�y5V��X�PK
    +Q�H��:�   �  0  org/bridj/demangling/Demangler$Annotations.class  �      �       �PMK1}�֮���gO��A� �RXA��[�K�5I�����*fW�-Tl ɼy3o���p�c�en13j��H�dJ'��7dsk�;�T�m"R��"�x��<w!�����	g�ˆh:ڄÄ]� �^<ף�3im4��ȪT�]�D�������wBk�-��0!ǣ���-��[M��	w���n��J{�/͜U�t��fS
���
�@q����6��
���t+��wPF�8�Q �A��PK
    +Q�H7�Ra�  6  -  org/bridj/demangling/Demangler$ClassRef.class  6      �      �V�sU���M�	�>h�j����6�
J[��P���Bi�<��mغٴ�-�" |�_,:0��q��`���t���sw�m�"u2�{����s���ϯO ��m���L2:���фHif���dt����.C�f��1������Ԅ�e9Æyr�vAc��|e^յ�P_�UOB��
���2�΅�.�HM�%:3I���kw�f��,=mfU��v�!RD�OK��w���(�0�f�HgIIb��]�턄� �PL�F����[1�PQ/�Jh��CC��Z?��5>��%�:��b��
E�'�5��}L		��`�l��A�ѣV�t��t#!2�#�UY������2�^ ���Oy�`�en!�ͫ�S!���	a&j�]�@��hD���թτ�ge����q�HvZ}��U���r���^�0TXݜKQ٨&M'���D���^GCI�Rt,��q^$����-jMNU��	����I}E(6�P�P��=N�#tP;�'C�x�MDyvYE�<�r.6a����NJ���~���3��Q��^�r�������T�'�mÅ����"G1臊cUn�4#'�\J�0C�5'=ۙ��IS5Dw&�"�eB#��)?Fpz�����c� kgvP�L}2'��M�E5�(2�yC�R[�@è�@���q��ַ�� $YŘsFt�Î���59r>��Х�q���
�Q�<=y�H�K�*�tl�I:���
N N"����@�;p�j�ݣ�=Eg���|�B+U-�gG8F"��L�5F.?�\ ��4mf��vh�]V�Jt|��r�	�ەN�F�q��2��A�����MїK���KٴX�Rq���\&.�u��1�P�CY�L�Q�ӧ�~4��+����}Cwڋ��Noݶ�?��p�l����������;i���7�|
��'*�%�M� �J2�y��d�r��#\^�G��j^�4*x͒	?¶Gx-�ׇk�a:��ϐ�1�Gq_���T+՞�����6o��)�;�Π���G�;o�H�y�=\����k�:g�6���uw�]�]?���e0�ftb�� ���=��8@;Q�z�%x8��C�"��5��TZ'��P�O����n~�\�a>���	Lr�)>�K\�U>��������<�{$�#��O<�<G>�E�[�(�ҧG���D�!���@��§���\��^Y�����Χ��)��{����+D���/�5z:��_$�Ef1���'Y�_y�)�3�T�Y$f����4��۔0��l��(�PV��x��Q���d��^c���b��I�C���^L�#�������T�6�
�<��F�H]$)�v����M��[X�o����m�+t�oH�f��*����'�Z���*d��S�t�l�H�>XR���B)��^7l�������w��w����-[߃�im%j�RE~�Xyk�����XE�ׇ
Z+i����� PK
    +Q�H 9)�  �  -  org/bridj/demangling/Demangler$Constant.class  �      �      �Q�n�@=�q��4)Mʣ-��
�AHQPRH���n��RG����~��H,� >
q���X̝��s�=���� �� RSo���̛���i�˩�4s���G2N�LL0���_p/���r4c��'"<x"zjjb���,=�x;0Qf(d5_O�(�OLT��E�q�.x0��W�2���O�04ۿ��!C��m4p��"6m��n��C19������f�<���W<d���sZnѮsJ��s�X���M�ң��m���:�F��$:Nu0l��e����Ş&�'���$>�`ȕ�G�8цa}�K�b��Zd*��\�ő����B��"�]R�Z���-�������à��~D��|��;���ne\�u �4��5QG�h�24Z7���Ua��ݹ��7K�;Ya	iQ��gѰ��K���M����ݺ��A/q�������[Tw�.�[�mO��M�JɢN���PK
    +Q�H<��>  0  8  org/bridj/demangling/Demangler$DemanglingException.class  0            �Q�nQ]�K�(B[��QQ�:m�O5��j�!��i�� '�4���|�F�-�&~�e�g �B_���>k������ la����=�����}��9��Y��V�����ٻ���sS B��~c[c�9 N�O�n���b���m�a)<�Ae���s���#���1�q�r���A�3�[;"���{�&�Ǿ��n;�ɲ�����za��y9�}���th�X!��E���UѮ����e\���@�]BӘ��hB�z�qCQ�$�tC�z������-V	B?��(e��B�ZK�BH�ޘ��b̲3�}T�A0�Z���!�:!ٱ�� �������Pz�9�}�懪�[������'����\�C���
ϱ�@��+T(�𹋁�H��ŧ'����6�a�k���u��<G���+�ĳ-����}��r�s)5ӬǪ���#\k�b��s��]���r�Zs�ƙ��0�z�DOuMl0�����'$�5|a|;bH�A��"�J��PK
    +Q�H��Y  \  4  org/bridj/demangling/Demangler$FunctionTypeRef.class  \      Y      �T]Sg~�l`I\SJ��Tm���5��P�@��p��&y	K7���Mg�W�^q��(u��Eo�����:}��"c/��:�<�9_���? ��{�ϯ*�]�)�d�r����ZG�_,5�jh{�_~�w�!p��M[Wl?��X?[��k�Q�~d�/0�nm�����!�fK�녖2	t':�6��V�L����P�_�];\�ν�Y~C@��7d0�FƩ�H n��6��P.Hf�.���coٲ�n5���\Y��Шp7�	q�i;5�7�ǊDE ��^����*57ykXau[��J�?_n9��b�p:
S��`0�pٱO�F�\4�1.���%�́�e�q*V�G�����3�v�vݵ*�,�^C`$���40�+i��~��������N#�U7-��:����nE2��|��T`�%+e�a�&�m�5W�#��R'�5|�@?8wT�b=�|�����L�8.͌�ꜝ+�����#��Y0�r�+H�W#N������^�AU��ۚ����s�q.{5ƙ){U�ٰ|[���Z�eە�M5�����j�!��zM�*K���.�!�,�4��?�5�$�|�u���	�i�w��S�0�o	|�u�%A�����y�=ER{�����gp6�����Pįm���K+�s�X%p��D�گ^�?�^�d����>���c\^���0s}��c\����d6����1�MKm-�z�e��jb_F^M,���ޤ~��-��S�ܠVK�D��6ΒAS�^`P{�amY�Ƶ�1��C}�5�<�]yP����A��{�� �ה�EZ}X�>I:��ϑ�w��I~��)JRJ��PK
    +Q�Hi��C�  �  *  org/bridj/demangling/Demangler$Ident.class  �      �      �SKOQ�n�>yU
�)�t�P)X���h}DJIL�tR�S���M�nLܸa���ф�ƅ���D=�-��׹�|�;߹����] c�e,عh�6��Ѭ�׬�iX����V���Ur�1��kϴ�I���̺�FV� �&>e<�]p24�/F�rB����0��~�ι�f����^߁ g���΄�[4�C����H.,��Z��(�)��0��:=[�hH�Q"���)K6%�+�����g�BB��h����~�" v�R�AD�N®H����/��?-k&��ʄ�~��Op�g`��٨��,w�P�ch���%�8l�+fV4P�BE;��66t+K�G�f->��FD�ʫBP���m�^��1�H�1ļ�a�a}���0��
D��/d+o����˚mhS_Csʰ�;�|F�k�b�l���q�/X�nϛZ���O��@r�
�t���f��� ��v�N+������E�BH�l����Ls_���]i��� t A� ���exxM\!�y-�wBqҚV�«~��%�|S��m�=B���ܵ;s�+a�q)(u�F��	J�Hu��!�7�~H�u��)��Ǡ`�t�{H
70D6�&�a��*�h�*F��Q4�|}||2����8O"�gp���>��9B��*}D�B��OPWvI�J���Ħ�&�m���ٶW�k�t��a�zn��V~!~����Xfh�$�zf��1������CS��7PK
    +Q�H��߭�   �   .  org/bridj/demangling/Demangler$IdentLike.class  �       �       ;�o�>CnF���t���̔,����ļ��̼t}3�H�3%5��'3;�����A +�,Q?(���\������W��gd��o(;#'�dF���Ң�T�� ��3//��9'��8�������8�$+��b ɱ3p�q PK
    +Q�H��$V  R	  0  org/bridj/demangling/Demangler$JavaTypeRef.class  R	      V      �T]SU~�IH���+��H	�V�(HiA0Z�ŏM���l6��t�{�^:���3�qҎ�t�������>g�Ib!-^���s�}��9��������}������3s�9��Z����,gxU�o}~h�5�#��W��@KU<q@����8Sw��[���f�.�u�@ P�Q]��ґ�E�c�[FڍK�-�zˎ{u�EK/�:&���Ij�3s4�Ϛ���	(��m�AE�t���b��W�tmYýS�-s�42kz��]��9��:4�Q4�����6Ti8�� ��_&]*Z�W�4i����:�!0 ���� ����а3��}>����kx=��)�pC$�5l�1�D��+������0�W���fFɩ1[��˖@�T�*����e�&���r=u@� �d���X]�v�Ӗ�]����Nr�j�D��0Ŧ��ٸ%�~����Zoc��Z�y�veqfZ_�	�]�f
3k�)�Xr�9���1v�ػXa7H���e�^�̷���"����B*c��[�JK��zS�&���u��/�O�CT7��r��T�0M�ѻ4��M���Y6ܦ�;�9�����]��ŗO͖$�@CB�\FR~&��b��ÉRY(9X+t��!�)��>�b>í#�O�ֶ���2'L�X+�R�S����p+��f�褍%S~h+6'�K�Q�?M|��E��1t|�I۩����)%qo�	��� :W�,Dz����KI�_\����Htt��{���x\�*�*�4�K��F���>�:�h��OJ}ܓe��Z�˴V�O}4V��Ƶ��GR�3�@�>^����.u�Gy		�1I6.�b������5U�^΄wj�{t��X�5�[��ϓ�4�=U�jU�J�iA^��Y�E�S	�[iưĈ�aY!^i�=�Jȿ���}�'\�y���ݸ{6�L��ꅯ0�V�L��a_	��s�P	��/T���^������g��!�QD'�%�<��=ǻ�.��1�K��i�{���Nv��<�^ګ�[��+-R�X%���_F��0�^*}��>��#��#w�k�� c�e8�� 45�PK
    +Q�H.^�  �'  .  org/bridj/demangling/Demangler$MemberRef.class  �'      �      �Y	|���?���d�AB �� sE��pE�B��#�̄�I�ŻoTh-n-�1�-�j�u�v��W������Z��۵�����Lf�I&���e��=���?��<o�S Ηg��X{��X�mGu�����C������+i4;���u�vD��#��s�z�fk�����9z]0;��{�L��[0m���	<An��mf$��iz0Z�M�0��]�`�\k��,�贉��H��.�!�P4RҜ��i������x�am$��FscZ�DA�"��$bJ��M��e����5�N�;��i�ssP~<���Sy}�Ѕ��e�bM��9�.�`��d$�����zc�ݝ|�7'��;�C�R����ZI��fl�`�iG������02?%��'�6m2_�eA[��x�\�\�Bd"Ԛ�pY46�n�7Ţ	���C�(�C�{g�-�=d�hx�'��`,ةq�l��%�%:b���D���JT�f�OD��Z�a����i���dH(�X�*-k�c!����Jt��#Pl*��lB�L�,�y�_I��"\��(,����Y|���,�w�Q�2M��;��)'�f!,k!��`��Ì���Ϣ��1s{�~Q���mb.&��6BG�c�����^LO++�>5���֡�/�3;�	V����.��G6���״�X�O�3��9�%Kt���¦U��v񵬴���`��P��[�(BЏ4jm2��ì��nMDc�ڡ�<�FiYztڄ���t�~�݉P�zxQ�`��oX�WP1�9���(�Nv�!<13���ă.���P�1:^RF�+�?��~���"��}��G0uX�xp�`�l҉�L�����Ҳ͛Gpܵ���\G�!�UfČ�ZS,�4YDfCiяp�fq�TH�miPS��k�ogn��f����qnն�ǻκ}h�L}F����.��8���C�KJ�D=���(��[��|�j�#��/,_̈��C>��(���L���R�V֠]lRvn���1i��c����f���~���0U���[�P�.!2Tl���HG�/�FWX:�L��	<���)^�L%2��;n��X���g��\���
�G��4�l��,����6����Ti� �+r�F�����DG���N'jՃ}�.n�?Q?�K��:ۏ�:Yy�52�^��e
����~|�zы������?��Gza\�6%��Ռ��ʰ�r9��5*.�n��q�,���r�����������F�fئh���P���M��1ϋ��Gize8d��/~��M��G����O���*Z�G���y�^�&O���:�/��K�Z����=���i��u���۲~��o4���o	������#uk׬r�����{u%�ރ_�v��R�����/�ׇ:���u7W�ؿ���������h�*�Ћ�,�T�{���i��&��C�]4��E;uj��~�~������t��c�5пɀ����z�[�ξ��E�n3*�]���ͼ>��|�|�a�:g��$ w�z\˶�z$Y����.(��/�����+���f3�v�g�3t�\qM��eu��n~R��1�W˺C�6:��|2Z� �5�b�EqG0�6ۊk��da���[��t�6���"�����|�v���n�&�����2�&�BVQ��=�I�$�����d����>�Jse��r�H.-o��c�Fľ�ݝV�6�N�ܝ �p�K7l�sx��l��s�5k�Mt�L��ڋe�u��8�ͶaSw4_��
fi���P����pP+�)OǗf)Ce�T3��yvU���e�Z��/s�J\.���ŝ�^O�B��V?Vb���"ݏG-vi�.��/����^Y�7}GoZl#hL��+s7Y�=�_��R�h�[�>67m�ۜ�,��=W�J��UI�^��ns[j�2�r�4��fK���؍�����3�{�r[���u���|԰A��)LT�'҂z��A��{1MX�V�`A���<�+�*m֫M�#�'��n�*2��0���hw{Gq�qV�{���u@BɂtpB1uB`5XJ�z1kb��	1��lY�t�]�G]A�r:v�G	�Mט�2��u*\��)tn�ڮݴki��B��B^�G�Mr�`~I��SHc�K�+� ��C,��+S�͌���z/J���h�-	��r���"���ٟ�f�(���V������2�:L}�_n�n8[菃�}�����+/S�,50s��)����mF�ͨ�nV�Ƚ��}4�66)C2`��0c�D¤auP��gf���0����䏧�����"M���I�E�L�ND[��fu]9R�6�"�n֙�����o�.,�?~'э�n�Fԏ��m�z��hw��\�8������q�`[� ��,E�F�(���γ
s��U�<�y��k=`��d���ZO菐ָ�,��B,�ȣ/]�F�˸��ŷaMb	���q����:���P�/&�Qz���%�觞h���֛� ��C̓��/�A@N��Ŝ@.�兩,���hݦYH ���4:��ನ��'q�Lԏ��^lH�C�cP��N��:a
6a�s��t	�_���� �L1�>�mG1��"���8ONq�<��rr6���5�Ϩ%�-6��s0\�-އ�%��Jb�i�ZS������7����_�.U�z�1����;�����-j�q�,\��SR�Zl\��=���g����c}��x�8�q.���8���=�-O��)�Z�9M�Vç��W��1Q5a��ej��z�W�N�`��B��4����PZ~����p ��qG�_r���U单��jT��z���jn�QQ��O�x\5y�y��#�p�ͭ��#���َ�˓c_��O����_��ɶ��8�g��$:�s8JS��cT��Q�o�-�����Q����m>u��}.�/���t�
ǹ
���K��d��z�g�k��=M�W��m�R��P��b�_¹��Q��<�5���Q�xz�s�k!��D#�����<Uc�B�,�
�ER+�^9
�>Q�d��:��*�?O�逧gcL�[��!��N������O��cM��9~�Gf���3=�sk$�pF������4��������s��=�W=~������~��c�ݨcحG��1�p'��4|-��L��_��RKR���7^<���W�{�+2����?^�JJ�e"�I	�,S^�N��kE�N��j��2U��f��Nwqc���b���e������!3e�e�R�9�I���{�����LW*
mn�0.�<�x�
c��d�D�Q�����P�b8_��	�E7��n\��`�ڋ�:t��q��7�q��	w�����[�ڇ�~�T��G�v���u�Uw��� �Sw�}u7>U��su���}2M�/e��V�Z��J�"�8ѾՉ�):�_C�!'�ɹ���ʇ�ؖ�l矨��c�y�?� x���j�!u�1��bh�|S�tE�T��1�3�T�uSp:��2�V���@��i�g��&�Bg��|F�(��뤆Nd]z!M�,��:с�Mxշ0��9_�@��A�z3���*O2M&	�����6}���\|��#)����'-M%�κ�.)�9�:)�����3���Y�K!틅�����X�Þ?'jU�Ii9�i�TF�s�T�WJƍ����)E�w��[C�#����moE%�=b+b.=��b�z�w�iz��T���&Z�[ج�FP����Oq�z����A'qR!:�2�F�jt��F��_Oո�B�l*T�����Zhle��˅��ڼ@�k��؀� �j��q=7�y@��d �4����Iٲ�<�^�q��>���9�HiI)-�#/I���Q�
�#��@�V)����󽲭�}|Ok�'15�ZژRh�v��^ٹ�R�`|�1�=8;��N�	�a	��f&����2��%]��&�j٥�pzd	�Up����c���lp�D���*N��ˀb�i��p�D�����Љ�2o�Ҽ��>�t�f��Q�>�y�WL>�a��5.S�A��-6�ϱ]}���v�/�iч�102�x���YÇ��x�����X����x���	�ȘD�$��)�����iG�4H��_��=]�8�{[��^No�ȟ�R�h�	�QN�()�������:8���7h:��i�8)���;4C�h�a�+4����^��"�4�L;G��Ϙ����6`G�y8$��y�d���Sg-cz�1y�4L4�c�Q����3Qm���F	���n�b�Q����hT�1��1�7�<,�d�����}LZn\����Y���:g3`,$�7�P �3�X�YB ��DzrYN��ف�H�  �	���ٛ`9by�!��E��q�S^�x1���X>��,`=Y�$��^B��M����Oz1�����ο��ɿ]3��a6�����PK
    +Q�H��i    1  org/bridj/demangling/Demangler$NamespaceRef.class              ��]OQ����nw��Z���P�Ѝ�X����&��n���f�m�[/�G�(M��(�쇅��bg��;�̙9�~�	�	LBs��H�o:b`��'}�|��"��Y1Y=�V� ��?
>����8���{��|}����ؒ��@�����:����|m�E/lrϥ/��J�
��%dj��EY��QР�!��1a���%W�o&�'��p"��v��~p�ˉ����3%��X��`��]1ޥ���f�pW��{��&,]s-��d�3��p�$j�p����U�h�Q�y��c%��x�����ΰgy]+��퉃��:�{��-�4��'AO���`��|�m��Ř�
?-@�����#��M�4��úi�3�ͯ(擂&�J�`@�E�&�E�@YAVY��T9�c��]�XE����r��7��4�>J�)��X��W�CV���"�[�I�}ƕQ^����3�eO�q��9�H��}��d}+κ�����*��x9*���PK
    +Q�H���|  =	  3  org/bridj/demangling/Demangler$PointerTypeRef.class  =	      |      �U�RG==��	��,6�b�A l�v��L,�X��x$5b@������?1���;�p��-�ʿ�R�=�hcH����v�sN�{��~��8����-=���f�򺑋OyKn�S�n8�Z�v�/�M���).������Bc��agMJ������pO��h�n�� C��@_�.\V�1�%�v�C{X�mn�0S����<��6��uCw�3��Ych苬�hC{ 2:T���	��"N�<��'�㜶,�B�@�8�������ӽ�Qׇ�.Ԛ��bQ��:��k
�H_�J��X����JlDN�bh#�A�{�L��U��<\��i��ܠ'M�L��\ �O)�i���Rr����a�9�����w<! ;�HYHo�s����")Qn��ǀ0wAs2[�23[j��<��E����p���-je�E1i9w�V�SӔ���<�,��=?��e�L�F<�P2Pq�v�,eq���1,!�!&�b�A�7q���?ᦑ����l 
Չ*����Z��(HRՒR��s�x�3�YP1�� �`�W�������@n��H骡�yJ��։C�����3]�nC�2VX�*C@�d�m����T|!�
�$�GkJ�F _�*�_�zև��yU��z$|�^(����*�r�!�sdDp;Z�IB��i�����T�ߩ��7�ɗ[^g�ۺų�>�L.E��n$oy��ɛ4�$/�43Z~M�t��1P����狅4�'�X6�V����C�3�����Uj{2�uI`��ݢu���,m�h��S:!��=Ĺ���GK��oѳ~��Dc������Kc�wq	pW�a��!�'C�F�)��t�v.�J�i�|hVb��K���z�3W@D%'���dɅo)A#u�2�{=��-�$w0�3zK��E�%�T)T�X��
��Fje��IH#�;�X�!�D�|{�ϾGkh�WLK�lo07z<PBj��{���ʂ�O�<OC�JȾDs������$ q�G�/��AE�G]��86]�;�a�N�1�H�nQ�7)��*���4�4����9\�#,%1 =A\Z���¼��ui	Ϥe<�V��6��W��L@[H)��/��	]"��&bC$�rE7¦�<ɑ)Q>Y��*��/H����PK
    +Q�H�,5  �  0  org/bridj/demangling/Demangler$SpecialName.class  �      5      ��y`U�o�$yI^���\M��h�ͱm�;G���M鶁�в�L�m7�aw�R� ��������S
�eEEDAE�R��*�a�7��n�M�?�3�����7�f�M�>t�� 0��$��ƶ�c���!s$�E��z����P �&0bf !��w{`<�c�[i���Z;Z?���!3���0[	L9�H�����3 +��f����{d�v��@f�"&��H<&�1��r�t�{D����N������N�1�f�%]c�̥;��ng,؅#�N�e�/_��V��J�����{��Q�o�@�?b���ߴ7&��􍚱 nv�㡭�X��N�O���xh�L�K��ѡ�pt���'���uW(�Jjå�R#�Kړ��Mm��H���PpM4�j�촱@8�*�6cx[(L:?6��]�@p����<t��.'u�b��N��V�����.W�U�`�q�>�9���qBAt٩�CC�������ݟ�gPΏKșq��7�ӌ�.����*�I�"fv���L�e�^wtd$ષ6`_�mf<?r��<d���Uę�'�9��#�ݨ��=����tE�o2�"�+Aw���>�xg����"�D(��F|*C���Ƞ}A2��;{7,�h�tl/���@x�ī⫫?��V�q����p>��p4�Cϯ�w�op;>��v-��}��7�9��^XZ7�4�m���%�Áx�u��G��q8�?��D<��P$���ej�Ѭ��6n���鞬q}?��d>�C,���f�a��u*��rk':�;Y"*{}�R�N���n��8Q�3�! v�ܘ�%G8���x�A.�\�c 8�3� �C��9���A�;�a``刹���i?� /А��g��2���ql��_�P ��
q���}�C�����Ȟ�ᄽH0��"�|�A����{�e�}S�0�z�\�a���2(�q%py�3�1����4��qg�)R�
n$��Z?�0M6��R��������P*����t\����mgp-��2���'4�ut0��a�odP�
}��fe2��A�+����e�;�z:\�?p���*]i[��P)ӿ0��*\��f����\�n���J��bP�
7c� �j>̠���1x�C�gP�D��P+��Թ:�c��8������×9���U^Wh�Xop���M���ƣ#fyW��d;��w84�f�1ht�h�	��C��à�5l/�����x4�:640�ơY�|�M�dq�ɐ3�媊>��d�����p�E�9̖Y!�9�ȝ�Z\s�ԁ�+��"������0Wf3�seՌ�p�'�:�]Y#�ˬ����32���a��ձ��y�l�E�g ;.�H�x�,vuldd	��2�d���XW�H�V.g���x&#�8���x�l3#k8��l-�W��?��m`���h�0r�%2��`������pX*�-:]��q�C��t�o�r�a�A��V�0̡[�����?�r{Cs͘����i�7����@,d�+���υ@b,��E��Er���G�bAsy���WE"f�Y#����xۧ�wa�ҩ����U�y������X�X�X�X�8U�Dq�b��t��e�����3��kk�������M�͊>�Y���(�(�U��8_q��B�E��[��;�(.U�T�R춉�������J����"�}���^�_z�*q��,�� �}�w-�r���} ۯ���\�3�Y��{��<v{��/��<�<����+�EP�m(�N�6�-�m/�i{!x]��4�9�eoٕ��e��L�Ks�V��,hҵ<��t��(��Iܩ����0��Ç{�hӼ�Ö�O!M��)h��w9l��s��O�\��+'����3�Cn�d��-8}v��-�зS=�i7Bd�:�4-%�H��ĸ#v���.G�����Y����َ��H׿��9����п��y���`���\��o�L��T��]��_��Ŏ����H�c.s̏�/W�
��T��?W��t�Ub�~�2�8��"W�N�=��^�enr�oD�~�2�9�v������1���Ge�r̟D�~�2�8毢@��2�9�~Q��S��oQ�?��#�yT���9��'�T�)e�q̳�D^�󒘦���k�y]���y�1o����ʼ���#e9�cQf"��2�&����.ST$[�馈J��t�1� �IW,��ׅ�H5MTd�reҕ��T*W%]��5H�r��yE�A�k��'�2[���
�A�+�P�E�� �ʵK�!�T�.�E�A�)�B���� �)�+�j�3H�r'H�N�2�z���;Q�6Ȁr��;Y�1�f�N�. ZTΔnX�5�6�K�C�3ȈrQ1�6�ԂQ��fA�?�f�� ݂]��v��g��s��C�� �i��|�_�ȶ�2��
D�W"�Xp"ׂ=a�M�<nC�܁0,��o�=��CZ� �ȂG�@L��D�/"�Y��Ԃ��-x1ÂC�2�PD�E��"9�J�舙)BTY�Qm�2D�E���G�Y�Qo���"iG4Z��d��f��"|91�"���ل�c�S-1s-�1�"Q�Xs]jM܏�8�!�>��ah��@}6��`�����p.= ��'��$�O���ix�>��g	�ϑ�<i�/��"YK_"��e����s��"����Nn�o�{�Ar��Iҷ<}�SH����w=��=O}��xv�=�я<��C�~�S���y(v���F�Z����:-�k���e��,z��Mo�8�[ˡ��)� ��T���1���#u���ʞ�_H���_PK
    +Q�H
+���    +  org/bridj/demangling/Demangler$Symbol.class        �      �W�{g~��e/J	X!@�	����p	��$$pvw�L�̦��	��7koڪ�&؊V������b[{�����ǟ�7||����f�!���3��}����=g�\���o��X�2�#1SO�FZ�jt'u�;�������'�b��B`~�:�F�܈��jqˋ�y��r_�f�mZ_L3�k]^����i/|��ɔ�aDv��Ͱ��Q�n�Hj^�X2�/�
��ʝ�6�xgn��x\�w-XXd�nӮ�`t�^��S[�j"aj鴀h(1eJ��[1:��d�j��]t�aR���yB�2�������E����s(z���hy�n�V�@C��fQ��ljj;��*�R�V������Q%�(�zt&�n��n'ЭY�l��jj��d9����rl��*X�J�."�W���(Z++�RZ~��HK��E4-B��J9��-�ޞѓ	���	����߯�x}��w�	i�����fO�Ƈm~������g'UV��.�p�\��Cɶ��Iz��ŸV"��f�ǋ=� �*��)�=��7؋���WZ�*����v]�ij�jR�;I;s��35���d8H�6�on�5Q�á)͉��w�Q}���f�֩�0�p+��l�e�W�J)(�1Fs.���RӖs��9B���EڗT�����N�郺�H:�e�cHЋ>���C���)�Ru#-�!ގ�l�n�hF\�A�S��9��rF�� �� �X/,����l6O�ɇ��:D�ԓ��������"m�ՓJ��&�s��9�G��
FM���(�w��=�l�23�ʱ���%;?0��*&˼��V/�AB�e����x?�$ڒ�����Р����T*��FBO���e��v����Dȝ(��ֻ�ʘ�.�4��!#e�l��-�g���GeL
�!<Nh�̄�F�;`�q&�L�N<eȚG;>���Q�xeę�`�Lу_	̱��PMEg��01����|6�����XJ��S�~�ݢ��t�RuY��,���ƆV�i���,A���A�4xZ��N�^�8�"_a��eG\�~��M+�&H��!��<I5��%[Q��Ř#�v��?�I�
�K��(h�l���wZ�,^�J|C~��Ơ�1�Mĺ`�5{3m����b7n�1\��<K;59l�NY�g�^����{���W��(��@�g�@������^�S����g��r�Բ�
>r��1�z��;R	M^�Rq���ew�"�ڞ�T���x�1f�n�۳���4�H첰[����}�=�1��.]�Tv�f���4���-�U���u
��������.�s��d�푗���=�|���z	���׍am�~5gl��|��m�"l;���	��t�����`�f��-��F�M<S�z7L�oiS>��Ws�g�u���W�6>ף���u���y=61�8��n>�����ݸ��M9�.VN�k|7:����8�d�6�`����%x�c��,��8-�~>[�7�^� �U�[���aò�N��1����
�V�9�'�$� ��C�?�o�Λ�'�P^IO�Y̷���H��Da���^��(G�ґ��2ץ�QI�EtH���q|wsã��a���U-��c��'`Q�r�����1���9�s��}�4�.�°���<=�2��I:���n��h^6�D^��B��Jt�Vt�B߃ыVq���$:D��E�¤^0���嶕.Q�M�G�9����Dz�d�n���q<�u�0n��Cؐ���=H�������&-T��8���|m��*9���p1��DÔB5o�Ü������]s=ǔ���˔�� [w���X$��2q���h�స��x��qq?o��2���Mn���)jןW_Gs^<BFxEs����I��tpj-y����ACԮ��U��(�BU�f/8�y�i�	�z0\:�Sg��KAVrFM�u)���Wk�0�A<J��b�4*�X*�DH<�B#,N�/�g�[������g�<�s<%��s��`�e�M����B�Wc/�I�&��������r���[.�kI���̿H�_&�0����j�(��9|n�����w��aL���B�`:��6vb�(��Y?	��p��\k]�%vE��#��'t��<��\��~��4&��kL�M��6�xk��L�]��{X/>p����]��Q�!�_"����b�L
� �����<
�����zW{�*<�4���k�w��w�W����N��h�䞟�?�ŏ��PK
    +Q�H6`��   v  0  org/bridj/demangling/Demangler$TemplateArg.class  v      �       ���JA��Ժ�Z��Ƀzp���b
�
z�nú��̌>�����
R<TsH�������;�k�	�]��2ԫƮ�e_��Wv����}v������u��Ų�2�F?��������.q�;2���{��pˤ�V2�a˩|�xǁ[Bq>��s2����#ap߽�Rnk'�潄�1JԼ=��)꫆#�F_}�:O�r�\)�0��PK
    +Q�H���+  �
  ,  org/bridj/demangling/Demangler$TypeRef.class  �
      +      �U�sU�}�&��[�
�]LӖ��bZ���\-�x�$�a�f6�~�U���q�A_ꌃO���E|���8�wv�$4-��d�����w����/��	�N1�s��d� J�]�L����/������8,&TaѤq��X,��M���"LH�΃(U,�CNQE���!�$�V�ځ�A�}�!�.��k��BG��dC�����$�S=�bQ
��{�d��蝡3���{�fX�)
cFI��F��q6��VA8'z�������yLT,O@G����N ����[�uKRsx�p/VI�ՌmQ��1�:AUs��i%�͟Ճ�c�C�U���l--���M����EF"��~�.G���U�.�i�AZ��K�T�*��E0Y�V���Mًe2���!��mU��;o�}��ؚ̓@�|7ޮϮ�;r�h���.�<r�)��*�֨8��J��C!1ہ�	�Q�a(#өV�<�k��pV	*v:9�&:����J[�niZq�ao{���`���i�(dƭ��6���	��$1�'t�)�8��ߕ5h8$��AfZ�5��Ū�)��l6�1>$�b8�)8�I^Ya{�Qhߙ�1����Y9t���y�� ^��X�.����4�!��X`T*��E�q�-&P���]3yc��\�b�9F�u�c��"gje��xGQؽ�r%Tf�膉w�Y�Laʜ���5&��2�	��c��o<���w�gk�l^�w�vW�8��Y����G��A*�{�Ge��cД�傐���5n8����Q�`������r�	v�oV�dA�H����^S~h#6a/9QU���P���k:�o����e�̈́F$}��x�����M,�~����UH�
�-��''��"�%��W�be��J�P��X�i��_3�,Wk���t�o=6���&G�;t��,��HǂHz��HMaq��R�o
�2%|yV �HG?6ye�\�� �_���!���2βK�p��� ��{e]��l6үG��5��rYW��u<~�٨��j]�ct��XV��zﳎ#�[�~�q����u<W��Uu��`'7L)7e�����Y�܎]�_R��%��ʮ�C���,T�5V\N�Kx�<(.PD�1γ^IL�%��t��^�k\��x��
����]{�W1��ŷ����1��Q�		���$�
�~�:��l�?�&�;�o�p���qt�g��� C��P����o���8㐌���^�s3����e�j5��5���P�5���U��q0��8J�����Y3����PK
    +Q�H�9���  �9  $  org/bridj/demangling/Demangler.class  �9      �      �Z	xT�>��L&3 d���0I�ʦc�A@-��'3qf�`�j醥U���*H��J Q�Z��պ�j����mݺ������f&�0��_��w�s���s��8ND��"������h�y}e����k+�M#�&f�]�������FS�M�����2�TrrRc��)��4ì:��ш.5Zܔ��_��V6�M�@hI��pSSNR��������Hx٦6Cs��4�['��T�C�XL/Ȕ���4&ú�f#�0�t3������Őu�d�f��ٰ�-��)���"���H07�6�����>��4�"��@�I��ɗ��-G±x@6Z�l�1�˰�=��m��ɯ6�6FBn���e�3�x���
čyѵn*���:�&gX���\���htS%S~����#�̍�i2�$ud���n��y��n���ţLy��|��b�,h.d����1qL��M��P�1�nb*�M�Xt�Zs��� ����� 4��f�Z��lA��tu:�	˱2ћ��)I�aS,n��i$��Ï
MZ�He=�A�����YT��t6Ӡ���C͒/k!��`8�j���h	��:�Gl/���̒lZ�9��6#!*J{ ��e��et�P�h#{�	X$e���J{UlO*�����V�S�ј����j����B�H�|�����AĀ��G�G�A����%��L��m�t����s�IG^Rؓ�!�z��KA����Ł���E��|�-�L���z����Q=*B&$)?�8��(Am�JuG��# i��F�@�\� ��=q-B7'���)!��L����LJ�9�/$��|�K3����yӢd[D����Rr�,H�n�C������F\o�ؑN�-1�'é�D[��E��iiO�,�F�ъm����*��%E_A�v=�7d���][�/U��Pi�e���T�94� ���'h��:R��=7}Sg�͢[�t�&-�r������	���ʆ�A���t�u��eZ�zR2d��jI�9MPU{�!ݚ{���ҝ��������	�%��n�a��'O*�J����_^�i7�0����F�������I���ESU�O��Zz n?S�y�M����`��H��#]&��=/l�w?����)�;^z��='	�a5H�>�2]�.M�N�է�A�����ݳGj����4��>�@���iUﰒjPjJpJ�|�$=#��l�(�F���(b���_��EN:7������8RQi��5V?���^ɡӫ]TR���SXj] ���׮��G��9�3�9�,��SwC��ޤ_ʼ�0OdH��l	
z�������M,H�>��������bӁ��5��л�������>�@�n�?`N�v���pu�����F�ib ���@L�G|��L�J3��ފ�zi������i�rJɩ'�db+}��G�z����M��B�ȥF��._��O��>����ǣ���nX�q���l�⁄0N�b��E��CF�~LC�_l�ShI ^�U��d� I�5'M�<P�1�ȏ#�B��E���'��C�8�r��d�A���H�u��i�4'������jP�T�K�Itpod�<�d����2�i�C2��k��^�r
A���R���!ӵ!jGO9<�qz�j���ޥ�ԠUQP�.F}]Ő���>D��r&��.�SS4��L�P���*/O�c΀n:q�'�<S��5�.d�B��g�)��$�f+�[3LS9vH�]�
��x2O/�IoP�>�U����bѯ�93[Υ<1�?�!j��d��D0������3���<>c�В0��zS�͒�W�ZEW�}���\�tM�eq_��_��
�s~��B�&1�)H]z̬�!��L����R|��`���|�x�ELUitf�e{�ݼt ^�R�Ϡ�=4T�����3��@{(�߀;/3��[S{�^u`Zr��[x�"��u��z�LB��J �#�Ғng��o�?�C<��h���٩��������%^*d8����oa�Uq/�q;S�)q�s|��]��y�<�o���bY"�N����rX�.5-=$�FMq!_�W��|u��}�l|���n�Y=�\�zsQ4�*uoz���f���#�G�-;tS�=F�h�x!���	�z����_8[��$��Ⱦkll_���le�B��{x+�ǟ�;��3�J���%}Z3���� @��#�m�0�ɠ�oe��_wӋ0V�@�&g� ��^��hk ���}�ڻ�����ϚQ˺��r� �(W���P����v��Ƿ𭢍oa�
���֠�3�x�!�ٝR,
Eq7��{��)7"�r��<�O��'��o�c��+I׺R;pf��x���&�jX����>ԍ`m$��͇=|D��>?	�����n��G����qP����䪃r���Q�YF�����Ni>~*�K��r>ʂ�P��5j׹Q�]>�%'?�:N`/�'���?�
�'�)���d�QNݮ�U�������?#��j1���5�>k��uxG�5�/�5>~�_�/�rE�$���07��+O�($SH���4�g`��e7���P�
�4��?�7S�I�YǼ�ZȺ6�����������¿�x�j3�~�&D����{+�5�Z+��������,I�˂�������\ۻ]�Aq���8GL�W�r������<�{5����d�������G>�'�K���&�xAyI�"D[���Y<.���pz3i�$�؈���M!�CUQ�F�f�D� ��c>���[e�L��9̫�4B�Ѡl���֫��%�������
�S��z�fyds���O��O���v-O����+�O��ښ���(�k<=^���!�<n{"��&cQP�	�~ѣF�9�9��E���0��S>-���tQ�`�@�{)yh>U+/P�m�ז��;|�N
��<�y�>y��V�s�:i�1Z������NZ�IM����Z��w����ImIӣzzܜ��Iz����{>�� ��* _t��S��9�ܐ�E��F���[�"�9�X���ӈ1���UaM��@�!ѕ%�C{"	�UX}�}
�.���3 ����M��vj�����M�Pc<=�h�J�a��~�� }� m��Y��tO�&�y��d�Io��}�}���l���OY�y�~k:�*pc:���[�,�~A����I�[�L�a�Jt4��w����h��������e��[l.%�\��v�x���Ҝ�h?�nw ѷ�?�"�G�0w7�l�����Oۺ��2�$�r���^����/�+?>�Q�,t�I��S�\�N�W�U�U��Ne�.o��X�;�w����u-�G��#>�Vo@>@ǀ���уh���:��Cx��l�nXn�v7	�z[=�t�8I)A�>�六t�j�~I2�fzؖ�����4sʖT�r:�\��B�N*�(tM��V����6� �m[�G!T�:�G���3���)"�߃ZD7@�`��p-���s	[�sM��[�ՓlwQу����Qh�ңI"z�I���K<��ܧˏг	70}�K��󚧗^��#x�%��L���������`A2�9��(��4�Y�<J�`꠱���\�;(�1wy��W��K2jZ�磗����1�����_�o ��ʡ����gظf ��4�&.����#�:T۝e�o-Ww!�U��p�y$����Ӡ�#���X�����^� rLmM"�ie������n��0/���Z��X�>�v��5��9�к�vr;�P�� ������m��'��*�?K�՜�+�+�}��bc��RU�pۦy�
yu6�02������iԫu��F4�m���[)�� e���h�J����
3���ӿ��YdҲ�s�t�y������_B����g��)Q�!}d	�(�9�ɺG�h3Ju:r����Շ�c��ל��X�:�L�IH9U�iB�  F"%�$Z�h�hG�ߎ��V�����Т��ۆg0[q;��mCsO|������b�TA�����<Ϳ���;mf�-�}V��&f�.�HS�¬a;h@�\NS��9�0Q;-��m�Jm��ډh�-�4vYM�j1�!}�ޏh(�0b�A�
�O�
'ur�%�,p_p�yh'{�ws����^�����G��4Be*��S2�~��"��U�mw���0�_"�ak���[�[�ľB+�܋�%9�9W�9g'�=A�|.�C��A�It�	+�84�P��0�5DNBI��T��,Kl���bJ�[^]����y8����ԙ����GE�O%(=��Y�E4���G�i�.���h�?�Gv��Gxd-d��;ُ�]v�+���z8O�J<s�P��tK�:Sq	��H���S,�Yyq�A��n����+󌇥L�-Ӝg�s]98�u�l�6gGR��*_�g�|�c��A�{�96�B�'�	�Ŭq4���(FU��6�;1.���^X@�5��K*NP�eЊ�|S>��ϵ�\��X��r�Ĩ��h�&M�y�D�E^8W�a�T�K�!i3g��.'W��'R!4��e|^z�:�*��V��J^�����e^�X�~E".!��ػ��A ��$_M����<{lMr��5��:P3��b��\Z#��h(,߸>�S�?��ض*�q�J�a⽢�_\�]��6�Rq��T�͡��-M�Km��aR���)[�S-T���Hu1�S!uPG����B�j�Q��cT�A���1�'�!Zt%_���6�-��͖'fېn�M|Y���-��&�e�Bc�Gy&*,�#<s?�Wt�|���E�~�	�u����N�B�Gߵ8���=ǝ�#�uu{h���|�o�+*7v��<'��x����~M���7��T�LA�u�������8IJt3��vosl�e����M�V���S����+i������4E}��kh��L���T}�V�-Ԫ��K�W,s�#4n�[����e� ��	1��:v2w����4���~�Z�p�tP�� ߹[$ݻͻus�4���ҼO7J�S7I�:��*ͣ�yD���1i>�����Sә���~T�}?�S�'Z� �z3{���"x��Ao7Bo7� �u��AcU��6���Ig�[��VZ�n���N!��.U��5j'mUߢ��.����{?t�
k����_'��\�}�'hj��U��ʏ�*���.<���0�ا{��z�O�}�*��uY@��aѽ��N$ʤ�d�ə����Ot���+����z���=��Q�n��.���ϰ�e!����h����H��p4V{)W�bu7U�{�R�ju����N����!?m��l��EC��(�s�l�<��6���4S��R���}��b�&� N��+�d7��/� �27{;�m�V�Ͽ:�o+��G�w����;��������̰���#�]GZ�Z�l@|�
��2K=����1�|ֆ�Y��cM��|�L@�H����^ ͱͱ�It���I�) z�_�b�l��3����r�K���I�sC���A����.��&���?H�O��g��ߤz�n� ��]4�w�@	{s�F]��`MC O�(BRu��~[�m�O�A#�(����g����r��4Q�@��K4W�L��+��רV�9�u���Z��՛Ԣޢ��mP����t��ݦ~O;Իt�z��Q`ky��b�|x��Q�ACY9b�����͍7׎�\��;Wǣ�}��$��3��w���e��<$*@��.;������s���0qd�R�}�/���""Q9� ���7��mp�'���ڕ:y��T���&諪��;�B'؟�X�?T:'����z�/w6+ ��L?�o|�g�Rrt�-����!������wQ�븛
�P��^�8@~�Or�OU�C���ٵU%���fԭp)W�[�%(Y��k�݇Z#Ou*OWv����4��L�!��x� u�n6��b��ׇg�3��+փ�����a<pKE�Y��<O�'f�-�Cc���x<K��M��xN�:�S�	傢�x��гq���� PK
    +Q�H��%`  �
  *  org/bridj/demangling/GCC4Demangler$1.class  �
      `      �UmWE~�l��i(4�JE[�P�@�R���J���FT�$CX�ٍ��*�7�����Zzʩ?�s���w6/	���̽��s_�;���W���öSJ����,�2�J�a��w��s��p�'T0�Bf�?�ɪg���n-��TMd�]2�9�L�eכ����bQX^�x,R��e8�v�
�!z ��҈�R��U���İ�SĦ
��Bg[��:�a����]�w}�Ak�b'���3zs{\�!U�����nًr�䞘qJ*�b8�"`�^�e�Vx�V��"����e���(�p�[��Дa�4�6v@|-�wqAG�c���"�#�a�i�Lb�+j�1���	�ލ�-�H��'�8�1��}��8�qU\��+��0[o9n%�-
^*~h@R$q-����@+U�݌�Îu�*���S)>�Թ���:�4��lG�-��5P�#y��ׯ��ON�;���v�����;4�-��sf0��S��)UD/ȥ���X~�M�ڄ����w�F�D��w6<����C����z����2���
��"�����1��shZFp��>=��3W����6�D�5R�`譫�/Ick���ib�!U�[�I����ߵ&���%jկ��f��T�'EThr��V����{�I�H5���*�sGΑ���a�$�+�;~�q�wc'N\��`K:Tz,�8��Y������f������M�*T��a��j9/��D�%�{U���]u
b��M�1/	o�&F-K8~Q��!�H���Y���h�C��$g��&�^�g&ƞ�Rb#����\`gs�x�5v1�}��/�ѣD�f�mN���m�S��Y��9�̿�gK�h|}9�,C���Y2���.�˭��6����>�p�`�S�dD��Z?�u�Ʊ(ީ2!�_��WZ}��w�	=P� �I������MZ)��(a�l���u���I��(n�!�ĿЕ��x�4��X���[�g6��G~�ʩ���	�w`h|�9j�v-��F�(��w�6#���c�+.y�+�"���
��\&��P�?�� v�w?�[�Fϟ��U�k�W�i�"���'J�7B:��Fp���>O�Az��PK
    +Q�H�/�e�  _3  (  org/bridj/demangling/GCC4Demangler.class  _3      �      �Z	|T�����$�	�@��b�I&!�� ,!H0$	Pqȼ$��83��U�K�Z�V��b���UDH@dq�j�.Ŷ�֥X[�vѶ�E�߽�͖&�+�7ｻ�{�Y������� ���Cᖲ�a�o]��h�[�`K�Y���-0_��"�v\�� 7e��u�^����0ՉLA�/1��g�5���YW�U0�������r�ى��"(�k����F�y�'	$5o_=�ub� C?
&�1�2��D���Y�����h[k����K�U0����U�����?t�$��4��?�D�j�c��֛��ǼZo�i�6�.*��[�����#ؤ4�{�K��=��v]������NL���(�=l4�7յ��Ѧ�h�-5*��:��@�o�L��ԖY�k����a�63i@�?�U�߈�Y���Hk�#�i��`�1�9j��i�R��3���Ԗ4�(���PҾ��{��6-}P���I��	�Z�9��G+���$Y�ި�Q�_��;g�^�h���l80��X�^�`�朞'�p��.�P.���"o���qb� ��NPK�fan�Sϙ{;#N��^��J�)���t^�v���Y���3�X��lTb!�Y��[
��ҋ�1�n��T)}v/��'��愥٨�27��].wc*���z�#��o'��f�Ȁ��x\�p�ζ�� a�����F0�6�6�h�^��8I-�b�Jø�1ʉ��H���&��K#�h��5X��7y��&�ػ�5��1����w�>U�Z���2AYu�Y�
�p8.�|1[�DÝ�T(�=�UԴ�A�Cia�@��d-J��T��-F���M1�V�{*�\����?� �j��6&e�#%���;�������T�7�b�g\�V����_"����_��(\Fi��ȉ;��3�gx̪�א2�W�Pؚ,\�ݣ�Ң��u�*��Nk�N\��kq=�>j�Kވ��j�s�M
f��i��#Ʋ�_9�gO᪢� �C���g-ʔQ\x"n�mJ���a
<;������>�S������ |w����\ޗ����V����V�bj�m���b˶�:�"]�t�U���k�4E�`������R8��~�<1^�&���6����&d��T�� ~���c�w�67��{8;>d��z5_#u���[��"�J
d�6E��=ܺ?����S�z�G�/{����LY�80n(]4l<��y��M�5Q5=b�i��Vr�Q�.V:+�U+��X���s*u������γd���/�E5�g��j�/gc,^���Go;�n�UIiZ��P�2����,�]ҷ��ʍ_�u��_�q�WO�a���V�.�3��ɂ7�Z�mz�I��ߙ�>*@~/�ޯ�z���̨
6�!�W�-������J-MM����"�m>�e�O,K�Nr!iaQ*y�R�_H��G�J�+���X)���Q�?9��t��*��df�������Xf$���NN��%.cr��l�d�c-��D�kɹό	*v;��'#KWD�F�]�B(�W��%C�)�Tk1����t�,��t0�C��\jUڵ\�����tP�x�$ D��:��2Xr� �23L�ܠ�Ou:H��2L��7xUʈl��HAUm��N��*��$����쉆�O��Ei8�[���jl�B�t�X/4>�'���e�h�`K�����p�)2Q�<ɍ��-eɢl�TrS�
�Mj�[JԸ�R�y}>��1���֗�Zgk�ԤSi���U�)<�d3Z�m�)��e�����S���{�n�٘ 3c���[���2��R߸��-sp�K*�gW�"H�U��"N�{���d�T*k/HQe~g�p�B����O�c�C���:��%�U���B�5!��&E��V뒥2ׅk����Q ��.��ѳ0��%+dn
�]� (8�\�4���i<�Ռچx*2Z��jI���Y15�T����}Z/�wZr�\�,����O�_���e�h�`���i�V�	U�[��Sd��Ē��3Qji��D�ؘ|��s�Z����
����Ɵ��''{�'�C���:�ӄ��͓��	_�v����m�h⫘��X
oAP�ʒ�C��1�-��1!i�t��	����$WӇxEi��}�J�
<�1kN����]҈ח�*��FG��</ة9�\���\Em)-��'b���>ݨ�b=���g$�����:�̷��ѦI�L�s��g�b�4C}��§A���Ԧ�U���V�*�s�~<�T�f6rM-���ؼSn�O��'$��[��|[}XD��$o'�I��ײ��3L�������|�,Q�+X�J�:�(���h�����խ)(l��#тP�(*)�O6&LZC
(w�/>߼@��N1���*�#\�qY�q�ܭoMh��x凚��v�`�%l-s"ZJB�,�ޔ����'�*bt�-�j����/�;�냡���w�Hz|���v��)��@I_N��L�Dv�0Ivr��$in�6�y��`iє�7+Ѥ�,yT�(�g��g�yL��~*��̽�FB���R��`���0��$$��f�5��i���I����Y�%?qKD��ԗm�7�~���k�����"V+��c�@b��o�{�4+�q
�_�WW|U�L"�]��^a�[^3w��j�A<R��_�o�:sH���0G�89�l���-o��oQ�Zc�[�1�ǈ�5�]��g��-ɻq��yu��ЗЅ�-�g�I^���}���3m�|�ᴱ�W��%�v�iGe�g�oq�&o`�7�W;��UT ��%�j�:���:��AE$��U_ޛ\U��#�������szV�b5�N[�(�?�L+r��&rmW�7�ʐ��`�ب�aD068 ^6�����o6xx��4�>�WYR��^L���n���z8a罼�Sҍ���l,�ƙ�1�ϳ�1�ў;�n����ݨasmc7�ٍ�b�n4<�����-0%aV��\4r5��
�9�>��L����r����E�9g�M}q�]kv+2���O�����-;�aT#U�S�u��.��t!�[��p�%������W�q�AJ�'iW׮W�kZ�
l�U���u̖+-}�y+��y��(���'(���R�[�\�=L+n܅�U�i�Y�lw"+���k)>*g�|�7*e�1����pS���q�Dk����@�9æN�����ʮsFmA6���pȒ�.l�e���]�+)݋mv�,݃�;Ԙ�՞���0{�	%*Lqqs��ݸ��HU~��I�b;~ą1�������؛��O�>�18��ka[+��9rfa}����<N�0o,v<��hϩi�-X�6T�;i�G��+�`���%c�������hͪ���0��1�=���ԍWw(!��s�a���s�ь�#x��ύ����o4͠75.��0�wgD��(�с؈��D=.I�ح���X�2��ɐ�J)�U/*�������!������S��3���Y��S�<�?y]�-�����v �,o[mՉ6��{N.ۋ�~e��������~?j^ieeX���u��y�'*�̶W��m�"��w��5:g͝x/�=������5�p
�z��O�搲P�g*�;6�e����୘�r������3��o�.���/�����[P���ToCn���6����F%7�t��Gӌ���nq�g�g>cMɌO!X�s�o�8��C=)1ݒ�����-��}�k,.)�+�,Ѿ�2�	h�L��;�3F�y��}���q�n��%��� G-X�����ţs�ަ�[{'�"W*��#��gI�ʓ.�l)b�j�����2��ڇ%��Z��p�Ӹ��[�L��	�%�2�L��2Ͼk�H%ώ=�%��e��s���Ǖ��U		��c~*П���Xq�u��Du�9I�$>���0�P`��6;�~��Bh�ä���r:���2�?��&'�SYG�ۊ�B�s��6K%�qv�2V�{��f���a��%$�|ډ�rg�BX�;�~��!��� �I32���3��U�>k+p�������׸���+���t|]F�:j}=�������o�B�(�&��[����*�6م��	l���ywP�m��9�o�{l#p�m�>r�?�.�5b�m=v�Bx�v)v۾�=��^�V�����Aj}ȶ�۞œ�7��<m�?�}����h���'�U�)��}
^���o��&-��<��ނw�p��`��hCbVY����1;�XxF3T� i�
�C�v"���v�^b���s���	VnvX>��z-�i1J�#�d��%�ʗ��\��W����|95ڗ6��8"_��bL��T�h��`�>`���.B>w2㨿��|L���B���OրO����^�
6��C�Ӵ��VG��[��ȰҲ�,���:��U���+3��1)�w��A����	 y�-�\fdjF��w*�x�<˓�e�X��`"���Xi����kl��v�~X�����J��L�'sl^��1qT��Kwē�<nr�JE'����:M�ùr-M��̑8�9�l�4�\GNc�W�z��4�K��98���OI�P�l���:Y�s�=�1@�F�Ŏ�@�db�da��P+H���:�E�ED��R�c�g���N&e���ǘ�O�Xfr�J�I9?�%\�t�LJ���u�M�/ 	(ޱC�rc����ڒ�X��-]r�Ut�c�����[�V��KS�{+��e�3�x�+Su��5<?SU.�/]f�ʌ� I�|�|j4�f�|�m��L2���v�<Nܫ# �����R�h<��q�UKaՒ�ES�I>� 郔b�L�����)8M��L9A���2���3��r�j&�7o��#�z��3^���m��2!Kv�ڬ)�be[={�{&Y�A���Q�Li�ʶ�L����:���ɦ��ڂ�s߫5�PѨ&�hKRi
��~��&��ҋA��M�z�Q�C�#�q8���{���.�����2��}_e���f{ȆR%<̉�bOB<0�:NƩ�S��&���(*t�C�2u���Yf�r{,0�dT�]W��b�m�Kk�4SF�%#�A]SJ��,�ƥX$�`�,'�ÅR�&i@XV�����e5��<���G�@FȅR ^/k���h��d.�G�4KDZY��r����<	���¬�2�����e�*M�Zl�N5_�;�k��4-޴7���3��;��uɁ�֜���)q����S�:��г�Y�K��Qx�!�L L=�?��}]����I����� �,a,i�xR��e��@
�	�\L����R\M�p��V҃;�r:d3��+���Sy�4,�Q�r�m�E�k�]�1�~�G��.y�ҷK~�ّ<f���ʜ����M�L�^W��c<꼺%7OC��K�xv�/�T�t꡾�FGN��1#gYCcf���_o��k.�4̛n���L=,��mT��#����1�=="q�r��ғz�:GŎN�/>c�z��}�=h>���y�S5�:��D+�y��T�)7��O�8y��.��;��x�JWn���<�{|ؐ�����xiN>zyE�4�s-Oai��P\e�G����t]$8�d���bD�5�9>>l}�I�R�,���K�$J%r#��MD���Xn!��6Z�Vt�m�Ln�����K�&F݃�e;�%uyI��+r?>����yH�&�p�-c�KN�n)�=R){�A����t�/7��&��nyV����������./ɻ�|,��\r$��[͐����	�?Gdg����@���ށ���>��y��}$�����}4e�����8���>��Sx��{����PK
    +Q�HA��D?  2  )  org/bridj/demangling/VC9Demangler$1.class  2      ?      �T�R�P�N��A���XZ ��`� �V�Q�*M�%ئ�$u��7pt�G/���u���_�{D�O�����$������K�|�@7��y'��+=��yΰ3Y��h�z���wZ�e0���9ㆡeI�M���%�����O��"=+�%-��_��y��
Y��CN&1@7Cd5~����d�^��a�֍##�P[0��w�p���Pm[�/��*Cl�4ela��o{��N�Jz=��l=r�����2��
��7k�-]�*�כJ�l�`h�n��mZ�VlC�N_T|o�.�f����o�Ѻ�h�S$���Ur�(��f-"d����b�볆3~�!���]Qъ
DBίu	��"��P�3(�ir���E鸰!~��q���Q}˟�$����4C}��Izq�q�A�{�fNf`&=:Q,�~��U������X���#�P�kNV�W��BM0HE��iN�̛Fv�p,#��S��P��l~��Kq�,i�ӌp���&"�I+c^�!��_��iZ�d��|�*a��l�%��ܛ�S��q�掞5\���K�`��h$"��~�>z�cIOҮ�,$Z�X�c���}I�魒i(J����D�Co�E>�	~Z�ޣe�5L�%�3��勋h{MH�1s<2�M���KHޠ�\�g�|�w��	��|�/�0��c�U8�>�4�}�ڱ2�я�3Rƻ$9N;��a�{!�vH��.=@��G�GHHO�KO1*=�(��ɧ�J��"C���C�4"��"�V�'�Fz����}/�!�.�T����^W�QS��C�]���PK
    +Q�H�sX"R  ,  B  org/bridj/demangling/VC9Demangler$AccessLevelAndStorageClass.class  ,      R      �QMK�@}kj���~�]<h�b-��Pzh���&Yӭi���˃�^�8I=x.��{3Û�ݷϗW g�g��*�\%�����PF��ίL����$��\�������<It0�ƔϹR�u�N�����?%N���?g�(3��P�ž��BfC�2q�J3�c�e2�d�C�+#������*�Jh�X�Y�Z&j��PJ'�{���t�/Zv����Jr7��1�m��l�
��1Fq�<q-sb�H�BH$8��J�IY�C��VDFF���M���L��fG{�Z�6)���梌MlQl�T�i��ݢs{E��QA�PK
    +Q�Ho�%b�    <  org/bridj/demangling/VC9Demangler$AnonymousTemplateArg.class        �      ��]kA�߳�d�tM��C[����loD��!R�
-��n����2�)��ԛ^XP/��(�l6$)],z1g�|�s�����O ����z�v���}5�=5p;�g�RO꽦
Շ EG28�E,�z`�KCq*\��ܷݡ��r�z&q��@���=J���+��P$�f�v�M��X�^�"����[�FX���ޅ~tJ��gbƚBṧ��a�v9�t��ӱ���2L��XF�7f|�q�����7���e�Nh��#��jd�3�j8�	���U��bMļB��M(�a*/��dii�¾LZ�=�w��DחG�!,�=%ߌ��ԓH�0�<��~���-_D��������A�8��W��v���0�.׿�z��7l��g`��z��&n�WB ��w�9�G�B	�9z�'̗|'Y�<����Ȕe`w�S��a�P�9�������D�����2�ip�}>���q��ߛ����(�
%��`�P�PK
    +Q�Hqn�A%  �  7  org/bridj/demangling/VC9Demangler$CVClassModifier.class  �      %      �OMK�@}�Ԧ�j?��G��P<���� �zPr�i�:%M`��y<��Q�lZA��Ûy�f�����;��	���p:S=Q�(�|�����f/��LY;(R~dm|�5V�*�D�&c=����sGNB������
!`+�*�4�u�=I\�g{��N	�3�yzN���V���&�:}bK8�����2�\��ʾ]�ϭ4��뛙3�`��bf���]Ѹ�smʅ�b�x����%���\�,t���+Z/�T�QJKmt7%j����*UK�
�V࣎�PK
    +Q�Hߙ�!�   �  4  org/bridj/demangling/VC9Demangler$DemanglingOp.class  �      �       �PMK�@�״ٶF��Cz�7?��*B޷�6�M�$��փ?�%n��R��aߛy3����\���)a���ύZ�|!_���#�2��� i.&[~�d ��<��M���t�0���M:�C����?*%���00����pU����
�2W�fh���1x�~������X���V�Z3i�F�0J�,-L(UbI�IkiƉ�2��@����cqע:衜��l:�����֞�jh��6��G�/PK
    +Q�H�G!  0G  '  org/bridj/demangling/VC9Demangler.class  0G      !      �{	|T���9�M2��$$@�a&1�l���0IX*�$If�̄E����n����H%QkݭK�Z���VZ�W��������f�ML��_?'��=��{���}��}��&�7�Ƅ#E�"��ӊ���PCS0�P����r��8��F�Hf�1��g}���iR���-/k�G��u���\*�i`�A��{_�<1���IL�}����%Jkk�he`C��4TWG�ŉ�L���3M���phss�5Zhni����'d����ޗ���L�~Z=y՛[K�N��^���2KLM;��c�����t#���*�������H���k��V�j���E�怓r��m��}+��Xep=��}�L�^f���-�Z-�q0<�H���C���ph��CyU��M�o��C�8�ǔ����r'��:��1��4I��z;��%��o�J��5^�e�ir/�$tަ�@�>�t��0����Z�M2$�)3y*e�)j���*���L��.C%�}󎙳19�$
�fC ��i�����@ep]��<S�߄�EU�֚9a�I�h��t�O�_��7K&�T�d�k�27ͥr��if	���5q�#{f�����٤a�:$��,C�ܝY��-�H4�S�lN���Y��p9�M��.X�jm�5�#��e&�DK�8u��ي�ؑ+LZF�30o0���`$e�ʤZ%1�q�`���5�ޤS�ةp�e�����P�_1��$9���F5G���%��["�089>�%�f'=�L��Q�<N���2����\)'2�m"J݃ub� �p��C�B��t���Cʙ)�.�G���������������zDb'�/k�R*Q�"�KH��V�{4xF@����6��sv���a��W��]��@ml��L:�Βӷ0���ӓ�h���a�ۃ�*ڡ�sS��4!���*,[���i8]��%XrTY����b�� �9b��~&p	��b�B�M�(&��1Qrz].9������]�IW�aAWC�!�a�HCTz���_�<eN�؞�m�n��Bƹ���j��jI$���`t��J%Q�@.L��:e�J�Jfl��)��S·�n�[��n���v_"���4��d�o��H�i���& j�M��-~wB%���`��ڠ��%�M�:�tݟA����]�N���
�ڔ�w����H�ډ��IQ���a�#�e��c�_�#r�]�?j�L��Ai7̥w'�Vsң�����*�ѣR�c8�	o������(��p��M��w���~2�~Km��z�nd�!��FBZ}vڸi�D�@L�Q�g�;�&l	�K�2���_D��4���d��[7�,����xK���UR�uѫ���--�P�r�2�!ևnG��-ވ�vQ����d�&�%y�SN~�O���r�wP_�w�{8h,�iL�@fŗ�C����S���n���p�$�"4H!�	�l�4��p�a�|XD��S����L�K<٩]�i2�-��c�N�^�n�4Q��|��/����i������=��Ťo��wH���í�d�/�D��O�Ql��M�����XkKS 7���(�u����.v�v�i�1c7�3�{����W��y]�GAt�O8r%-D���S����䁲V�6I%8��
��`7{8�%ں.�(��z0��&�a��o���^7����D�(5�Y<<s���)�%=NʥBVm=�Α�c`:<`��*��hU��J�V��{�9�I%9A����`0�%�*A�	���-ᐪ����YM��	p@�"v���J�U&p�����&-�Œ�;"�g$P��/J��d�#(��j-b�)<����4T�:w�,�ڧ��4�>���L�M��M.�m��g��%p�`���i��`�X7�ƋS��e(N1=ho�<_-�6|�I�h����wThRZ&W�FH�BLk
�b�&/�CK�h����@]n,�k~�����ST�����������޴h�-A��.ͣu$(!�Z�����f�S��ْv���nu�i���c���>Q�Ԗ%�}�p�<�i�T����1iu~�f��1it���Z�s#j�2~�lr�V�f�|:^7o��r��!��r�����O$AE]�6�,�n���UU���8!�k��!��o�
6�T&��%1xi�r	�UeV�[- ��O���{?I�F�����0��\��-�V�\����n��|a_ԥ�jGbN�Y_Bd �>�2�2,s��|�DQ�fd΢���x��R���0��r�5|����C����3x��N��q����Aof:j|�̭S�v|�J��(�ñ�u��fY#��q�v=�U�>ܭ)���C�g�R�K�W/._����!0Ԇ�8w�b��wAZ��!ZQo�=�]���н�	����m: �+3�^C;�Ҿ7�}7����Ã��A`�ʿ���r����b�+\����F�+ �s�`�A��.������ʠ#VW ��#�d@ҵk)����P�kd�E��1b^sKl����P�t��C�-kY�If3�������ð�w���O�o��k~Zf�C\u�r����t?"KF~�M�Y����F�_�;��C(�_Sf��ې"���K���
�ڏ������`�a�ZR]������-"[�jR#�}��܊@e݈�����!�f��=�Gת�i�{��y_޴�`|~E*�I6�GR�D諗�K]�GZkcaT�e����-$�����/�M>�������ޙ���ν�%�c^iTFy��G��aC-�j��L�Z����*-Է%��*��]�_��m޼�akQ�Ш`��`}=ra(f
VX��aX[����\d���X�M��n:NR�N�S#Ђ�O1�.�n��g�uakS,�Ҵ��5r����P-j2ŐGc��$��;Ć�R�,��4MB�Cuu����#lҙ�����Ѩ���P�FL1Zcsm˃�uS�ը#m(D�֦�)�Ҩq6�T�7���3q'c�J�4� Q4�_	�i�ܣ5�1�.>{���l��C��S4f�m�%~i ��h3�k��TI��5�&ӕ���b��m�S��9S��P���4��vB���k��-ƭ�rQ�IN����.���X��Gt��8�bM��}H�J�K5A��@+6N�L,�h���56��)�5��6m�q�S5����p�x�Ư��J�c�4�͹|~��D�k�cs�����z������zb��@�r=D3Dd[�-��tU����=E5��֐.{Pl�Bux���\y�� ���dƮ�M��,3�qB�8�_Ww�{�U��"�F@�0��Cj�yZ��Lq�ɿ��&[�U�O�X���E���F-�F@fx�yn����%.�=p/Y�P�1�en�!.G�D}�Cp�+�Q/����rѰː��*7�L���!�%�Ii���y�upn}
U�Z���Mq��Q
�x����)��e�@]C+{����4y#��1�+�L"o�b�q+���n7�Su#v T$(�W�ieH
0ػ�ŻW܃Ļ��5���P�V��jþO������/@8�L>��AXV�T���c(cGĿnZ�	P�ǿ��.Y���sA�h�unr��WԦs�� �ߣ�|{Q��J�Ě5�$��@�����+��-���h�={��.��/�y'Nd:�O>p8��&=G�K���݄-2d�G�/��p]@�U�!�xע�tXY�F�	���K���¢��Z������>�1-)�.�a�í�u]<�J�}�=��0�?���cݸ���3��*���J��P �ڬ@�Ɛ 1��f�g�$���06�fc�9��$���
:i�w/ͭ�y�h�Ò^<�������
"�t��V,�A��(���/� :{-���a�=�~���X~I�����W��\��
�ɂs-�Ă-�ۂ,xĂ�ւ�[�-�N�/m�l��|�z8_����6jM��i�F�SQ��yL��BX�'$^@:K��b�ϓ�
ԀE::���>CQ������kOHz���%i�zj���|��<�-!���Ms �R���1>�n���s4s4��?�?DK!�*���8�����oh5=O'�K��^���&��m������O)H�Q}A��5��[:��M��� �6��6q:���Y�Ep�%� ���������[-7Wz;���[����쥢_A�, �����\��It�EŎ,G�n�����f9:�,����d3E�i�&����bo7��:X���4��	;�˼�n&�xɒ���>Au#V�R^���z��B`/��˰���U)'�k{N��f�G�}��u<�Vcx�,���F�����8�r7�l#�'�س�WXh�|�u��	k�*9y;����_�ѝ������z8E*�h8���=q/�M?ν��g�Y�_�cR>	��%��q%�T�Q�^[��ov�l;U�-�s+E`i��� �h��F,�� ���^~��>�lx�8@��+��V�2��+�_��{�z����>^:�N��]�?r5��?选*��E�{iD��� ^��9�{ir���ۻ�N�{�z.QgI\��w���羚��^و��]��~��}��F��,��(������`N�Vp��62�&C��w�6s!40�Kq�d��N��2��p�P念h��C�yf�+��'�z�>���Hz��<_J/���@����2�-P�;-�K�j:٬�>�<s:xȬ�[6�?���45�v��qCR9r:x8|+��s|r,Ǳ��G��#���k��Y�X����*�aD�[Tx��l����4FF�.R8_!�A�����I�i\������FC��n���2��L ҟ�Ӳ����i�\p;��J�ђ,����	*vf9��m�/˹���шx �;{�CȰ�RS��"�: f��3�#�kq�7+�Ї�\��u�8�"�IwP?o&W!���%c�d�9��j^�Osx9� '�}���.M�DTȐjH�V�̳�F�C���U��r=��U��N�T^J����S�T��	4N��b��54����Ґ.����6"�;���ޣ	ଔ>�e�!r�'������)�����8�gt1��%0�+����������j��,�Mo�X�Gv1� ���f��4���"��܏��?����H�(���Z+k��5��+�fep������pR����e�@C���4a�R��%#R�6f��qڴ����Y2L���m4P���9#=����9;(�x�r�bG��4IR3�Sz'��Yr7e��̹�2��y<#=�u��������L�up��9R.����i��Y�}(������rz<�9��`�K�l>L��7���DB��7"������IG%�dѕ�*z3�?�V�|&�&qR�S	�"qe�:��)�s��G��b1�F��|>�N�q�s��^��}t�(lKBa-�@r8JJ�$[I0Se�lp���vN�xà��u�CꏗY�Z�#dj�I
���chO�a<�rxz����J�+���-�[<Mi*a��*\��Jwk�H�~��o6�V�0,�A�g�:����|i�o �N��z��:[�}��BW�٭���[�ςxa��-��a���|�UM;�h�N����ɗ�^���+m�K2�j�k�N���:Y��2_v���l��;�F�k�Wt�}��4I���EH_Jrٞ�=�&ݖݑ|�Ӷ��j�l���Ed��3[&p+����V����ۆ���ʱ*Q�!)�}�h�ujt��aZ������Nc�k�kh�]����R��[]���Aw�/� r�L]���JG��KSk��C
�����7���}MZ0ՂY�Rp$W��F���72��C�_ryD�E._��"�a��p�n�o+����7w��(U�rJ�hw�n��:�/���2^�����5t�� ����7��)�h@xX�t�x@4���* ���	Ua{�f�YP��{����\��n	e�,��sȃq��J^ Ύ�>��\�x1��K�B��k�ɯG��+�n�ᇐ�w��8�)�8���!���~~���c��������A����C�U��M��g��|���g�
>O,���b�*V�Eb_,|���W���Zq_'����^�A<�7�]|���7����2l��M|·�����)~��m���7f�/�Y�Kc?l�����X���c,�G������'����76� ����
�AoyS0��4b`�$�������5z���_JA���ZBJ�%z�F��,�&~���4���L~A_�D+y������c{���{�m�$�=�;�E�<���C�c�!��(�grկa�L�Od�|~�/�Y�M��&�3�{#�+�.Z4�o��o�xނ������ˠ�G��k�
��3Sˏ��k�~��������U����*S�iTq��I&E��C��(�i����?����x��H��{�V��JҥO���f�;�B�vvY��Aͤ*fG�bnC5�@AV�����=�ce[���m4�z�OC�e�x-�%wZa��N�n�Ғ�3[s�(�P����J[���Q�OP];�lDY]�%�MS���Q��3(� ��o��/��/i(�}CH�k�;Z/���]t:髄;��z/�Tc ��&��dJ�rQj�+��o�| @���Z߅}�J�9��^_"�4:Ա�q����x8 �+Ӵ49@��1�lR�:"!��;g�*K ��Y	8����v'�����/_�	�_���w
�t@�dF� � �^@!`"��4����q���y��'NjOʘvX2^�JP��;˳H�Yn�p9�j��(zN_�f��֝�{� ��X����&@��|�}"~7��T��m�MQ����Co���B�a�1�>#�ȡ/�(�J�ҷb,}/��8v�|v!{�� }��<DL��b2�)�+�q������D	O�y
2�1�KD9��\�;�+E%/��Z,�b)�,�y�X�ub%��,�8�?���b-*��AQ�_�z�J4��4�^4�Y	�h.�!�.���V���+��ꭐ]iż��Z`��<5�dU���|9�U;��7�C�%��Um���Jo��M_�q.BFۏ/*:�j6rd�m����@US4�Xq�Ļm:U��q"Z��Q�B���,:B�M��9T"Υ9�<*Љb+-R���j�%�F\Ju�n���JȣX�<�a�5�NqA��p?m��=6kIW�sM�����i��u�A��$=��V������?��>����N�Ҍ�饝�}>4��
��{�*	)�KF��o�p
@���np�=�Se�{)G<@G�����pJ�v�R�8���G!ydR��W�+^��֛�t�Ȱ��Q>%� TBF}9Ht�`��F�G���s,ɜ��gd˥U��A�[���[ȓ�SV��Z]�b0;���p1#��U�r2��Q�>A��ƈ��N�H���,Dj~��(�z��Ou�Z��mq��}a�OuIq�y;�-q�8�J./��(�z�s�@9�Ku�S)C�*nSG�M�}�J�v�X�R�>,zs�(�9���c��d�mSP�L������-o�_������?��UKI�C �������%k$U�xJwȫ7q�
��m*��-�T�� �Kݲ&>_�3���B�](ޣQ�}�T >�S1Z��ħ)�{�j�P>���GI"1�G�3�"��H�����7!ͪ�k~%a�DM�(��P�=�(�)~���fɇ{�0E><��|�%�ʇ��e�0~���G��C�� ��Z�\��t���]��l���u�
B�s>�J�%��?h��
*��V�oi5��Sſh��7b�ԀE��@UjP��F�Im6�t�a��?�k����.6�UƐ�*tk]A_��{�{�Y�)�(��2�ҍ��<ς	�@o̲��R���c�O�nA�'��S��x7�����}�n�~�s�����3v��6:�6�P#Mj$Y
M�LN~wm�x	r��ڨD�Z��`$O���G�&Yv��k�G�c�hZ���W0,Y���#���	E��<�h#������������L�y�x&(���hr�4�ȣ��x�n��1
��1���=�8�G�y�q"��<Ml���'���6��ƨ操�GC[o�p�X�c-oDs{����1�ը�K��^n�c=�j4�SF��1Z�E�t~ٰ�0�SVd*"V�#���y:A0%O#��"������ꨃ�+K�[�Kw��Ȭ.�{��2��ѹ8h�#��,ʠl����7�z�@�s�������Ǹ�
��Ex�����=�S�;�3�{,��PK
    +Q�H�˲T�   �   /  org/bridj/dyncall/DyncallLibrary$DCCallVM.class  �       �       ;�o�>CnF���t���̔,��ʼ�Ĝ}퓙T�XT�������3022d%�%��$���'e�&��3032�j�)bdP d4;#�|F���Ң�T�̜TFϼ��"�����b�:&`b���\@��$�����	 PK
    +Q�H"���   �   /  org/bridj/dyncall/DyncallLibrary$DCstruct.class  �       �       ;�o�>CnF���t���̔,��ʼ�Ĝ}퓙T�XT���\\RT�\����� ��X��������
efdFբR�Ƞ@�hv6F���\���Eɩn�9��<�yy�E�9��ũ�@uL,���	&Y��4H����� PK
    +Q�H�^�H7  �  &  org/bridj/dyncall/DyncallLibrary.class  �      7      ����f�5is4i��W�]�t�lm)�
�d'2�e{�8�b���#Y��8l�l܌��a�kc��a+Ǹ�͟<��J�_���q?G��y������蕬���}��5�	�:����k����g��h�+�Y+��I��k�ic�aث���5�����aϫ������a��uA�ͧ�F��#5vz[�g���C����s�K�
E��*�!�*�p@�E6=�Ef��F2©+rUW���D�����<��wB�I��	M��U%�N�5bT���pc� <P��ǈi�5���
��K�+jS��՜3hH��b���˅B�XJ)�l^I��IpI;2�ijAW�j%QL�t��i��ؑ�U�E��2�e������b�~R�$�Ө0&L%�\����դ��s,>X.���S�؇�3KRȣb�H,����U�&4u)�M�J,a�tB/Q٥\Y�	�XF%���:�S9\�%b��W�*���p���/9/���i��<@l�%�&��#[\�e�45W���`8;%_Nj)b��:�,���!b
u�^He��	���WZ.g���[Ã�bY����L;zW��l"��kCLH�3\��Gbl�j�n����-����O�L|�4�����NwLP��Z��2/X��.�'���YV����-�15��/��z����I0�/�\>��&+��P�l3�}i�@8��ok�\p�
�TZ��W�Jk���c=6��v�baŉySG�H	%���򲒒i�H]v(Z=Z,�"�m�ʗi�AO1��ӱ��Sd?%��E˶����U��%��Q��I0蝴���i绡��jk��3onA�f3sBT��l�t�m:r,x��z-�&�����H0T�ͦ�Q߬SG��q�*q���j�q�w���v�H��Q꥟t\���N܆��j{���ث]2$`gd�2	�	��h���O7���i"���)Nk��m�7F��S�@��e����@��cd�=���Oy�c�:c�,�U��*�s�*d��90I�I�����H���=��޵�Ȃ�|��Y*MkM"���9T�]HBy�,�{i���������M��K��r]��S��Fd�{6�Ƨ��gNi�l`��n'jƿ(��J��a�dIN�|ǂQt릮�6�d��hX���i�X�+R�3�y²���X���/��&?Ѷ'�of��v�\���;�!����8ٱ��a{�SfP������_1\���+��&4L,�Z_1]�̈�1���������y�+�'��Q��>��Q�jZ8D�p�uu��x�Y�d����Q�hucd�#�o�Lfcd�#Cou�/Z&&~?낻���K<�=���̈́/��5з5Q���죶�G�L��}�����/����ݧ�w�m��D%{]�SȣKR��&�5�癋�w.xy����U���~��<����(�0�;-�f�-�3�ڶ����4�p9l��� G`&a
$�>yQ ��;`'�]Ȼރ<#�%H�F�	���
�8�_��O��#_!���(�G�$�g���~�+#�?92��|��W#_#��B~���i���終�:�����t�~�?9!pY��`O#/	���
��g	v2�&p9'p� �?�(��\�����G>&�G�!��s~.��"�z��U�D���W�kבM�O �
|��֐_(py]��~
�E��M�=��F�_�|F�	�]"������A<J���{��g����Pvn�W��G��?Z [oP�F���*����p����� 4�
�����c��D���:�?A~}�� �q�)���F�?C~S����'�Mfd�ߗ7�tނ���!���8����ο@~'���/��ws�_���[p���j�7��>x?��  >�����s��G"�����c�y|m���ȟ�Or�=��Ӝ����,�?">ϵ�������g��E��/�o����4�K�e����q��SO�9�_���p�\��{����I�^�����H�9{�y�_�o�7�ퟡT��~~��'8x/|�,ͺ}�\�S]�Ͽ��f�7���~Ʒ����h���D���#�KF�PK
    +Q�H�b;��   �     org/bridj/func/Fun0.class  �       �       ;�o�>CF���t���̔,��Ҽd}��<vFF�+��ĲD��ļt}�����k;L!Ft1vFN�Qz )F�Ă��JFMlpg��%����jh�� Ÿ��K��S�2sR��X@�h0;P�����37�f PK
    +Q�H#e�\�   	    org/bridj/func/Fun1.class  	      �       ;�o�>CF���t���̔,��Ҽd}��<CvFF[�+��ĲD��ļt}�����kGC,�v�B��b�,�� ��@R���9��j��5������XRZ�
dk�8Zk�� Ź��K��S�2sR��X@�h;P-�����37�f PK
    +Q�H�2G�   4    org/bridj/func/Fun2.class  4      �       ;�o�>CF���t���̔,��Ҽd}��<#vFF� �+��ĲD��ļt}�����kGCl�FX�0����X8A�ꁤX
r*,40�c�hb��383=/���(���W#���:���Z3$(��_Z��ꖙ�������� �@G�3p0 �yL\@a13p�i6 PK
    +Q�H�s6    5  org/bridj/jawt/JAWT$FreeDrawingSurface_callback.class        6      �PMK�@}Ӧ����*x<�=��RP�-�X6�Z7�l��wy<��Q�$�Pf��}og����@72s�3j��X&�����x`�<7b��|��[�˩/���}D�}��_|�`g��@,��¸�2��wB���Jz�b�5q`�Z��u��ܩ���s�{*���%�������N��&lޏfܯ#�M�Q��8K�����*}��d쑚k�����
�������򋫣(5���׹�Z�~(�X��
��l@�Gp���H���'8�y���� ��M�:G9g���m�w�{��*a�1�-��5�~PK
    +Q�H� ;�`  �  /  org/bridj/jawt/JAWT$GetComponent_callback.class  �      `      �PMK1}S�]�֯���A��*X<�dQQ�-�(�kjM$���)O��?J����+�����7�yy}z��5B��n%��W�ۨr�{�*��7�7FK�uD��Ε"���O~���u�=1�B������KX�Y���+�]���pO]x���\L2�jJ��N�(�s��tfNt�B�V�ߟ����Cs%	Սou'F�H�jUNืo�Y$�0��V��/[�#L7��ǃ�@��k����2�H�[���_;����m֓�iB�i�#�U<A�Pki��C:�H�
��e?Ϸ
G��|����y�}�D��l�s��Pd�4�]f[�4V9���b��e�IxoPK
    +Q�H�f�m  �  4  org/bridj/jawt/JAWT$GetDrawingSurface_callback.class  �      m      �P�NA���u_�F=�p@�g��G$��@�Hfa�A�M��'�9�L<�~���/���LwMMwMO��=� 8�!�n�5����ĝ��]62g�?6�N�n}h�D[�ڢ�wE��R�=�/>Jp��\O�a9D�F���.N���š�\#�}�R;?�#kL/�1K��2(*��!��k&1��,,,�Z��}���J��I(d4_xJ��B���({IU=�n
��ۗ� �J���֕�qꪫ�?4�B�-N�c¸B)d��~)l�I9�����#$��д�
�L�k-M�/9�va���s\�S�3q��?a�q|��1�A"�e���c�cV��xs\��5F1lsN1��ƌ� �*sp�PK
    +Q�H
|�#L  E  '  org/bridj/jawt/JAWT$Lock_callback.class  E      L      �PMO�@}�ZѢ��"�`㹄�M 1���lK��5ۂ�gy2���G���0n2��μ}��o�/� �p�P�ذ�M�	������f����gsg��1�߲�W=͠���	�s��
+Y��/�wR��-�|�u{��Bc��-S�ΐ]h�4�/�C��汁b
6��V��ֿC��"�y0u����@��+�Ɛ�����:��ސK�m�ĉ�h	����lW~V���<�I��
��ҫ���l%����L:m��we��a�J)5^)�xr�e���0s򌭧��K9�(BG�p�"�T��m��O����epH�KAŚ�!G.hPK
    +Q�H�{�EO  K  )  org/bridj/jawt/JAWT$Unlock_callback.class  K      O      �P�JA=��ۚeiYY=D�CK�+BH�"h��:��6�j�Y==�}Ttw�
5h`�9s�g������s2�z`�Z����?v��S�Q�����繼72��?��w>�`�gC>��%f&��9G��y)��t5�O�F�~��&,���2�ə�HE*T�r7�udR0��`�r�p��Ǡ�H5�G�!_��q�K픻dX��T�6}j�r-��NhΦT�5yp���Xm9P<�h����»>©F����D�ĕm�u���y|<c�16\1�pv�y:ل�0q���稼C1=K"��.�d��[�&�i��#��a�X&V)rY��	PK
    +Q�H�\�"Z  L	    org/bridj/jawt/JAWT.class  L	      Z      ��moE��;�ڹ�>�iKCC��}�@ҤI����i�	��%������T��H�(
R_���=��|g�,�����vvg�����; ��L��U[���_ݗ���������cE3��p���ڡ��@�X-��C)p�ql(��6�V ��5��C�u�@ހ.'�>T:t}M����f��S4���n]z�@9%��u���_}M��۴k��K���T���4�3���}�)��Ħ�\�k�����I�j��Z��j _�z��~�m�9/0;�@`!�-2����l���ተ0+p)���U�=2�Xt�.	�J��1WD� �n�yi��n}��a��s����*o��cC`���5���l�lT�Yc�\`zPoaA`rO��#���� �W�5��ظ��ETq��/9��';�ī�DǼɗ�o�_	^��@^x�R�IO}W�*�.��b��V|�+�pl|�%�C��`��cƘ/S�f�֟���Y����2{㴮��|�N�ۑ�+[��6n�Z=��T��luY9j���X���)%H���ivڭ���bZ�Tm���4��"ԃ�Q'�����Ή�O���=���/��~7h�5פ�v�VAݓ���`���7=�Sl36/G�����d��n�a
�9ڽM�����/R�'�7�n�S��r�m��'���p����G��v���8�y��A9Bދ��<�f���G����=�BOC��&���q��iG<@��F�?�������͓$z�b%=>z+Fo&я(�艑��c��$z���5���c�F���>5Z��$z��f��6�:���|R��<Ky��T�E��˔Wp-�DH�3GY6D�LØ�PK
    +Q�H	{]�  �     org/bridj/jawt/JAWTUtils$1.class  �      �      uRMo�@}��qBk�BK)�B��T­ĭ	E �B����6�*��]W�M8 �OH $� ~bքri���f������'�<"�ef�J��X|�a����Ъ4��� B0S�B�·ñ���2a{n� ��d���/2-�}7�ZS�c��x	{�V��Q%�F��	��r_J�J�$�����kv7����9�T�#-�t*O�V�a�{m5���Jh�]X���M�gOUNX��]�2͒�����_LX�
ś.X)�����f�d="=F9�,��{��4�L�}61�|����Y��荴�YBh��Z�~*�\��f��	@A�t�g(�	p����{±��{[���}ǭ/��w�1\�
V�n���|���lB�<���W������m�]~��;X/&Tq��Q�w�?��g�?(�}<d��:�5g,]g���+�?PK
    +Q�Hwq@��   
  6  org/bridj/jawt/JAWTUtils$LockedComponentRunnable.class  
      �       u���@��UZ�;���am%	�H����DZ5#Ӗw�� Jt,��Ž'��9��~<��$��>�@�Q�~��rz���8�z+�E4S���B�BJ���	�q�ryb� a��"�~�����؄Ο��Y���o�q���rp x[U�P�cC�)���<�DV�VP��\x�����5���`u�� PK
    +Q�H����      org/bridj/jawt/JAWTUtils.class        �      �W�[������0x,Y8*�T"�*	�]�	�!���� ��fv�6��i��>��Wl�mmc ���Jڴ�����y���>��3�r�`H�a������z����g��������^�L6�nSG���Ά!������n�7��;h$�0��6�{���cR���CF���ؖa���X�ޛ6�(X>ϥ��y�m#"�z�=?	��ѝu��ca���F�B���h�wt����V׈ӧ'����;�n��G�z:ݫ'��X"���ل��>/�M�
�!|�@e M���	�#7�r��VT�	4/��A+=�O���9@�� ��8�1����� 0��L�tw���X�:!��f��I̗m["��;�%�����G��i$��h�d��*6b��h��_��
T4��@* �_��B�HKn�
W�:zf�Lf�m:�5�B�v���3�T��f=��W�lQpZ�<����I#㚶�6`��Y�k3��a8Yʹ���6l��Me�Ǘ����u����w)؎V�XW���#�gK����b7�H��K�ئ�N��˝6��`�����f�-�N�oDBA��{���"Q@ Iލ
�)z�����1Ç]��L)͵5*�I�Z�礭.�A�hehx)pson/����Gj|?��^k���28�N(�*�
�H��4��`�FMw�o�8�������d��D������r
��U�ل�?���_�C�٧}ߞN�z�����4#��l�3���b�خ6��`f��$�`Hƙ�w��LZ?!�Ta��3��Zj��j�cx�R����BX�ڛ�{�t�6n��SpU��͊ٵ��%�%Lu'd��d�3�c�Q�.���oSP���tv��3�oK���<t��,�3�7����#f:%��<&_�M��e=�|C��o�����Z�I��LưR^)lo����.�[
z�ʼ��G�>I�~�2��/����|ć$�YɲT|T���
�@}�t�'��'V�\ ���}��9=p�Q�/�@<P�<������,c��c����T���g;þ�R����u�'�n�3ہ/��9#���C����J9��*���$*������vH�~EA-���R8����_�V�Z�%{�[`[}m�ׄK2&�������� ����`��!:��>�On$�瘒AfL��h���[6�W^D��e�-h��׳5���R��tL/�8@g�ӭ��jy`f��Q���=�أ�??UQ�E���[q�����ɍ��R��eI���o8+gX�n��hw;^z�NN�/��2��Pt����i�*��ь�JO��C�cJx���	�2:G�{'���v"3��t�#N��cʃ�nY��u`#�D/�p-J8�q����<��UHh�8�_��W���	q�矴h&�=�H'��ͱ-���3���q�S<
���cs	�����6��gQ1��=�;Ǳ��$�{���5�}��	t�o�0�{�I���q��aG�C��P�)����&��kV���5X����J�#g��	��ղ� [�a�p��b�I�mԘ�5.z�&.�I͔nz*�D��aIu<�d=�F[B�c8�)Z����h�m)����Zi�$���>>������i\��#�l)������a���=�,z��l�O͡&ͧ�K���X�G�T�%�<5�>)/y�.y�b�S�p���ʟ��$����ZI�͋�n���U\��cd���_��Es`�E׮�s��/�B_���z�)�E�Y#V�5Ǔ��%�b�1+��p�ˌ�������Y����kxNFP4�"/w~�����LWPB\(�!�����y�J`����J���_��y��y�W)��q5��R�Ld^	j�����+�0��Y8��y����Q����Q�a�gv]b~M��M}�6@I&m����?L_�E9l���f��x��������	j.Ko�~.���CW�;74LB��8�_O���.'�?D.{�X��x)W���g�?>���P�(����Q��r��S�����A2��;I�S��y�&���G��^3)�=�NR�y*+�Г��^Ī��g��!$�W#�u%�7r�床�j�ׄ"�PK
    +Q�H��g=  d  H  org/bridj/jawt/JAWT_DrawingSurface$FreeDrawingSurfaceInfo_callback.class  d      =      �P]KA=���m_V�[=X-=+R)�!(�(��h�������)�Џ��n�܏9w�{�����3�.�;��É3��й�����ϥw#3�8j!~Cm5����˽i�����������>��˥s�2�/�g�֤�a�!]9��ȣP��U+��C���)�$#�LOC���FK
S=�^C�^�h���Fr���1lt��ѽ+�'��ʱ�ad(?_@Y�C�q��z"^���x�%cn���0����h!�I���!�E7�"��9y�������kX��M�M����&�;��]�R�e�G1�M!�+�PK
    +Q�HP�O�D  �  G  org/bridj/jawt/JAWT_DrawingSurface$GetDrawingSurfaceInfo_callback.class  �      D      �P[KA�FWM�nv�)(zPZzV�(�@�G�]G�favW�[==��Q��-��RB�|g�������3�STھ�X����5�кl��g�/���"=�8��O�������pwV c(�؟|����w2�s�p�w����g�7��a�![�LQ*��*��ʀ���{�U�j��C��M�ڗ*�QK��QF��Ѐk�O�cǰѕJ\Ew��L�''�����>�Hs�9��V�Ɍ�l�RϏ�+�eܓ�QJh��A ��l|2`��o��"d���#̇�L�|'��u�m�|����$w���(�}�X6�V��PK
    +Q�H�=��5  *  6  org/bridj/jawt/JAWT_DrawingSurface$Lock_callback.class  *      5      �P]KA=WWM[��2_����zU�0C"P�Qf��F�Y�����S�C?��ݢ����ιsΝ;/�O� NP#f�F���T,"���f0:7b����[�Ƀ^��F��}Wx��P�Ru>�,��D~4sA���QyB�G7B����ڄl�1�QD��+�S!���	�l��<�IB��M~(I�ltٽ��^a����(��r��zOiy߻�|0ž�hņ�����l��K� 6��P����Z��/�P��2<z�2��'8n��a$���#쇴\�h��(c�q�w>e��#`������j��˘�fP��U|PK
    +Q�HC�^7  0  8  org/bridj/jawt/JAWT_DrawingSurface$Unlock_callback.class  0      7      �PMK�@}ۦ���+j�U��zhP��$"(E��z,�t���]�$���$x����I)�3o��Λ�}y}zp�Ñ6c�7r4q'|�'7���s�ƽ���@�_�P�a��������|�y�|���@�9�3ΰ�{��k?�1�RɸÐ�76ʨT`a����d�p���-��j����Z�&p����i5���坮��7���觎��J%.�{_��ܓc���P�^ ��Ø�Nָ�Ӊ	ęLu�s���BE"�v���ӓK����\BFX8x������;��n�3fn�
X�x+{�MV͢vS�JX��oPK
    +Q�Ha Z��  t  (  org/bridj/jawt/JAWT_DrawingSurface.class  t      �      ��kOA�ߡ-KKE�* V-U)WoE�5��E4C��P��d�-�_ib4�?�e<�4�.�l����s�9�s����� �C�aʲ�ɂ-K��}~�$_�}��ݰ��T�|���Ea�1����Zt�
���0�4Y4��k�a8w��+��ɂ���C��ͪ`�c����jB9�R;���;Ǧ�#���4�;Q�2���n�x��@���cdX�A��B4��j�:C�c��İ�#�+�M��0�>�a�G�\��2\�5��x�j��hc`���2t/K%��@|z'��� �	�
竬0�r�7L�Uc�O�	kI�������Ha�R�`��@���٭T�������Sϔ�SO�Rf��X'7%�m��(b&�H�a8�&��]��>t��E_д��I�o�ywio��']�g!���{?����m����}KN*�Y=,�n}W���Y�dXS�r��!U&��eŝ�Mq�f��t���Z�b}�0�}����w��.�ͅ�?�K�䭪]�+�*%��+Q�-jʠn_ЯY_S4[ e�Љ_���[�4FO��l��9=� K9"�m�h������$�����D�P�]�*Vh��;�Y�%�k��Bf��y�B� C���x�Ɯ��"�Rt�/t��^��<n�6|�?���^���-�=��_����`�+���	�K4��
�U�k��C�ä�����.J�t
���������PK
    +Q�H��t�H  #  ,  org/bridj/jawt/JAWT_DrawingSurfaceInfo.class  #      H      ���oAƿ�-,^ji�R/P�Z/4&��d͆���'cp�2�,�4�7������g�(�@�K�<�ٙ�~�;g��o���1Ú��uO6;�?��/�^�}��C�ڵ�k�T�5���gk�4��zG4|Q��a����a�k�Re[�=0���	CL�gHlJ%���|a��<�IĐ�}���1����<p��r���g��Ǵ�\�|�ѱL�ڶN���!"I�h��v*&.`qd&�,3�m�h@e(�'X�&V��ܙX��$.�2Yi��)��D�T������q;v	�U��2"T�r_��0����ln�+��u�Жn2������\Ñ5�An��~赤ȏ���Ȟb�2qwu�{�4L#b4�6	�`���sO�#��@}��ՠ[�hee7P��}ٓ�����SU��.&kn�5Ķtrt�1}�H����q����x�+�Ϻ�x@�9\Dg(n�d�=2�stJ�":XM�`�=B�S��� l�
H��<}��
�S����/��+����d�L��#����ajz�ZSs�(�h4q�����#��S��}��'���,�wK5z��PK
    +Q�HY�h�  �  #  org/bridj/jawt/JAWT_Rectangle.class  �      �      ��[k�@��g�ll6Z�ެ��z��A_"b�`�-�G������NZ��|D�?�J<I�b��}�s��~����� ��C���a��j0����v��>Ⱦz�JDX�L94y�7�ɘ\X���ũ �ŗ%B� VI.��������lFh�TZ�W���� σ���HM[��c }��#�J�鞒� �xQ*#,��M�������
�=w�Fh����������"a��X�-7q�g;/���350��h��#��#SZ|@�M6�{��/ҞȕHRyT
�b��|_�$2��Y?(�Q'��&��ZgF�i��w�y_�Tb��������|V���
XS��~����X�N\�5��5+�3����Ye�sX���~�j����O5�7Ex�G,[���ύ�f�9iυ��;��f �����Ȼ��g �s!�֑���qU�����W~PK
    +Q�H�gh�8    '  org/bridj/jawt/JawtLibrary$JNIEnv.class        8      ��[KA�����fy++_B����_��e� �z�u��ݘ]?VOB}�>Ttv�2�2g���;g��_^��J�����h厚#�6-6�r�гC��=���P�j���{�+/��@�PXќ��T��Sd���3婰MHխ�AY�&RX�Dx���-�!\Wˀ���e�+�妭��K��<�㻒P����V��~dy[y�7yp�^f�+���BEA��yRw�"d�<':	P�)�����d�s��z�m�_�b��*�<
��aߌk}�q�����B�8���7k��Y���ƚ4��
�o`�PK
    +Q�H��K  E     org/bridj/jawt/JawtLibrary.class  E      K      }T�NA=C��R("EQ�ʊ�� A�R�u�b5񥙖M���&�[�_�O� ?�x�T�	`��;�Ι3�޹�_������߲�:m[m�)��4�j�����j�siu�nY�F�m�q���6C`�(I�����ȹ�t]�as�eb��Cu�8ٱ���S\)�
y}Ǹ���Z`��{\w��ۺ�����\�0�/ 
1�=d�7�Z�R-�K�������������@�zR9�����FpL = �+�rńټ�Ax�|RگF����U��;ֲ�nc1�a�a.�G,:ח�ƌ��ݐN �ayJ���}E(�A`l���_�0�h�q�p�w[* ;�G&��X��=�R���{��)ݴ�5e�&}%���:J���Y����DU���>��������3o�^Q��s����d���M�@�R�]��� p��L�j*PL0���P�D,c�� �"�I�9Y37�"����7#x��V��E�<q&�`拯N�����Y���_{�Ǵ�� �p��	�I� /��;�`���x��o`�	������w�I�����]�W��5��;>�g=yv�h	~$�����TO�E�?PK
    +Q�H����7�  �� -  org/bridj/lib/darwin_universal/libbridj.dylib  ��     7�      �}y|E�xO��E�\A�QI\� ��h��h���rIf�hb22M3�UTTt#�kvE�(� &�E��%J���!r�ｪ��N���������|z���ޫ���uu�<}�|[��Dr�..k��r�����8a���1\�o���pr�p�g�&���Cٌ�j:���B�QZ�Q\��q\�gRn��JN��Yͳ�R+��F�o�Ԭi��f��[�;�7YB�-җ�랝3cJ3��<E�;/=k���&�3'=�9az�{ꌌ�Ya�fv����[��9-#7�a���@�{�p�|��y|�3g�5�z|c(�8ͳ������x"g��	93�g��+c��#����˚:!{66�)}�X
�tO�9�|(g%Q�'�6ƦIP�+����^��5y��Z:���j�[�k)3ݺg=�X�/Q�Ň�u�~ZƄܹ�'͜6a�{v��/�z��C~����_qE��yn����bZN�ۈ���j���}`�r�gL�®g�Wk���FY0�Oaڈ���K���[n_*��Sfge��Ϥ�&j�/���_~��_|������Z6��3��]����l�/_����/��٦���յ�O%����k�[Ɨ9s���3��W2��k�t:->�D=%<N��w���Λ�rN�?���>�5�����8C����Y�s�̜�����)9Ifd�sϚ�3)w�#�g����9Y���Ι|��ٙ�g��0;+w�gv&$̜=e�$H|3��1�?� @3;7cF��@]�L��i��X���a�r7��WH�� ���k`�^󢅻��@�׍��.añ/W�4��9e�q�~H�XG��ۮ=��),/�f���55��;�p�蹹��7Wx�_G�
p�Y�������M�3g?�;������rfθ![�p/T���Ig��tq\��F��d��ސ�%��M������E��F̜��2m6CS�qF�Pbo����f���k��m��g����������������6���qͱ`�6:ط��������@1��ğl���w8�o�IA<#HC��	oq��p~�8Ν1��k����鑆:$w�8���C��<���'dpn�S�o�H�'r��i�U�8����`A��v����o��=l�0>0;qͳ
�AW��qj��v���m�#j
{����J�8����Q��Rr�|�t������$��/ /π2����D[���j���
��ոӄ��(S~�=Gb�ª���-�GqA*p���O�^JCΤ���)�R���_������\|>��X�����I�sN��`�A�"x��㔘�|�A�Q�%P"d���o�
�Z�ƓZ���Jm��I��6iOV�_�:L�ۭXjP�q/k�櫁��X?(|�4�S<&�yK�}���2�F'p��o��	��gX{��Ǥ�*���z��۫����J����v�^�_��ky�m/�X�w:�]�w�d6�'�:m�䯠.��8{�6R��h�:�rC妁��_(<��ı���ٯ�������
L�5��z��-�V(y<��-5�=�m5�;d���5b!��+R^���֮��U����F���:~7����r���H�����
��� �j�Z���j���?:]��C܍l�M�y]r��,?����)�l�k��������2�)�N�쮈k�4���6����Y���!��l-t���X�g�%��ߒ]�>N�^-����x�!Ӥ�N)7�!�&����_��y ��ڽG��l��Fy�����;��[��F���QX�=�.�k}�Cze}
�('}S���xit:6Dy��~�%�tH�$�U�nsO2G?$H����)wOp�ہT
y�cەC'$OM�����g��P��V;����
t�%�V�*+�z<��Ւry$f :����������Zi��bf��}��+I����׿v��<ΠWfDiz�m{�z��^����N��^q�r4��_߹�3�rP�oa�����oTo%'��
0�4&!U�O7ЦE�v��U���)�g���wPm�ìD|g�_��闶]�*w@�Z3�N���kL�HM5�~oP0����0	��?�����5p�zZװز¤P�����X���?@���i���J�,�h��U��#g�hVwu���E$��߽�m�nj_<�6�!V;*�x��A�G�pX��$�%���r �|�8�2m/j�D�&�E �1ҁC�	�'���8��2,'A�v�:��w�Pp�qů���r�h7��T�m8r��C��'Y�����m�\� ]GS��`qJ4`/؊	E��I�Ƿ%
��F�B<�,�!yR�S�3j�^�!��I.o����9<;x�nʡ4��!X��w����omD2����(c���j��S�5T���.6�B��-x�Vk7�oQA�/�����O9�V��K���=�xOv��Ι=��o�h�*m�]��-J���)<l��������������Gp�	mS�ס��������=���ӈ�MV��F$m��E<N#�7E��,�����-Q��e���'l�s�O�D���%�w���&���JwYEۻ��GTday
 ���wS|���n��BGj�n$$�2�����>S^��S�LY��5��r�+�3ePb�xb�>���A+�ZB�o��$���s��ph��$�g/:�/+O��U�*�GP7�T����t���S1Q'��s(*����R��� ޸�j0^����C��pnA����U���B]5b�b��%I�Ӧ��8ړ��϶ݷb�V�kiz�����(����T?���䯣)�Nij\� B�h�2S�r�Q�Jy�!����<^ǸЩ�c�y,��d���F#�ը��O��H6� �7}+6�h�+�	V49��~�1�G�:�D�B�x>X<1��Z����[��9����h���J�ՅM���g!ʑU���K�՝�oő���kQgP�??N��cZ���S�Á�Kx���*!v(	�P��ΐ��Qm"�z#�J¥!�2DU�$\���g��ٛE�^bQ�0j<0	Ք�lۈ2��?�Bil� ��%�@�ڡ��˻��U$�j�ܳ�R�:��C�����j�?�gE��@��,F��~fr�_��<�$(!�K����嗖���T��2���`r9�GH�:_j�z���Z����"v�pY���ep]��&�;�7�_w۔��Sʄ��C��%t~�RT�j"nNe[�NO\}n8Xe!3�@�T� 6����&�)�n��(o��5M!n��a�L��0��oP�b��[�(�[���*�F����A�nuL�p��i��b�4�X�;f��@E�E�
10�zǨ���N$���>B�����Z(w����{�X�O�Z\�Pq0`�JJ��lR���GE���{�+ه9��F"��Y}����ٞ	eK��,����,�
��}����#b����\׫X�A$ctM�	���.�V��.Ve���� �(�I�wnUp�����z���i\;诽�.\#�
��p}�+��C�7�?��m�Cj�@�/�-n��ur*G���>0��a|b;�j���#̺�����8brw:żq�V��08Ϋ�~%Hw�t���ŧ@��sC��O�h_
��tp
�[D�Z[ᡈ41k�)�}���iK$�P��U]-�0o-G(�����{�/:MħR..�~1��?T�/T�d5;Z@�˫C��mk�D2��&�_�t,����`H�� ��2H��{�/�����z%�谜ɘs����JO��b�W 5UmX��Lk#���o�\o��Ӽ��Ќ����c:�I�$NV�xp+}��;���6%���c�� ��m�bSFZqA��e@q#��዆Rnː�㽰B*�D �} �J��ԫ�dq���l��ؓq`^�-��C�=���!"�9R��L]3u��*+aC��U���β� �,����H�̏r�]�}���
MqJYeL����̈́�S�] �&�R`��]M�,M�Z�]���24�,�_��X^I��QJ'�Ya�X������Y~<0�����.bX����$��E&4 }����be=�5Ԗ�B)�mK��I�)�cJf��#���N�i-�t�N��� �#C��z(5�/�)5Mf��b��#Y��n% (:/W(�j�e�HN�)��X�K���t��-������Հ��� ��<!c��6BT�G�*c������8(07��������h]�P���ge`A��ĄE uh�(���̤���O�&����+�-�Q���P�P��������_uv{�E���<Gf(G'��r�5�12����w�r�0��1�$�ż�i�U�8�8�b�m(���B9�6�Q�[����h{�S^#V��>G�m[E�׏ҧ�X�����ۭT��{���X|�2�ƾ8N�}Q��L�؂[mC��h�9tq�~~�P{1�x�H�}�?K:}+�(��a �V��w_y��T姏���q��d�����=�B�~`�3���f��Jy�Q� Z��3*6�\^���bH��T0���w�}\��8E�->��>p��d3\�a,��i�x��\8Sx���*��ނ��):\xF�Ԡ�2��"z�Q	��l�UVw_��=��⋖D �r}=ԛ8".P�H��~�Fi����H��@P`��"�ET ��h��|n�-$3�X����e��qLލ���6)�@��dND&�zd)zdCY�EE6�G�|�vi��<�c%ϫqH?��Ş�Q7b��N6а�J������{�/J!�B��+���au�I �gP��	�<��	|̑�Q9�N�;|�Ro�E�����a�hC�.��7�-y3�]��x$�˸g��$���`MF�bgf����bY���!��-�td��=�;�5H�'J��/���6ց�2���;
*��>V(�z�3\���k\_����|��ѫ7�qxu\p��������8\�̿��\���fd# h�#Ú�tX#G5`dhL�Nۚ���U���zZ�o4�w��{r�֭�O��@׾!��fu���Α̣���Z�(�L�p�C8w<6F7��ܗ;��S1�Ȯ�VGUTU�Ma������.�)��v_풲��{`L��S�t78y�#����ǐ}����ۓ8�o�����SPE�권��V�rl1]m�|�~ᔢ?HF��e-�pe�7�X9�ܯ�?�� �V�겄dܯ]o���G�ͿP|��oŗv��������o�;py�|>��>�e|_'|��.��Z��
ŷ"�5�fQ|�Z��I�Mn_*�7�|�)��Z�*�.Z�wb �wr@k��Q|_0ǗO��A�P|����_Wym���p|e�+��+����v�E|5_f8>�i�������w�fTYi�\*�K &�����������ͨI����(�&n&���J,�Pq6�3�U
�y����� u k��n=_����s����	������c-����BO�l��ԗ8�~��+�Z����'��Veo�ȀtX���
~O�z�:���jJ�W�����������S�F���7֨o�~�3B�'�[Ƞ_O/Y�,-ሗ6�BY�3��nA�^k�t��4�f�o�v�i6�u�H�����8�_�fF�)�aS�(���F���7���}$�p�p��I��P
/a��,7�d[ӟn^������ǔ����k,矦�[*g�Z����^�Pc93L�I`���L,'U3�\��Py�Z��ג�l����P�@��_�_��U�y���V�c_�u�Y'���׾M�����������m/o���L�KP�{����Iy�Z���HyE���g(�mZ��~Jyٴ�i&�}�O)�UZ�]��I��n5-ϭ�w#-o�Iy��촼�������v��uW��c#)�����ڪ�M$���VޞDCy_l4+ok�R�FZ����OT�[F�{3��BcyKMˋ�ڐ-�4�7}�5���1۽��zL��2b��4�ȾJm܃!�^���~Bs+�6D�ז�;����j�Aj������W���Vpg5k)�zh)V���e�>OP����?��:�-��j����n���滟����;b�7O��O��'�/�A_+��,4ߏVY�{�<?�!y*�k����c�'�*�j�`%���YIiz�@�a5_��m����H֭j֛i֧���1������#A��)Y7hD��v������4�Ca����� <<�J����q�a{R�L
��:���W����O�`�W`�2��
롰O���W�e���T�G(l��?��߮b�96I���V/w��c�'k��	�*
�&VT`�d�e*�ޡ�ꏩ	�}�7�����Wa��* ��9v��������R��(l��+�L��(6��FS%6#��N
���[�2��v��7����`-T�ʋT؅���1�]�j����Ma
���a�v0��L��La���am
��v�����Ja�acX'�]�¾��������`G2؉*��v6�m��;��&��WQ��)�ea�
�$+���ܓ�>Ka����z�v5�]AaǆöS`E;K��Aa�Aa�_ޯz2���@��d@�Q P1(e_���}��G��]=ȣa ��d���x�I�=ؠ�hv?���O$S��r�`��ZA���2ȅ��N0	�}.h�4u�b���=�<J,%�Lw�
�t���=l~�QT,K�U��|H��,H<�������7V�-ǣ�N)��i�N!�;p_��|��9�{��A��h��
�Ò�5���o��_q�4 �b=��b-م��|���� ��_�=e�U��VQ��ﴙ�-�����3N��9A�SH�����&N_��	�A��INt�u��J� �}�H1���B��Bp	u�� �7�'o��pQ6F۽G���B���t�Ž#�>�b &M<&g�A��l��Np�� ��H\q�E���q�*_�#]L��7�ٕϬ�葖J�U��)�K���xO"�㽅�T������K����V�adZZNZ�od��q#;=�����N�^���j���,-z��{�s94�X��%��jܑ@��ے��V�@D����cU��p�6Y4�B����ĕF���Hh/��ry��}w�P�U��cH&����X)_�p*�Vcqղ�-⾔T�ؕ
�t�yd�_���xZ%@� -Cbi�S"��������:�
:[�H
��������d�7(?:�nl�'�
���-�{`=�CD���ک߯��h'X���о�+�<�O���l�w���e���6���Rt�+�� �/�1�k�Œ+���k^_�����ՠ�;X�N���%�����4��ض��ǵ5��p��ib�����`0�~�'��?Eů������[��=썧�ވ�����?Ot�Rw��"�����hC�J�wh'�L��.z���:�YJe�};>���)l~{�$_3����I��(�R�'�A��Nu�*r��[���O�݃�4r�ݫ䢗�'�M�gܽE)�o���h2}�NrV5�s���������WL��Lޣ��hG��׾�`+���?R4�t��4�P�l�:��=��}��G��׽B��}SH=��8l�N���;� ݬ�h�ct}0��6d�g-�$dX�U�w���R��*-)��]�J�!*�O�#��6��,�Bm6�<3�OU���q�����A?�b��J�2[խ�@�O�]��x�����M�z2��-��6��'����I-��~��kA*���T�p|`�[�<t��N�oO\^��T�
�/��Kg�_�y�:�����`���F��i��J3�O@򯥹���|�tr�����}?����!����1��%�N���Y����%�s��ׯg�Gp *�<"jC��N�hoı� �Ȳ�X��jm�o��|��;��OT��ǧ+��I|ڎO� �6n#�8���KB��*s�[�ܕ��!�Em��}�F�8ĝ�38�?�&
��Ri|\�4=�h�mxfYɽC�W�D�r��NH��e61-!�&>�`���%��$G�9��p�|�88i	��'�$y��ĀC,.��$ �o稂<ȈK�I���L''9�2>���3B����\Ke����%���w�S�+uJ�K��r��ӷt��w_dq�!�	Ȍ����w�T.�C�M܇��i��{m(������{����ߎQ3搜	���&�m����9�PI\��UQՈ��E<���z�,̟����0��s�
L�.+4��e��?�d�8��>[��S��]U��B���0�P�����hmN�Bw��-M��=��]hܔb<�G8T�iN�K)Ҙ*8a���5�B�
m���R�z����%y�#��
��2�P�UО�8�Lif�o���-7 �mZ`?�&��[v �����Wp��n��1� ��a�/p��t�^�*X��,�V�P?5<��	/��έP5K�aP%��O��>����LL�c4�5�q��O��	�j�p�&\Fǀ���k	\Oh����������K/d��R���E7��������O%<U������M|�&\�	�k�D������Vx+��!=+x��h�a����c�_��^#n�2E6G�!�xdC�Rߖ�Qb� {"�@,�=�8�Wr����!G�h����7��M��:Z�9���⤕��!�9R��F��&61R��G_JS*�SJh�ea�c	4�W8X5M�Ѥ�{}�*�p��1��&|�I��Ѿ�&��hLXA�P�|�.��bͱ<bd싈���P{��ن�ct7Nl����g/3Cr�Qe�H:J�}���������I��������new��ܗ�|��_��^n��oA2�>�W�����E>�"��C��@��-�W�|���p�H��v��M��`'����tB$Ӂ�r׬�4��pX�����z<� tK��I�|�?c{t(���	VɾH�JP�%=xV����^�&�V�u�8�����(��$L�����QQPQ�RQnQQ�WQz�������Z9�����������;Az�l+\_���a���:�.�|� O4��YL�_T׌��ب��,)���2�UVh~�5}V�R3��p�2:���� P��~>Ĩϖ}�t�u�{h-�D�șل�9+ꢜ����w��R�غ0XMnp�}\�����b!B�=��7��ݗ��!6kE�?�-��FU�khʭ�)L�}��T���r���F�Bf
��>�I�jk-M���1�)aGxA%�~3�WP�u}:mCr+:���EM�:�XfH���'i�&�,-�A�+<W%��������t��X?*Կ%�&N�w�_]�-�z���r�/���Z�(�bE��"���T�
�B��|���|�	��P!���u��v(ܚ��vC���/ȁ|��@�,׫��M��]dU�,��+��#���m�b�\v�=~�{��������]���L:�K9�.��D<oc�9�.�`�B9-V�U�0�/e����<�]�{p��Kbb��yr�D����'��X��W5.ጯ2�ǀ��)���D2�xFn_.�އ�E��A�SQ�__B�8� ��,aR<�L9nH׌��`,����b�E�d�����&���)$vOx~���|�rEx
S$1���H�"��0��w�bQ��ٌN8��L�w�
t��f�I��0���4��3U�7�L/E������:M�+�3U�(���hTO�-�ꉬ�����e��� Y䨔�S ��s���q�������h]�#}��u���f�����a�92Ob��)���9�tHO��<k�[�"P��C���DP<�q��8��9:3�YQdP\9UaH#(�+?	ݗ�o�
���?����3�M� �t�gQ���J��\�a�ȝ���#u�h���H?!
�T�N��΃Vr�p�t�Z�ݣ&:�j"�y�����N�^�^�x~ݠ�����zE�MG���)5\�N�����iԢ��b�N-��sZ׏ݟkE?NY�ӏ��~�3ޭ�ǐ��|�+��:U;�7Վ��GU��b�o�.�,�U����C���CsZ��P��e�yN-\QM,�~C������ )e����X���Ŕ��JYҾsƤ-�8���nӤR-����:oLY�R�/l�R?�ġ})�Ʉ��9�(��;�ϰ��]'<�.����T,�����\���Ov�9��õF��?S��3>E�K�?���3K����K�*g��J����1�f�4~{pːW�鮥Nͬf��.��?_�C�;\�ߖ������V��o��o.�.D~KT��,W�_��L��Qv=zj*��g��N�����Iew�vxB�[+���p~�t�"�bx�"	�gL��l8�"���$E�o
KBAU�8��Qװ���R|,%ʘB�"K�-lK���P
u����N�i.pY����"�����44ـ
�&x����\/$E��8]\2y��dNlQm��c�dxUe�؜�(�4)e:b���tD�FG�����TGLe:b�n�#&RQb�͌���ÿC�a5�(��G�J�V���Δō�V�B��uZ�O���8S}����{GqJ��,��9�'��oIdm������p?.���Ԉ=Ɓ�n\�������g5��L�����C�q��dгd'>$>˶O�������������U�6ڌ�ݢ�ש5��k�;���w̫���?T�F](}_�T��Fߊ�}�y[���5��k��oX���.��dB��H�S�F�ήa�}Y����	}���3�ㄬ��04��by�=��n�л��ާ�� �
T�r��5����m���(e��I
e��Z����z�mNq��y!��>�>��B�2�F%ӝ�q-��6�[\G��0z��wF��V�-[��7�H/��'D���.�^�B/t��a)H�'��T�+����V3��z&D�m��t��{h�T����;!y�|�3ĺ�`�}��x��U���f~:>|<G���y�!�.��Ì=w�B���L�ޥ�՗($���}G�"��q�{�j���n�ןw�d������E��4��K�0cy�]F�}��5��W����_w������Pu�}X��`>E�#D��LzL��t�`���J��!�א���A4-�Ba^5瞀���U>�N�u�4����ұ���������<�ı�6�Ny dK���-w_���?�2����G=�H��mgҽc�����|G����v��>,z���zk8�D��0�&8Ń8jO�߃�tu��=8JaR(?�����rP�?|�[BS5��F#���G�7G��A/� ��w�
5�.��.�_w��bl�
~�숊���v��G�k��l���-��K�K{��h7ķ�~Z���c�G���LO�7*�0�o�d��J��Flⳤ;�ۤ�?9�Ŵ?���BQ����w��!��c/@l�
j�����7݅�T&
��ط��?��Ap�������o�e��+߈����}#"�����L�O�g�����5	��_�9� ��Rd�S���B}o��4���(!$s�y���C�/�?�p5��ʯ���M׃Ho�c��1��0T�}G��0���?�#�-N��R��O	C��n���q�`���U��%6~'2ԓ�Ud�wT�6��ۡjA����k�6��a�����'O��?�6�@���(��̕�*�Os �B����˕-�ʦ�ci�~4�Ԇ�PX5�o���)��m�a�n��H5�U�T�2u/
v� ��7�볊1�4Ooٺ�0w�[�W�he
�K����/M�%M���m���4�_�T��I1q՛�ϰ�W����{������`n��0�-��@���{X����$F��wt$ݿՖ�EmT�j�����8�؈{҈�#��*�
�W��"q����Ild�
e�v�Cw�w��h;��h?����E�4�:TK�ޢc�%�`e/��:m�����4qqv�Z���dZ�}���j[���r�$�1��9)��s���VC>ê�;��I-�x:�X�i�F?j�>�p��Fo|�C8�~
� ����:����A&=�hO4��l��E�^��6V��Y��R$h�}�:��<
�F�m��@�IxP��Br��/�D����m������l�MS�][b�ޑ��y���N��KA�'T�O��ǨD�]5�FBl<����8��$vv�@d[�Z�4S�ؖ��~��g^#�lF�0�a�>���}�l%���'�����}�{���
` ����ܺR��C���C��O�;B業;��Kg��r�}�oD�B�7���}#�,����h�Ϫ���0;���by���;���Q'�Q'��?�����1qS�����Z�`�s�}/a������}� �U��ijW�J���Q�)�]�����Q��]u�;�����"��5��Gn4����`_�=�����u�{�L}{<��׷V��ו��וF���5�-O��bJg_�'�۲�1��ݺ}�|�U�:�h_��CUIҾ�tPo_���!�
�aWn��5�j_7��ו�}�/�,������M��n$ъv$)�~$)��$)��$)�%�J
��
�-�p�̺5ͼ�C���M��WT�4i��y�{\�_g��}{��/}Yc��f���^�����`0��r|Y��5{����f�����U�x��b
���� �ȊP�c|P���P�_���~i�,�"`�d.I\�K"��J�DD�!G��MB�E�3`%� ��L�?�Z�G���͝?�(����������%��;���W췂1���^n:���s����9��/)�|�>՞W�7���̞w�ժ=(J+��s�C���U{�s����a�f��j�,�6~�Nfә�Sz}n���T�u��aƺ�%Ŝ�7Sgή27g�/�
m����+�ٰw�rՊ��a�J^��?~P���0��������טӿe�Y����J��[�K*'�_kΉ��4�=���=~��N�Ǿ���O�[�Ǘ.������b�=^�j���^�=�����+Q��_�1��[��7-m�����e*C���I{������5:f.e<�M��cc��e�]B'u31�š���������]+��v٢k����M��m��i�.U��Չ�C[���&������쮫��s�����腎g]/@C;���`��,����-�wgW�[�E��Am��ی����'^cf�����د���_���/�z��;U���׸��y�E�����_e"c_��޾0!��
�G�^PŨ�/���V�ͯ'<Z�)�xe	Ƶ���:h�2��H�-�hF�<H����WI��D���O��ߪo���OЉwq1�2kj��w�s��7�y��oԿ����%\��=��\���G���1�|SZ׿���S��wx���G}Z׿)o�-o\��b�\`k�?�_�?*7Y��������E���7����a�?������������š���@>�S��G-���.����o��+��5Y�/�^�/������g����q��*���ӿd�B����/.�Z��8Y����+���	�t"]'1��0�u}upa���5��|F}��H��^���e����c.Ra�vR�����V��`�W/H*Cm{�I��/����:n[�x�lR����y��?�/�Z��Sc���'ք�����?D����^��]��(���b��r����_��h�e�P�����-l��e�ׄV��7�5���bTލ�����P�EߕF��B՞�[�;>�/�-PI������/}�׿����{Ⳍ�A��3���wN��w�Q�|Vejܕ�7o7׿z�
���q�[׿���S���s��]���Ų��������H7���i&�ա0��3�`3�.Y�Z#�i~F�n����oe��e��T>z�ଟ�?,
w�b�ay�F'rg!s"W=�u"��9�_3��O������ɾ�<Q�:�G��o����ꗠnh�}B�U���6��v�����ωW�e�n8�r�z.��e��3���)�(W��C/Q��u�s�y@Y��ޅAD���9d��W�.�Ώ�oqk���!y{	7u��~����A�&P �������2Oɫ��3B�M���W��t�$�q3 ��"����#�HC(�
�ϟQ9��rE���Q�}T��o��t* ���������
���[I���Ĩ�"�Q���.��T�뷫�̽�Ϙ�3�u���ӭ귩F�vc����.�����!^���×�x��4�a�}��|���7%�K�oJZ��1_u�
.��S�Y����Y��zJ�z�P��ռ�3�?�c}Z�����G�o䋶��-�A{x�T|�뼐=��8Õ�e�Ņ�l������ޞ�%�t�jQ��S�)~���SK�ў>=���1cZ���g��Ğ��q0���<՞��B �^���Ӷ�a`O�ݹv�ߛ��E��ɥ���>?�Y��ѭ��eO��=N�,�Ss���[���|؆�Ts�J��f_��~"��L�;���x���RA�.��S����O2�|���]c��Gs�����*�jL�5��41
Z�<�ߊKt���wW����1���O*�_G^��׹����y�[������ט���Znn����:W���~�_�jg������g��n���;����Q����j3�hqN���sJ/`�k�j�6w���s�6ra�s�������{����?��O�ϙ�����oWk����fN�E�IA�=P��As���5N��B�i���4<6�}��ae8Or3.V�~��]w)"����n���SCޟ.�[�'۷
R^�S�i��ρ�O��iBAi�,7��t�PX�"��D��GfTzRn�+�+QcrA���s;#��X��;��K�B�r�P�$�~<^ʍ����:#��|�K�G(&]>�ʍ�=s�Џ#H��1i|��|�|TR���Sb	ٌ�Ō�w���#�]��{���R��6p-}/3��͟�B~�ȇ�}�-�=@�M�}����f����) �7J�tLͦ����O9�}߈|ڠ����P*���P杦e�U˴A��?�n�L��[�J��b��bG?��%�����"�1-r�'�lif�@���>!ĹXNi��h��Oh����WE�ߟ3��%0��QPO��FЦ�4����h�O��=��o�T^�W+Hѧ�P/��?�6�%o�(�Ry�x����^ajT��������Lr�����sB���K�*�<}�x�ȥd4�K�)r�K�uL�6;����x��xW��f�K�c�	��kq�)�6l>��i��uh����_|�*/��@[���|d"����
��2(�f�8�2��,�H�KJ�rJ�?�1i��!R�QR�{�@�����-w��&�}/��u�/�ꊞ�!������:!�(�]ί%�����g6!c��>��ůh���5��� |wڏg�y�^K:~9ZO��_�=�T��k	[�)�W����ߟ6ړ2|q��^�=G��n�_-���>����`d6ţ���V��J�n�t���g*wH#�lX�k�SQx$}$yQ�xL(��?,TU���ކD��J����)n??�)�R���׏0rB�з��t���d�h��p~�T��؉�%7��J�>9b(pM,����/q���#^��$}�C6����
}���{���bA�>@P�"��O#h��	�~��8?k_��]�����6�A� k|`r���:�Þ&y�<,M�:���Z~a�K�R-�N����d"�K��T��#(�5#ȤCDvO�P�"C�6��%P�	՜N��<I��G�zƜ�,�R,�B�7X�QL�9w~�����(Y��|T��A_ ������;�[�A#T�;�9��E�����C��w���1U��������ۆ����E&"F�K񇇓������9�`�?��� ����W��t�`�7�|B�GFm��c�;�<�:�Q�z�	�_�7��j��eK�b�C�Y�g�B	�(��}O���Q��O����oE�$��������z������O�9�?�%~�{��1G�BrE6C�q'���G�R�;����dN.���A�r��Z�=�#�[��=�����(�u��F��y�8��j#�:R��6	���|�A�$H��B$~�al<��i�^�/('�j�x�i�X0`����~ThK����L%K��2/�	������յ����IcC�Db�Ek�Ec �V%B�"1�J����)P�Hce����i	���&mV��T��'!/K�N���]��R���'�ԏ��m����ԀZ�I��`��w�y�ۚɮ|_��H<�='CE�"�1b�L�d�d�Cf�q�|��Q��B(�i}!�N~�R\r����q |�H�E{cA��&O�A~��'�������T�I�O��Вzd���B. >�?��%?r�Kvf<����eCߐׄ���ܟ�_��Π&R��NU��I�S�|�S/�����˛�?z�YW��|�rLP,g8B��)��9��]�E�/�H��	_r���	|����.��v�$��x�E �@tՒї���K��c�[��J��Q߈y'ŦB9�B1�_ԗ��s��wF3^�L߷w���F��+����e]�o1�r/ᵑ6**I�(����Q�㩕��
,��'8I�m��Я�P���U{%��5���1[��*U�3����
�o2��1��m~�����j(�'��#���G��*Պ�ܴ�z{��9)��df�M���3ye&,�ў���g� Z�'�zB�K{�|��e���C�S���_ñ1#��42N�]�������ϡ�����̶ު4��@?!]	q*�#�+_�
�o!���6���
��n%����~���'%���y�fBKzw!������pb���%�%{���H���Qq�*L�仓�������C'M�#)�^+~z��bEG������iⷐZ+� :il�P�5i]�ɠ��t�d�����_������H�&��a'M�m��Ba�D�`p�����NZ��k���~�&�
���dP�D$�8�~D{]��dǉA��iW�2��8NS��XP��Ȫ��޲�!mؒ><s�4@�f>G��~��6ԅ1�h���@������X��?�2��/'�K���)BaU/��pܭB��~����U�t� ͆�ƝqNix�S���Q����ׂx��[����~����a�X}b�C�:�t�K�\Rj,�+�����������	�O<2�auPH�+8R��ZcR�d��B�YC���x0XJv���0\�N]�����L�7�/b���;�"�t�}�0N~Y�ϵc�}G���F����M+
8�(����]�Յ�p��E?��F��O��cPt�ݎō�e�s6]>�h_�]����|!�g�6�\�]rHP��/�K��������ס�g�,n�h_i���h_��Y�X��W�Gz��X�/�|j%�@#Y�qk������$����g�x�n|+���+���2�2���
6co�?��9��j%-VA�Iħe���y7�c��|��� ��U��4�l�� o��c���SicF���e\s���IVhLR���B����4�R�RM�4��44�)QCSJs4%R�C4�2�>n �SmLi��4��.����t�MVMq��d�4Y	M�"��˓��I�Dq����H����0���aD��CD���D�$��7�(���W��"ڔ���ZB�.-Q�*Q�̈��U�QՔ(�a�&���Hέ��Sr�9k�䔩�5#�DCNYs�PrJr�4��c �~�)9+)9�	9K��,W�YjF�OC�����Qr�����7��^���Sz�z�Zz����虪�gNs�L��LU����NH�s�����3��3FK�8��1f�z�5G�@�Tz�8��(�#�u�'��3PKO�J�@3z5��4GO"�'Q�������z�.\U�����+�J��ő�?)\֑Px#S7*�5�q�$�� �i�k�P������'����ʱ�Fi�9Bi�����C�4��B)F(%��R���B)���}o��!�X�<)�f1m�J^5���zN���*][ϙ�q�����*���1'� =gJO)���гJKO�J�*3z�k�)i��唞�*=X��W�M��mJ5�F��y�/�q)i�b��!�?��ht㼋0�h�Ő2B��H�=�"F�RF��"�m��C���<#�;E�|��Ԙ��ER�`JoM9���M��s������!L9j	�L���a�S	�j,��u/����5�}���rq_%ݍ�|A�,/��\�s��}O��&p�6�M�k�M�0�6�8��D�h��$��i�z����r��ϴ�,� 	k�	�~	%,�&��@<�M��$dh�c	'�NmwhSF���r�6e��eڄ	��`+���������o�/aw��?��34�xUi�_��s!��O���������`0��������L(\�����0~�,*��Q׫߇����WGnoא۫�䶬���+��[L�����?�ܨ���ȍ�g�C4�|�d�3	@�8����%��>���*�NS"#%+�Od�M/����|"c �ts:���g4%��e�4�C�2���ӏ��������69EeE�cY�T����0�8ųc�t�lk��(�>�����RpJgY\�.�Z�����ǯRA��	Cq�Ϗn�m�`�i,�i����ueu~��|ݖ��l�9����(�#l�D�#�N\�&��dz#��X�8!�L�a8�e'3BN^��w�!,@�����|�,F�8��%�| ��KV�Æ����R�~ �������\�q��f^����:+��!��%#�}��Z,��j!�K��4I)b��&��m�`��bO�J�G'̦&JB��+N�\��9�2��25�ђ���%�_�'����x�����B���ryoC�,3=^��g���Q��U4���8�&A%�-�P�t2�F뜆�ȤTU*a��*��Y���K7�QKf3jt��d6c;_t �,,n�h���fԒٌ�|�^]ܝdv�;]��̎�b]|��ّ��|����<bٔ�I8;b�� ��D�c\h6c%Nu,x�Tn�vR����%���9��p�-xQ��W^Mqk"�w2��� 6c�$c�"�#n�劣�AxF��b��-ţ@=����o���xᄋ��_���M��������	-W9ɒ��=�(�/�D�y����g�i$�[~#�W���l�ch5���A���0n�m�<Gd�l��/[b��#
(O�%��5�<a�a�|(�s~Y�*�t�O�$u�n�Ӻ|��}=��R��Y���/����ͤ�>��z�����:�4�lfj�Z�Cmq�����-� �q!�Ҁ�#E��h�)�n���F�s���1j�D��N[�&i�-������)u��g�4J]P*_�RWeo`T6�����Z�(P���S�cR0���{�"����x���2b��ŒY��*d�3�2TN,����T��vE(%.�66�jK�G���V��FGZ	[�t*���i4����8�%��t� ��c�h\�d��V�Y�
�JA|�X�RZ/!M
��m8um�d��B��X2i�߁�����!Jܭ��u^X���7��
����;h��j\ӡ�?a�뱥��
\�4�]��]�-�@����~�y+G?; �;�c:#�^�;����?\��I���X�?h�/@����������`�T�"�|��|�%^�'�և����͓� %����()�#)��u\H�h���
���B��(ܓc�=Y��!�J]�2?0+�� �b^3+*�Z������J,]Q�����1�]Q��BWTJuqcpE��~��A���nF�*�r���hc1_e9F�9:��lMVYiV"�T�/`��8u��FJ�_���k���IrF��FnJ��`�z�� ί� rF�1D���LM�	>���c�K�3T�f��C���/�:�oד��:�~��:^�<���T�P�y�`o��R��õ	�y��0�F�p�&~�0����Ϗ��}$�������h?$d������يn~
��xE���AJ�K^�{���9Xp�j=��x�����(z��FT�f�_OxͬƳN�g����ыt�h�w������׃׷縐
��y�&9�Q�,֘�Q�2�I���S�֠J������#{l5���ND|;�%Y��6R��yT6PT�Q�_e'�'@v	m"�~�@sײae-���*{�8څ�4[��OT�0v}��(x[*0)d��
|��!q7UF]NΆ(;yj�*�S�l��bB���)6������XiL'�� �t��y�6��C�m��.S�n���gi���c�]���6�CO�E�)�|i�h�-~�5��u6�8MU����f� sN��a�<d�t�݃F^���d~m"M�����VM�G�P���,���.<��ۻ����N�����_�u�_~~��U%Ȕ���5�:�~���{*�D�C~��׾�Tc���_Ђδ}����Q� e'��O3;3W��Cߦ�m�2�sj3��U���Μ2C���Ϊp�B$����V�ّj�`BF�1͔S���53Yֈ��b#��D��%
��I/q5)���kɡ��������F�����XX�&u��l?\��b�g���X�m!N�U��V����{�Qnⶸd�� 4QA�V΂{zv[��QA����<�v�:�y�����Mȸw�D^u�~�O1f�T�>���\�r���0#cBŇ�RY9uXc��4�@؞$��r|�PRi_�Ao_�}8��� ���
�/��r���J�qRQ�-UL���S�m��	1�iF���Ad��Ŋ����4ԋ7��&��jSv�D%��c��ud��^�+�e�� P�k�cM�x�\	��v�Q������^�D3�(�{J�~=��v�$�I�īƩ6$��.�� iμbt�#�ѻ%����S!i`���cֲ�.S]��6�l�uy�d?4�^�.���8�A�p�<�4�9�F�<�c�~UC�+ȫ�ͣ����j{MA���G��E�ī��9�NA}jK������S�-�+�I��$��?�Pr���%�e	tO0t�*�V�����p�ZV�r���El�N��b�RrNQmY��	J�U*�L�����_�ab���}�S�}:e�]����NK�8�G,��"9�$�D�����Zi	D�O��φ�9ML��C�8�.t��.C���BE]$\ڵ��1H�zUN�g��ipF����}ށ�ra#��\xq�B~���;��@�*�6ʬ�Q薥i�ץ�ߣ�!2�Y�[�lxi�|��p�&.���,;��@�tO���7��6��K%�Y��;O�ڄ�	�L��'��A�krH��$�#ƈBm�<�tO��S�(��P�U�Ry�Rhid��Cʠ��YL�� ���}޴7b)���%�<M� �[[˩&1�o�&���*h
��X�!ȴvje�l�X�I9.UA������&��O�S�4j����TF�+���W6����N;.�!��~��.X��؞��΂�R�4��#!�3�T�4�8�����<�0�Tʘ�I���)0�V�W�q�%R*K���P��̷�I��.�����#�z<�Bxb��6Ny<d�R����/��̢0u�:!�`?fPd�J]J�&E�`�.[]s��v��	�?W�j7T�_�:XS�۩�n��Cs�d���i�|Z*�ǫ�1
�J��6��N+(�h&My��RCgJC����A������s�T��:�
��8��Qc��!�:��cd����2[��������۠�9º���kh�7�*~��?�������I�ZC'��dA�r&-N/{�qj��j6�}589ź��yBσ��X!V�fX�P�1���6���*��4����l���T�����bqr�v�T~iejc��O�\��y~��B/�ï+o�<-M����=�[�ߡ���s��s�h	�m�t��O���c�t4�ʤ�����s'��1��cgD~<	k�o&	e�L^�שQe��������h�[���DC��4�ATQ�ȷ��C5�3w�:9��ED���5��6��(��>��L��d�wī=<�8�i~B
����ZB"�ON������LB,�;�����!F����G�������G8r���%��q��l}��l�7x䟞L�<[QN^��(��5�����S���#�A�㖆���)����t3�Um��4��t��c5
n�]�/� ����\%HC���x�FC��d�ٰ�qx������� Ef�3���_��
������J��y�(frW�qJ�B9�$x�sڜ�k����_�*�;EO��G���_��дoZBBX���I�_:��;/�c6�[��o��2���`߅��."���1���/%�/�����e���F�W��7��*���/!�������_J��E�ג�u俌��'�����俜�o&�[�%��&��������!�_��]�7��%�ߓ����k�z����ۛz�������p��v#�<7��\�a�ki�1o���.�����,��p�W��x���.���C�#1<��]�H���a;��a���$����8N�pG������+I�/�e��4��54��[i���h����p�W�p;/��h�h؂��4|.�R�Ói�w����0��N�� �B�ݘ�ssfL�wό�̘6->#~�n����h|Ό\wƌ̬����3��Ysfee� �$�Ԭ�$#bx<g�ۓ1-~�̜����I�0����iY���)Y�x�Ԭ��Y�3'��gϜN�
�-~D��J��\w����I3=3&�?��
����S
�sfC���S<ӳf��gfǻ��ʊ�6R{s#�~���͜��:����i��*Uf����$�n(RV�,2�bΌ�gff�s���ܽ�=#�����sr)e��G2�0-cƔ�<3�9ӳ�s2�f!Rh!����1%+>q�=i���3Ϙ�39T��ɢ�Л˞9m��'��Ț�5;'�N�=�5+g'd̘<�����qnUe�73�2�[�P �B�B�
����3:e:��i�B%�Inf�fr�M�� B�.V1�]�P0*�V�jpq�;*h_��AQq_v��UE�?V��9�{��;�����~>�M��=�{��s���ޛ�fziD3��k�
�J�PX�LV�QYm�ݒ��GO��3�P�����2U-�2|`j"�d�M-��ll�O��T�*��2-�M�3C�RnJ�YL��U������7d{����Imћ���ሮ�-ޮ����l�Aw�4�5�gM<�\kQ�e`u�ʦK��spـ��Z��E���7�����&M��%��mZ�mc��$�#/賑D����M�m$��bW��njT~eE���e-2(�T%͕AVJ�5�����^��ךDP�i֏ftm��Q)�km�)�P��0z8�H��ݨ��X�LF[S������i�R	۵�vk�˚�3a�3Z��U�:��Nk:A���0���Q!T���ÚJ��M����d�"etC2;l	ʁ��Y�0�o��1�����Ng6��ajf6)�����t�N�{���у:�Q�撲�S��F�[��6���t Yk�����Nh�P�g��l�J�R��ZZϔK���e%�"Vˮ�%'͋o���j-������v9(Qi���N���"��c	�Fկ����v#/F�"��f#Z9&�	i}��}/c%g�"�FX]���V�զNO�����.�Hy��@�d4RV]S��T]Kztx�H���9�u$���&�6�Vc�U�#'Ug[�'Z�V���Fe봲�6�����-P�����P�i10��l��nꪭ�N��R��%���F��/f�{�fT�����:;��>,���Q}��.+�QO��[b1L�j�p���e]PU*{�JX]u<�ZIMeS��4�Y��������M^���b_˂�`"�毓%R--����8�����3�hO�7w0��W]�@��G�_�ۧP�k3C�<���g#����n7�{h���)`
���v#��&e(!mf2T$�͡%yO�U>���%�f����-�$�h���M�!1!�,s�蚐Y6O,��ӵ�d��R�A�ӆ�,饝i<�l.�b�\���'����MU��*ӫ�22g�5���P0��05�%��a��-[W�J;2��!=�˔�آ:P��'�C�˵�-jZl}�Kҳ��e��EF����	�A���E��}��^^m��ɕF򪛫�|�@n>U�[q��e`�,FaےCb[-��x�����ԙMF�1t���\A�m�`R/�Ñ�.��}PI�r��Юo�ɚ&�7m�L�k�av�=+o�[\��a�i��Ȩf+l�a��Z�h�-U���+X�x]������F�A��u���5����}�u)�i�j�[EA��'N6��o+HO��ԩ�,�e%.�Y#�[�!v���f���,�$���e�e7��q[6�;i�M
�G�rU��;yTҢ�I�<PX�\�-�����aǈ6\��"-��R_zɵ�v��X�O	YrmR�y�֬��u�S�,�B�#�C�%�嚟�Ԅ�֕⩪�3[�v�y�\H��+�(�ް< �p��R�Q��`�:��������tw >3��u�ܖ4��:��C*�1��ftK��h\�,�w��~��{���۩w��"�ſK��_�Կt�Yڌ,�����e�Ià��̰�e�8��Q�B��8�B&u�>a�pT'�0"]r� �Խ!�g���[5���%p:e$ir6�
��4�_y0\yE��j�y�ͷ�%w�|pb��=���W�|kh�!����b��g�����\��e`��Z@^���H�Қ#����*G5r���o�*�D{9ޫ��	(��l�.��
�lWo�l���gv��uZ�'�i�x4�g���I��4-����W%�����l�V�Gh��#U��G��5�fhZa��ɝJ�T
��i�Yڌ�,�yr��4v�6�8[k�NF��yh�h��H�_@�iM���4�j�"
[�y�WQI�Қ�WkZ�5ZK��3��ү&�Fk�XC%\�y�֒�k5O�Z�e�Z��Z���R$9�<���N�y���o�4������'�S�QةiŝZ�/De��]Q���u�-FiwiM�H�n�ɛ�<�	��<�&I���I���Q��0�ic$���-������$o'=w��;)o��}d�]ZS�=TO�њ��j}��?���8�P]��ܽd��Ŀ���~�E� ���|)�A������֒z��� �y��rH��}H�ri-��fz�Z�S<LuJ��a��Ô_�d�l*h́���մ�g������bB�9�O����^���}������9�!�-[5ψ��}Jk�y~v�#�xJ�`��^���]M�(�v��v�;g���gqO��;>��8�k�MR����Pw�"�I�ﯪV��G'��3�;��67�����ޝ��4�8	��p�{�[�������c��OwΏ����Z�6��Dz�:��<`���iL9Y/?yt���ol����3��|�"C�{~��V{s;q{�;E�wV�v��\�!���;��ŝҔ{�)����mC�s]���ž��z��W��}л�YoM?�`?�=��zꎧ��1�]�Q�$����g�?N�~����Oio���}D=��I���X����O'��U���N�Op�K~-��}�������@�q�'���Z�c�qnSc�S�86K�}��^��S�+O��E�A�-��s�;��\���fG����qa!��I�}�s=����z�}g8��z���������n\	���X�z�\ ��9�#��~�y�����?�G,|7���M�4�϶���k,��F��w��������w���hr�{��7��n��$��4��m���8�ǧ�����F�|c���m��E�����]�?��4��n)�]�?��o���^
L��;G����x������va���
�M.�^8�<ޞ}�zv��OR/�z/�c��G,�:�LW��H�������g����?I/�]���/t�|f�>.s�?a����O)�g��󺽛��J�JG~��X���tǑ�j����u��<�_,����G̡��ҝꢞ:���]�3�?8��d��v{���~1�y.�+��c�����4� �J������ۦaϫğ��u�bM��
�m�|���Y�������U��+��Ok����Ӱ���h��_d���V�o�����)��8��X�j>�V�̙M�1�}c�za�;��7�����6�l��x_9>=F�!�����D��o���<��a?��4��?��K�ޏ����SK��;H>M|�2��k���y>'�Ok����s���*?�\�n>��"��G^Cy^��@����/���z����\-���پi�� �����q�� ��U�x����h]-�~���{�ع����WI�k��K�߬��,����i��|���=�㑳^S��D��#}�}��sh5����:��������k]�8}-���}��F}�}�� �}�Yߴ�_������-��q�R�?5P�N�[���7P�c�w^�����;{.ͷ��ig��o������ �b�Kz��޷8�~~��>��v���5�P}A�j�� �=�_w�{�;_"}C�R_��7��/khq<�ǜ�No�'�;��z4p�>Az���F=���1��/�{�kl/��%}�]R��s�'��;ߗ���J���Ｎv�:h�}��w�7�~p���6I�?x��*ڟ�mj|?�FZy}���!�[�����WI��n�7� ��^���x��q�������O�������}D���{���C���M˿!�Ǡ�����li|�;��kK�����J���Z.��z� {ٿv����������������/��~��]������m��q������[�ϓ�����!��
����6�]�����ǹǈ�|��Fi�K~#ƹ4�po�ǹ�I������K�w_��k�x�ƏsH�ȶƏs'H�{�ǹ��i���q�� �k���8��Ono�87g!�G74~�K������'H��?�Ϳ���;׮	�W��~�;D�<���᳽O[���k�W��R��B�{�5����<�=�o�<���̻��~4��Ϲ���Y����$�6r?�8靀�F�����a����}�������0�����O�l���Y�iCo�����]�}������v����GHO����}-����;Ioz����z��}�/����o2����=�{z�o���=
��� �����yΉ����\O��_�o��|�=��=K�����8�s��[�Կ��ɹ<,*�������������9��@�q��|��5Ο��>�towN�x�~%�F��G��L�>��bz�h���C�ou�cJ{��T�}�d?
���x�~|���i�y.����϶��>�Q�%�V=�@=�@�F��+�O���>�����؏اH��n��u�V��zϧq~�Fσ�b���������9PK�yu��q�ߧɁ?�{���[+���s��>����s�u��b��V�u5��,G��N�G�:���-D~�!�߫�֝Ὣ����.��1?�H�u7��ڭ
/A�c��/��L���|y��<^�xc���sm���� ^ ��x;������T�~9�o�޳�+�ȗ�:
޵�����}��;3<���w�x��[��{�x�����{C]��P��w�[C��(��.xw��c��ˁ���,)��\�Wo�Іl�f�qb#x�9�x��w��ǉ�s��8��"����ԁ��D�E<'�ȗǉx;�x�8�-<'���ǁ���x�t��81��/��vI^��D?x�8�x��Q��ng����g៙>���^=���y�������g���}���L����6�ۨ�v����>�~oy�U?;v��=���~�{��}�!_�g+�-y�<�gy<�g���}Sm�3�.����>�g��́'�c�k��{���C>��C]<n�"x�x?���:���_�_ٞ1��x�'�������^��t�>�5��~8�W��r��~��n�{ơ߱N~@�u�'��<����p��8��7�+y�<�>9xr��x?t������G��~�!1��Wk^��HA�|��7��c����]��cm�i������s౿��}x�^;�9���_繰��U�ש��_[]��X�sʗ�U�׉'������}�ۍ�'�ߒ<^����z~����Z���x�#�9���/s��]�W�n�g���~�-�u�ygS�t��tBz�B���2E�R�T�<�+)���C�|r��IȖ_K酜��2 ��2
���r?���ȣ�O@�C>y�UH�̆����r#dd?drrd�� N���T��:A�l��?=a��G*����~N̮����3���A��5dꈌ� _��&�Y�/Ex /�܆� ���'ށ�~���CY&P�<^6�w�Xzk��m��܇�Ճa����V�lêU{)y4�lϸK{'��N&��q)���qH�R�!�!��A:H^/@��X�������?�^���y��������}�~8�f 7B������r29�����<Y�<Y�<
9yr�9�	�㐓�'!ysȲ�9���\	�����9����AH�p9H����}��q�g.�ˀyM2�`��?<f���z�~��>��ޏ�"|#�_�p?�ǀ�I��&��gq�6Iy�I���,y+!7B����5�r�,Bo�9��-Ҿ<�~��d
r�rdr#d r%���9��
�A�l�r�8���sf�{rME���R���qO�Sh����S���'��z�'�&Z&f�rgO����=)���o����e����z�~���<�q�w�HQt����N��Lz
�|����1I�&�E�����?yO�����O��ǟbS�)�񥊞	��!M�f
�s��KI�z��1���m�}^��[l��s-���1���+?מ�z߸�_�&���@�O�j�����2ReP��������+4�=�3�Φ��	7F=���������ZR�LxTsd~��������6Ur��?;;cƖ@�����oo]���o�~	�ϟ����z�չXX���X��}X�}X�{�
�mܠ�p�<�#�:׹X��X����y� �:��X����::�΃����y��U~�'��9��M��80&����J�����;XN��8��?�x�����������&�7�ǁ��J�p �+�)�o
����?f��T_8��>��-�%. �>|px.�3��K�����ώ���?����K�G�������p����W��]���}�_V����_��[y�h+�ߌ����5-��[g�=-��Ɇ�Z*�;�RY�}6|oKeyn�,�[*�����w�i�,��������~ ��v�ĞO ~p7����/"�"��xxpzv �� ��HQ�1����
��}J?��Ok���Ee�����x��E�?�OUz<�+e�u��D�`<�<����x<(�x|����)�(�/8��!ڂ�<_ ������+*?8�Y� =n�]�K�c��Ń,O��x1���%nk��xa+�/��
��p
��'�>8��S�x��x �8�p�x�!�ߪ�~����
~��"�9�$��%^�� .B�!��A��?�����7�{��� �=� �;�W|<��y�%~؇>u6��P�M��}��'��C�c��_T�������o	��/�@��S�J� ��V�����W��G���I�s����p �a���x/*|V�?$�K�~��<���r� �	O⁷�xV�O ��`�׀�wH|B�{���{Q^��u��_J��һ�'��}��ў?�ßN=����9<`q=p 8�> 4%��7-�S���?T�3kg����^L^<};��/r�A��G���_U|��F{����c;p��b��0�� �7��[�"���9�/�>� �Kx�?�C�p?<1<���G� ~H��H ��������+>�˓�����$p�G%^x�?�\8$q\�%~XC��*p���>��S�����핸x��v���c��wK�,���/��s�<��K;��{�>���$. ����wTz<��'� �+ބ�xA`+��#*��I�׾�!���^`߹(��8����p
���a��;�s���M�:��sW�'��s[�C~X� ��b�<���;�S����X �b=�a�"��~�*��2�8�7�}��{�X_�P�����9e>�Ǖ��xQ�7�P�k��x@r���<~�ķ�x�ϫ��O���Q�^��*p�g?\����+��?R������ʞ�x���,�"�\�I��*� �#�Z�G���^<@}�JT�]*�=J�?K�x��%~�ҏ�}@�?��?�������q�����#�'J?���%�[/��S��?(�x�6 {�#qp�$��~	`?ؿx�X�yN��Q��}R�a��=c�F�o+�0��� �Y"=������ OB��G�&��oK|��e��*�?H����;���>T�'%���s>��q��E��SJ��V��/({P��(��4��ON!�\� ��E�+�ǁ;���[�s�J�Cy������'�Q�_��Q��'��K��E��i����Z�ޟ�>�ǰ��x?X�
8 |�҇�x�'����C����C���� .���'�=?���4�OF=� <�xxx�E?<��/>���T<�u�c�7� ��8<����?<2(�׀s�ǁ�ϽX��п �$����~`��<���ۀo��<���V�?<�"�������Q>�E�c�k��|� >�n����~��|X�.�I�
�n��|��*������C��){��+{����������p+�O�ې��R��9�^e/�I��&�V���)�O
8�.���~�� �s��)�����ߗ�7?���� �ρ��͋���M���g)p x=�J��TP���J?���A�ǁ�(�S�G���	�����w���Ն�|��{3�Fી�A�&����"�.���w������? >
���x����+������y��ƴg<���"ď�>޲��O����x�8<�g���<�
�<��������w�������J�z��͘�?8|5p 翽��G��8_4����XCy������>���T<�Ϗ){P?���~�p���*�S/��/H|>��=��cx9��ZŇ}������a��8��}p?|� ��`/֧���K?y���߂�Ҟ����(�ry%�c×���*n���pȆ�a��l�6��Ά�n��%��_��K*����96|�/��6|��Ն7�p�o��m8f�I�k�w��_����T�σ6�9�?������6�;>si%���R�"[�2^e��m�ǆ����6���ԗ=�GI�@r�H��HO�<���_!9�#�Ҥ��@�y#���)�I���C��L���8}쑿{�S����?��/��K��J�_������G>��[��������$������}:~���M��?OE�V��J�YM���N����=��^~��I>����&o@���ߤ�'�m���_l�i��D4��dB�d4�鉔nj����e��P�0vgS��z8�o�վ>aDv�Ŀ��c��-��#��12�'�♡�=�v������L8�W�����	RQ3̽a3�EZ#�L�H��!#�L�3YS�4�^=�G2�i#�z:e$��>�BXj�*����P�r�3����z�5���{��B���#Q%�}(lV	�2�)�)�+Y-�۠6�\#�3a��i�0��j��x2�W55cf#St%��*��Ne3����o�5��05]�c�%���� Ud2OS��9)_���Qq-���2ɮ_ƸHY��h%LW���(��M��� Wt|8��2{��UW�rE(�ȦCA,ĥ�Z�uTOG�x��&�N��q��p"4�0�	�s��B��É�^B�����޷#��&w#86u�pCi�0���*�/���Q*%�c-2GdӺg��N�2� ��o]��!##�դ�lJ9���T�Z%do<I�Q�N���b�|���Y�H;,�"r
�7F�{�᤼��⢝{���n*.d���+��$Kt�}���'����|���h�c�7�|UCC����Ʈ��"dS4�eh$�A����h�ѓ��g�:i�}�pJvI�C�VZ]�gh8r�B�:����xBu�pmO�a��6�t��$��p����>����a�r��2�ji��Y�v�$�6TIZ%ʚ��*����L6��iP����A؀���'�4�+����l(��&:�A�pG�N�q��<(�c*�N�݈GU�'K���~'�ͽ��4KO�x���1�zx�3/F��;:<`$����3l���������k5#J�^.��7�`��S�j[&:�/KW[M�G���;ٴ8Xa��R��:��nH��4��T̃�+"O��q�����X�:I4J�DW��p*�g�� s����1�W���+%4���mھ�V��a͚�r��+fh�����B�ìЁ'N�uUD���)֕
�B�iMk�Q�ԣ��aF��q��kam:9����b�1���V�4�uG�'�Ⱥ֕9�3tGL�e�Sl]�,$�y�c��Z�1��}V�4��K��:͌�x�QnX�`8D�d�&X	b�\��G���3ś�Q��e�(��E�NWo:&{��*��jQI}/�DW�X��`#B�U���ĢZ���4iuN�W��jE��U�n� �����v5߃�n��崝�7m�]N�i�i;�f�N;N�i7Ӷ�Tw�I����u��i{*m:9��֞�Ӯ��)�id�Zk�N����Ӝ��n��㴝v3m�I��tǬ=m�]M�SX�ȶ>5c&����H�ZT7�dL�0�V��Վ5��p&f��������p*�!q���Vq�R"��Q;��$��j��V*cF�1�p�Qv�!f���{�P5�i슄��|�S��w{���ܦwk�z��*�����Z~Mh���<=�^>�B[�oj�w���-��@x��u[��Kw�˷��ټ�o]��[�t�0uqw�W�}f8Uے��h��d&.q$-��%.ձ� 8���hZ\Y�xZ^�jq�#�m��Ȇ��.:@��3����t�����dT�-��i�����^M�]�'u3�t>S����W3K�U���
��N���"�4Q�;ĥ��KY��Rգ �Gq��Vɻj�K,��@�dy�cJؖ4�������ke_��a�Y�P�1�i�a�1�ڊ-�1,�'@�>F��o��.�%@�HA���b���Ԅ���u�x҂;Ź�������Ƅl���hd���u]Q��@݉����a�.NQ����⎜S�T�U;�hD��2^ٖ�:�z"Z��'��@ق�6ݮG։�d��:@kg�H�����,n<`��
G�z�@ٕ,�<`s�Jo��3�m֬�Yn�j�fW���D݆�Ǹ@m��F����X�m*8@�m�X=�7����+V2����qH��9�U��,��d=�&����h�xi�L+A9�K�%[E\˓��58�6/b�ݍ�����+O�e4c�uu*ףA��$��&�g��]�hLv+�]q*-O�	c�i��|���v��+�L�����)�M�
�$әJ"@e�r�5z[J�"��Ł��-O�+�2�:C��>�/l��o4�3�z@I3]��V!V��N����*5U*��YT�ѥ+�n�G�}C�t�����8L�n$��K���[z6��GaveR)B,s-x�F�N�8�n&�i�V��˾k���ޖ��L8�X�vU�~Ep����K�[
�d�=��ĩ�F���F�JQ��Җ�I9<63i^�r[Y#,7K�^@UճG�2�JF����}ar�-򱎐�K�bP�Y� �cQ7��.g���ikE����Q��mE����p�94�(c�rJ��Pq�i�TG*i�1(�ekKd�4&�A�3u̩6���w%c�J��[~��4�T*����������@)e9�J���ݬ��k>�&Yt��MA��o��׼�R�5�L�-#��$KUӻ��T��WϔZ������`PY�� K�˝QE3[��n�¥�L�E��A)Ȓ����DT&*Y%���X��'�c�e�V��iag�D@��ԥmZ�`���k��"K�o#O�ڙbu�7b{��+�\�09�VƔ��a�떆rK�	$�%�ʪ΃
ؓ���σ�?]�厞o�ꉘZ�1��hl޸~l�����-b%���+=����	g�6��L���eIԛÑ���.�Z��p8N+G�ڎ�=}D<�8OS9������qˬ�{)�-!&����������^bO<ME0�����^u�c�)E9*$�ލ|{ V��em��6(Fg !3��gJ�B������<�4��PL<hf�Ҹ'���,%/Ͳ.�2�ыs������O&�Ó��d����<>�jϐ�pdH�ړ	�}T"L�f�����M)>P�&h2��v��=��c��T�����{p�V��]��ͩq�;g�6��p���I!�i�i^����7���+B��H��SaʢTFx5�N:�G�1^c����(P�a�
b�o��DɷeO �(`:>��sC���)*+dj��Y��W��y��j��PK
    +Q�H`4�].�  �� %  org/bridj/lib/linux_armhf/libbridj.so  ��     .�      �}\U��?>QI��FFyT**�c�RQ��S�abYY��B!�Rѽ�XT��hv���ެk�-+�jQYyov��������PTjT���{f6{8?������Mk��Yk�Z3{�>�8��p�/PD	�6�"0���[�p�nȋ����K��!C7FJ�̗i�P���`!�u>���O�X�6����6#D�`�M��?f�09!&L�&�����K^�汃��vwkրk���D>�p e��F!<��JC�ա��8�mN���"ܠ'b�>��G�cLP��BX��T�8����x�.����M�~�+8�Cu��fi<ژ����~��KFx�J�IHx=�a!�#�	0a?�D�W"T_�P��E��~/�=u��n0hhEx��M�i���4�n�����/��T�;�����!�~��r�/�xO� �8�x,`����؁�ˏ@Hr(y���Ep��!�H�!a8�,�� ���� 
�,��t;� ����!��;�Pn��� ��A�W ���Ql���\#\�0�c5�{P�9�����X���#�q�w�>D�G���t;��!\����'��?��6k�ġtCB�!���Eǿ@��+��Ju�4�G!�|ੀ��t~Ҋ5~�xĩ�n^�0�ψ�Q��!?�f�_/�4L���_��Ӏ'�� �8T��0�-q�41���)s5¿���_���p����YC���:fp=�x#�2_��0�/���B�����"� ~�x����_R&!$ �B�~F�!���2�}a�t����E? ��g��NAXb�[�0ӧ� ���x,�.�'n>J�j�����lߠ�Y�����2���y��Ku(;d�-5�}��H�p�>]�� ?�������.l�=���N<�ȫ@���^_���~��a�N?W����׍�'#�4�J��B���I�g��CK�r�#,��s#������e{h|�1h�a�n�:����x�H]��鲷ix�A_	=��@��a�W#�7��7��gnF�x�g�#���u�Oݟ���-���΍����R����i�_԰IC�Xh|��!�����p6`w#=ԧ\9B"�LFx�H_�p�w4~맿���'�?����~����0a����^���
��N�a>�e:�
y�'�=�?����.m8��x������1c*�SK�C?I]��2~T����ԇ����W��!��\�B����<u�Y�ό�Q7q���Qxi�_���1� ���]8!/�&�� W@ȹ�~��Ʈ��yvOWvIB}OIxI��vA��*_�s��[N{�1%��{N�Y�_�&�q,y��I�KJ\�""*>A��<�4X�黸��yO.^(J����yq����Sr���ߦibM|�C�N��y�c�p��=9<���3���O��������G��[v������Jz_��-n�}MK������������_i,�H�<Θ��5�B�-�I�G7N�mޕ_)�Wq�F�Oh�^�SSoЏ溴|�(�����-�?A������!�S��4�1�k�>��(Ô}�E��-ٱ|`���=��h��'m,m}��5��}X�~��t�<u���:��M�sig�sR/��+qC�B��~�����}�^�k韛k�k�ӷ����w���^�����hg����H�{P�S�&S_[v������+��t����G�Aߋ:��/�%�!�;P�p��}��|��I�?��rD;�־m�-kG߉���u�>�4}���}ە��4���q�T�}��ץ/�=��Υ�r���n�����o5�eG�w�^��f��������E?�{S���sr�}���
���*��0������g�4/_���r�?ʖ�r����4X���w�y+i��v�Y[�9�×�����Y��&2��+۳�����_7~4�����}*#�>�?���?J�Q5��?�����Q��}�rY��L�勞�eYӫ�m_\�3�1i�go���#�3g}԰;���}|c�CY}��'ya�+o:����'={ٺ���������e���xw~~���<Qq�lZV���n�o~�vY����?������m;�¬Wo}�Ao=�$$�v��{f�x���ě_�3`��^���O�[n�����E����=����K��eD�M�V�x~Щ/?s�ɕ�o��u�G����3S����த��Y�e�U7^tI�揧����/\���w�7lC⢁��s��S��m�>�������)��kB��~ ll��1���y���Z��l�w�i��Q��W���`ص��~��?���w{M���;��\��	O{`���/UO��f�y��}bȨ���^[[V\vϘq��~��}���7:w�|N����ߤ�Z~g߹�=�A�2���u�E��7f\���ٳ��>��/V����C?+�h�{W�z�o?��E��>gڮ/�q��o��ׅ&uo;��K��;glU�����R}���^tઑ�9�֝:�Nׂ个�����ykd���{z��3gʠ�c
wݞ[�V�ؼl�k[W��~����u���?�]��y7��²�JS'4~���㊫k�<�|��A�����[X�|��򆖼�ї~~�ŉ�����v̛6�[�BLk�̌�b�.|���}��[>���I,���2��z�rcj����z�m
|��ˣ���i����0�|m���/j����GΞִ䲝	���|D[��9�_��[��7o�g��w�==�$��a7]��Q�<?����o|����}�����ޟ.}���Kyj�G���\Y��޿+��~��ߍ������<%�׍�<�F�e[^�p|�o\^�Zŏ��yoB��>=������d�<0p������7��~V�pm�i�=Z���������K�׌|o����Q[2!i����[p��Q=����^u���M7�s�����碤7��u7M��g��1�/lw��Lcn�#5~���=�s�]�뤇'�'�}Ũ��f|s������~�`C�}}N����ۧG��[�i/�rFC����{m�����_���8�ۏZ���<<zmҁ>+Zw��K���O�aH�3[�Q�Ӳe�?=���O�p��S2˂��������_m���?"��X�,k�'	����r�JG��V�)�����~x1�o�k.��~��}����?��퍿>�?bQ�G-Au�N�õ#�����=��˟.|�R�s�{um⾖{G�4�����Nz�������#��=�̢�)�ur�=�.�j�y�����+#����/
��ꪌ����u�긟�KRR8�շ�<g������n����zt�O�_�Ƀ�C����m���~`N����������?���ٴd����9_��?o������~�}YN��?u_�ޓ��;`>��##g_x�_��^���97:�V�\�8WL��ᬵO�9�ˑ3'�*_�/��aJ���_��1cn����|�ޑ�W슮|4n�]IQ?�^19�ʿ.�j�i����u����퍮��5�]�p�?�^z۟�R,���OQ0P�x��ء���y'��x>��������<;9ӧ�@;*ϒb|�/��.:�����'��'~v�O{���������|�9�G�x�O��gW���O��}���_�9>�g<��Lo���v�o�鯻O�7�����s���v���v��:6�:��˧���X��{��n���۪΃�?�3ƫ@��@��3N���Oꜛ�;!�[�;�9B_HϪJ�����WA��3r���fo�Q~4�Up�����/i���I8�!�/���!�;?�sȽ�o�f;Ө�g��վ����Q����ho�Q~kd�s�}�/��O-�3�Ǣ�ˈ�ўˠ/	HT�:Gb� ��n��s��Y�'b�f{�Y.�b��q���߆�c��*�|%?����W ��!����7��O��=zCz���8�q�|�K��!�y	������G�plβU�k�G�=y(3���=����� o�>R��ǣ��(7�y6�|����A�$ k���,ꃱ�b�����C��OG���|L�"��@��0�A�1F��N}�r����o7��n�;��0�����_�5X��/������(Ԩ_��������U{��3�>�Yz\��bދ��W���}j�'�������p�Q����
�/5�C}|����[���};�����!��F��Bv�;:�ť��dȫ%߂ު"� 򸩗C�_��k�c���P�'��ǯ���������������"G�<�7��[k�o�|���{�{Qt��d�����4���O�g��=���P>��7�÷<��H�?�c��:�A�K���������ۍ���a~k�|��,��_0��_�����!����T���2�!�92y�>�!�t��G�����/�h�㳞~B���������ly~F�o���Oo9:�s*�U���3�/�ǻ�I�;�e��ǋ�Y������M����u.#��P�h��`��"my���������Vлn�:�g|<�k�0��6�w*���!��|u���!�[�O₴=D�[�m���Y�\t�w.��j��=0�C?_F{$:��ר����f�����^�6���o��~>�=i�%:�?���!�Ť����)���0(�U�=�|�_`�ׇ���V�?���5�߃���萿(����X�_D�=�����ՙ��K����A~,}��+��,�{c}l6�{�G�C��ϕ��+�O�۶�g�^�_�]�<����R��u���
�ﺏm��y���]��A|6k�w��ǰ�|��\��B�O�&-RϬ�FE��w����U=b�!�ذ̎?KF��@����B{ی�����O��DG�>�w51����Q�~�r�z��^� ��E�<Uc���7���m��~E]jۧO}����Z�D�>;�����R�@^k���+�>c�-ϛ�^�ϴ��s�C�� yp��<����ǀ�c�b�^a���nC����~��|���d.��־��u2�y}l�p���ϥZ_�y�a�ש�߼����a>�~���`��0GG<�3��c}�����ٿ���4�c�;����o. �¾�����({}4c=��Tg���`�z�OjB�������	��j��|������(~^ݭ���}���~�$q#�I6��*}E�{a�ϴ�ު��0��>��/�ۋ�j�� F�U�ی���%]l뇵o�uV�x1	Zo��O�����=������2������f�����Ч�C��?���a��n����F���^��d�����m�~.	�����Xc������,�1�}�-��b�%�a��?Ag�v{�1>�G�����v�=��p?1����z6о<o��q=���t��_d�^l�2���@��d�/����[ �̜g���ۡ/�u������l�����J{=O�?��d��k�>B=�9�\_,��.��krl�%�}e�_����݌�E���'������!U_��r��g\��O���b{���s�O����;���h�?{%�|����c/#�q�zV%�����{�;�E[>� �/�y�@�UF�[��j~���O�������_���y��V�'��Hs�8t~#�{�+6?�Q~�˖�8�L(C�?��_�!�~�����ي�[!�z���;a#d��ϒ�([�tG����=8�!}�u��?�[e��r�#��/_���^���}j��|=�����|�����h��mF��#�X˱>�M��o�?@~��3��y�5`\��� $�(�#�g�|c���(�f�?�1?�o�f����6�WѱY�������Ǡ7��o�3�;�&9��7������~����_����
�a����^�(�Vt��7@�A���^��X�qa�C��V�������-G=Gd����NG{����g�A�k��D#��%F|�G���? [�5�j7��Q�O^n���b|aF{O`>ۍ���盰?���N�_l�� �H4���1�5F�(ʛi/P���_������F~.��4�S�^�s�x�">��k(/�v{�З%Q��l��/_�xÍ��q���}�%�?Π�w
��	�B���_�ܶ�����z^{^~@t��y�m�O��b�V{�<��v��c?��'̰�����w���z}z��o���ps��7�b���/k_���(�f����0_���7��_7��O�Ç��τ�}p�m�.�>�ɱ� �]�d��H^����r�í��Ø�A�����l��ɐ��nvP>�(O;\i��{@>2_��w��W��v�<�
{�x{�z��o��2gnnNJAaZ~aJ�H������YEiDӲ���)W�O�6cNVAaF��촂��169�ʴ�icӲ�'��gg�L�7S�Ϻ:7=`t���ܬ��Pf���Y�Y�922!#'#?kVGZ���F������fe���#;2
������LN�O˛�5D�����[�扼|4:�0m�mȝ�!feg����3�]�QP���aՔݫȸ���|1')?�0cVaF�����s2
�|��[Qp|n��¬�ֈ�U�'��Ӓ��ڲ�8�4f���r��e������e_�Q���>>?wnrfV���)Ϸ�ٹ�ٹ�����q*Z%%�o��ْ��i�j~SR2��srS�sg�I��uvFL�%�t$Hi���
�8%7N�����[S:2RP*!�`V~�������9�����/��du��E+*������S��1W�����y�
Evn�
�P�:�є)�,=���B�"
�椩u0	mia���d�HQ�j��S�'�`�^z�0�����oRN��[D��g��$��Ą�y3�3��1����``��*ylfZ>���Qh�����/[U�w|vڜ�Ҳ��V�B�$+�����Vh�#���k��2����dD�54-g��DT))�)�Ӳ�I�.��aUP�����em����%�t�#���B�A%g�2Gv�D&u˝�(W� fw��P���˹�k.0��)F�p0�#�y�\��8G���[ىX���f��1�����2rҕ~�h� St[��T'����
3�)�i�$nI_��(�Ɇя�:cFe)���ؤc��Q5��i\f1v"�P�g�����Sl�R|�lKK�iV�d�O);�J���S�N�R0v�2VJ��<��#Z���KQG���i�)ԑ�����j�F�]I1�����d%H���Ӭ�M�bF�N���u:yR�59��i(r�uW��y�`����������rr�l�r��e���r���	����3;�5F���5@�x3vC��2��W�ţ�
�&����e����M�X�R&���ˁSdR��њL��"Q)
�h�����t�W���$���r+�"�a��;9}��Ă;���͞�6�Hˑ���N�+��\p�%V�����񩛗��6�@Ny�yFN~���ȱ3f��/H�O�H��JG�|�(M�I�(:"5�<�f�lj�N��a�:R�,�/�0v%#1=+?cV�YhlR��3>pa�,c���P�J/�#}�䌌��1B����A����͙W��
����BL�\�?�$)tR�5��ip}�5�B
k�&�"e��K#D�!W_b�̤��LiW2�gO��"ҳ!3��w��2���rz6=��O˿14Q0Ie�;/�¥d�K�_ ��=�l��r�|;�j���)�s�o���g�N�U�_vNƂ	ٹ3�E����T�q�"h����ۺ��q�q/7l϶<4�h�G:6v��� %v̼ٳQC)�.����6+��E�;q3��>��f�gd����c��$�/�F��(�����I�j�=[�����|�Z�r��u�E������^iL����t�d�~��_%9G��\s�&��VjV�T�������ϝ;Wm`hF��z��)����ZG���s��n;���Ghoέ������ѳ��}�EB�Pl&8fl�Y��ʰG��Z�Q��h�����I7M{tzZ�2�������\�h�j�A��]�V̲	Gi�.rB-w:�8j�J������Y��egg�/t6���-�*��<$���X���u�*8J䷗�����j6��͝�J�~�9s��9�Э9JGG�d;'e8�1�5��R�ä�O�*ȅ���V9��م����2<-??��l��O+���Ċ�u��F��쌹��ʲ޸v����\]�<�0����.�ǂ��m�KL8��4�(�U6t�������.͒,yԱt!����+tDK]bǉT��Żʐ��t����h<ZfG��M�q�p�]V��J�fe��wI X��7��]o��SƷ�.	�	����*�TVɈ>E;�|=߬\1;n1J�*�ea�bqI�l�uIdɣ��]��x�v�BG��%�;�
�	�w�']+,�N���]�,U���R�	tt<��ԑmu�1'T��[Y����B�c���;3���2�y?�\a��.�[�T����g͞ݕ��|��B���ӊ����iyyY���I���qt���d^(�v�F����k6N�w�g�y�2�r[�z�/�$g\�qGG()�˘�5;kVGZ��&���ٯ�rBZa��Κ�k�_�{�[=�������m:�xT�>���>�F��%��3��sSfB>�Y��2f��n�ԭ����q!��9[�/�Hzv.
���-�s�剹�rҳ�������f?���'J�z�(#F�i�S�����h�q��n�$g�˱�ǲ����)�i�<RE1�
2��$�ea��Y��|`_PU����씔����y�E�0_א�7!qҘ�)�o}lF����Z��)�#G��z*O�
������������9D���;jaYY'q���3���*_t�t�����"7]���,Ӱ\�J�4\�a��5�j�Fõ�i�NC�C��!��"�pߥ�w'a;�%�.D8a�CD>�����$��Q�3��&��!܄�B�9D�,�q�"��j!Ov����	�Hx�I����^��	K��A����B�v�L�MX�y�7QHx�C&;D1a�%��;D���Mx+��|�7a�CTN�|���&<�!j��|�;��ØoB��:����!��q���:��'�W�M�����!�����J�Y�m�OBl'�;�<8��0�!�	s���<!��v����k�h'L� !?69�A���?����
x'�O8�!������� ��'|�'��^�ф#�p.s����?�:!�/�e�� �BL$Ls�D�=�?��?�x��'�(D*��H�q�0�'�T�<­�?�T��]!�	���7��������4ܬ��j�M����У�Ob`�#�	�$���nao�'!�M@�M�"�y�O��(!��$\�e�8D9a0䓰���.�|b�V�}@x�C�^�$�$��u�1�O�ȧ��A�����'��I�w�	{A>	�@>	�|�
����Ax�̈́�!��� ���
�FM��p�SΛC$�#�~�$��Ix�C��}J����*�'a�'��O�A)Ӆ�"��|�B>	O�|VK�0��3!�	��U�O�^�OB(�$¾|��7�8�'���?a5�Ox���#!��S��<�($��	�C>	�|�{@������>�&����;�*B�j¿�������= <�'��#|�����?!���	w����`=���@��_��M�7��r���ǅ�΀~��
��ys�=��������t�h���	���O������D��'仅����+���t���?���?�$�'��|��
���;�0�'<��p8�O����'��I���Ʉ���	����o����������|O�0�'���w��,��r��m�?��X��X��/����a�s��	ǂ����X��i�?a&�O��0�'����g��r��9?�?a$�?�j��+�����0�'��?�#�?�����C���O8��� ~ǟ�]`��R��5�s�7ȳ��۳�������}oI���.o,�y���<���|��'x��'x���x��Gx���x�����l|���1�f�i��|��o2�����x��Wx���x��x��gx���0�dO4��3��6�H�0�05� ?��1�����|��o3�-���7�:_k�^m�U^n�^l���m��>���<��<��c<��#<���<����`�1�����|��o3�-���7�:_k�^m�U^n�^l���m��>���<��<��c<��#<���<���4>������o6������&�`��|���x��Wx���x��x����O6�DO0�8�1�h�4�3�P2�����7�=�l�;|��o1�M�����Z�5�j�2�r/5�b/4�lO7��l���`�q��_M��/hs����V{�K<���Me�����]y��gb�5��\K<�(/\��B\�"܍|�n�=#Q&P�nx����WM�,�z�K����x����"_���!UB,�D�>*�>B>���>�Qwފ�@g�;�kB�^�(�j���&�ɫiH�i(:|x��]�ep�z��?�q��
��Y�mӸ�^���ɲp��h[�A��U�n��Wx��5��5M����� ���~B�V4���r��eYN�/�Z��꫽��%���Çw�̩���;���A���\���ol����.~�ڍ1Fc|��
o������`�Ǽ�Ί�Q�q=�%oB{�CV{#�c^�Ή���s/�:C�%�6�ʽ�E�?�����>%��n$�t�E���}�G�l7����B�0��u�=����=�S��ض�&�Y�HS �}ǹ�{�?�Ԉ-vO3/^煠m�Y3� ^sH�1H|�Ɯ�1�L'�/��o1o�7�~�c��ޝ�"�2o�˽m�6LD��P�2S�+㷷FCf +!���#ef�!��
9�Y(yS%yBތ��z�����f��@=Q�U�7J��� �z���+�����W�=%K����*�#��gck�6���������w��B�����k����������5������:# <�,��N�Ro ���εF��%_�#�|r�O����<<�->9���|"�N�4��?��
�殖�	E�0���"o��7ԫ�.�fac�xR�Z�Y��y��C4�̇<բ�T�ZOUw�-���φ�j��!�.������99��T�h˰�8�s\���:: ���uQ7b^ ��� ���˽��T����T� `y���j��>���R�)��u������$��(�5��{��i�:m6�������h�
����M�\H�P�1@^ܕ�ג*ohj���uE����/p^�{%�pj��A_�~���I��.��
o����,uD^R����^��"=��%�'�� O�%��0-2���DZ�4�)�*�ߣ��"��$Ȅ�o��֞(WrP��(��/(��~�;����6��8���v{�]7ڵ�C����C�?齑��Z��!{��ӎ�V�9�?_+W��y�8��r^��@�V���Z��]��M3;�#�#��"ڠ}{��{�;tk;�Z�=]ڝ��P)sU�7Ю�ǮPg�v%�ۮ8��4жk��ϛ1��i>ؙ7���u�<���y���7K���L�&*����)\7n��O�6'��Y_!��`��#�!Č&�G ��3ȩuT�g�7	s.ܕ��e-�]�ZB=u�k�Wx*��Ӡ�������!���o���a�*��m+[Agx�C�	���Mk�v&h �A�Rٗ���w���t9Ǘ�}�����BG�'.{:�T�:n��Rk�h�O�s1���L��ߧ/|�A],S}���W>���bL���C �����J0�%���EIc�Oy��u-��~���J��mU�X�u`m���:Å��,�m�b��F���L��8��6�d>my�9ސ�����%�v�^�E��-�O�����T�'P���X �A�ثԯ���Zb�?(�� ��?���x���O7��=�Æ����q܃Y>�-�Z<���!
 ���ٶ�sPi����7�h,IZ�]�y*F�ݒ�x��rߵ�%H��^��P�-K��ơ��]���5V��_P
��)Fǳ[�_@t4E����e��(�+�|����,9t*�����t�+w�J���A�����w �Y:�~�!�����޿S�j����Ҝ�����^���S�N��J��k�� ��������)(����?�����a�^��֑ԃq�s�Q��z�Ұ�����g�"��á#�+c07�ѝX�a(��q��@9��8�R�G����TtґC��0�򯅸�i�ԍ�N?�}1Hk��q��Ǉ�ޜk�7���kQ&L�1E�_�/���.�,��F�w*ڜԏy�~��ϢƔ�T�{��O�t�DR�#?�����ޏ����N�Q�*��T�X�Ֆ_U��B�Sh#�^��[��񅺿h�ҹ�1P,m[�F���^n��&����Jo����"����3�N҅jM�QrM�L����L��S5�I�0�I��;�?/����p��=��	�����!v�A�a6����i�&!�F�G��F8a��ف]#LG������/�4��<P��-�T}9�q뵞��+m��G��F�W�ְ��W<�e�7~��Te�'Y�!��{�h��7���#��gY���ߕ��~ =;0�L���'K�o���H7�u�ͯ�ql��#P>��·�{�W���Λ��=�l]����W;/����u��9�k{��l��_�����5:~���7��'��~��|�=�KA���B�x�i�:BשB���砫׾��eС}�@��k4?\O���=k �%�=�~q���(2v���~'#T#T !���5a�4����AG�:��+!�?���h_�Q�Q)�aΙ����1���:�p�E���,���r��F��C�,�2s��m��>��@�!z&��&�C����e�_���s���g�^�_�'�h{ m�n;D�&V�+t��X6ȵ�1ĵػ�h'�W�N����a�����u���~ʷ��^4ҟ���{���f���H�]�ס��'Qs+u��t��$5]L��D��r�	;^���Ɵ�ޭ>?G��)�5p�����W��9�y�ߋz���Ӿՠ��v{m�|�m=��ۍyz�({�A�T���n����"B)BҶ���w���By���uy�W�[�		�})}�}C׮��^�?��6��P�G�<"*e�*�}a+X��a�����p�X������:�B�D�A(D���w�Cؓ�J�?C�����ԣ���*�o�\;�����d�Ր�����~��������'��wg�x�54���m���Q�ʶ��=�����w��e���T�)�W�f��ۋŭ_�׳����] �,���6���!��d�9�]�i�g��͏}��F���6k�6�����O�y��:k�:]�-�/T�Qe�Ļ�0�n�����Ǒ����W='m��0�2��n��xo%򪍼�t=�s������ȋ2�N�<�χ,�f�%D��!��lY�)�_̳T�{w�V�`�\�U��.0]��D��F���P���{�Pn�Q�*��ɿ�宧.3�E���҇�~�_첉Ҟ����G�{���&����e�"�r~�%���Ɠj(�Z��yQ~��yC��qR�ZV�A~�>�y���]��B��Ytv�V�j?2��彩�{��󰯤��}$}�@���+�g{ܣ,'.ϧ�oy�v;I��y��O�����D�9�>"�8�d�H�*�ٴ���i��!"�{%�=~/�KGB'��Y-�!��H%U�!�y���q �k��g@c�+ >:�;(�~���|H�0K�ChA��������5�z�yO ��u�]�c��E�ep��7l�����:m1�e���|��.�gRa���#������\	�e<��Sw�|���ޭ�����m����_w�|�2�w�Αg�*��סo��g^R�A�o:�H���Ƕ~�ZӅr�i�H���O@��}����7�c�I�u��9�ʄ�����c�g<���0_�縉'yF�s$iVzO�Ct� ��)��R�?��{����(�yh�9y�>�����)S��S����-c������D�J�K��5Њ<s\�c\ɺ�u��Jo'}�w@�5V��?���@}6�����K��v=��H?Hѵ���"m� �9u�J9�������A��t����1|�AF��>��4��y��ܢI׽��<S��q2�W}ڈC[�6X�}=����E�S�{���F�L-�x�l����ߌ��"B�m'�0�yj^Iˏ��3T���y0�aKd;�%=?H���p��Q���������ܾŷ?��#�tn�>��
�>��32��k���s���������C��J>C�{ķ;~��}ڽ��C���N�S�?h'���΋h��hgbڙ�3�.�K$/�Vv�K@7��}���<��vФu�m�Y:HɺZ{�mo��b�?	���O;����E����ȧ�T�7"��t����4���"{�9�w:�a+ڍ����2��~�(ǹ��~����-�e
�,�o����KS�_�_�-u�=��G;e]h�/x�ޅr�|�[a��0�����>#�T�#(�ƙ��=����G~����<����F����������M;�]���t7�ڏ�NB;EF�-���Iv�m|����6��V��g�0i���%�޻nY�2�M��zY=[��P�Roh�Ro$l��ߦZ�[�<�u6��;�=��z��gN�o[wX�����.�i��<mF`��T��g���6��I�k�|V�1�]�‿ʱv������=�}�����������7�����M�����x��-�����k0Ou�ۥ�w	���Z� ������hc�p�o`<|������@�܍��"�=5Q_�6��luW�g��9�!v�|,h`ߤ�Ϧ�|f�ᳶꖠx�w������ʻy����F;�?��վQ���8�ut4l�!��4T�U�~l�!u��y�v��6���8D{���=��o;��i��Jg8�+Z�?��z������G��~xp{��#���I�1h��~�C�C�А`���HC�������ό@��з[��ؿ���Uh�:��tT���:�]��p��E�ԫk�A�Z:��"u�P6I���}8���O�����=�$�d�2��i�S�ćҎ�ާ�h�9b)ڧ���kՅ~\>4�4hr�ߓ���p���zM٣誖t��E��\���(��t��t���t���6�?�m�zv_��}.�w��'���L�!%K<���3�T��U�.�֫;ֳ�x�U�˽��W˻"��<e���iMlc�<_��~C���A��M���I��n~�cZ�<�6��������5��v�o��D[������ϰ��}�2�Fݖ<OJ������6���EcO��q��Ht���;~������X{e�y��
���9����#�"y�{�7D������`[��MkiyzM��3����F��3)��Z�"�aʵ���3j�g�8CHj��ȳK��}7'ϹTY��G���.T_���΢~�3��֪�w�5W�V�i� ���+Z�ދ��%B�%��9D2O�!&"�!��\�r/L�o}��]�5�'�ݮ]��}����~D����(���u���&o�m\X�@�W�����O+������a�O+߰�oB�A������-uS>c`%uw�ߔ�O���%�c�϶������*s;��:n�_�n\�W�w� �!P�����Q�U~i��k=�JO��7��Ɠ�Z�V,�oxM�Uw����`�lx9��)���lEh��a�N߃��J;uz�.�ߕ[
X	XB�X�P<0��XG_�wf�]O��3��D���3����eJ��q��7=!D�n#���'O~J��Z6�G��L�?�X���pl��B�+Ǒ�C�蹈|J��{$�X�v"�w5��^<:H�����3��6P�������9�u����[��tͫ�[�f+�}�g3������`oX�������UP�&�)���`u����(�ō�C�8]��%BQo"��]N�qēO.Pexǥ{��X$�9����K�~L��헢m�+��+�]����WK��yG��%ʼ�3a�+�Ww%v���(O=�_�"��s�)��Yv�[�^E�`����
-�1]�%m'�t��"�+:AZjO��-h{KiiC���%��ވ3P���wشcД0`�7᢮є�r�N�����>?���.��A9�	�:��L5?Α]������1#�F�t��>��h*E�RMSYiZ�>�v���(��i:�:5MbT�h�<y�7rT�h��rO>1�
Q��,ESQi�F�]����O��=��G���E���ab�FS,�ņ�M験�hʌ�M�裼�4ա\ݱh��Lm�N��i�	�gs�����ԫ��z�ubQ'�5~U��u�Q'�u�:�u�Sٹ���+Q��u�:��������Q�k�Y��|��#q�|[�iF~3��_�����w�3��#��.�%��sX���|�Oy��n�u˲�d��KLZ��j���Y���G�_���F{��io�W����5�)��d��e�MG)o��A�G���s�1w���۹���9�RUN�k��1����$	�I��<�~���:E(Stng>�����V�
�Q��%J���eG�߄�7��rJv��,�5�e��#�ӆ�=+Z�]�W�W�q����G��r��w�.�t�z�b�[R�,?	m�r˽��t{nu�!��z�t�b�^��zU>��zk�zu~���������v���ǧ^��'γ�\vd���:�K����z1~�%�ԻXכn�K�S/ϧޙ�^�Q��O�j�z�u�:��z?�6����N�^��z�|���w?Bη�9/?������v�z1F�8?�}꽯��2��+�N�+7�U��W�S�	]o�Q��O��>�����z{��;�S�.]�y�]/��#�E]ѹ^��g�K�S/٧�4]/Ө��^�O�1�^�Q��O��>�.���z�����S/��d�՝�Z%u����}�WK},\+U=��N�3Ӊ�����W�vߑ��=�g�?�k�q�Z������Zc�=���޵�H[��#��H[�W�))2�����!�F�}H[�{�F�B��	i�;w#�6�Wf�!m:��3�
�6���i9H���B��,���Q�Yp:�B��j�� �W��v#�F�}���F�4�}���FZ��9F�UH{i����H���i��v�ϳ�8�"-�H��4��>ߍi}L�t��=�ί�۞�����9!��F�H���BLGh{\�R�0�����Z�Y��%�D�[�/�K�����=5�L�,�<#dY�]W�j�}����s�$��֓� xOђ��g���y7�zw˪�v�� �17m{ԝ�u�Mt���|%}�x��-|	�����|G�S�u�����:�w��{t���,a�ҏ�\�w^�Q�眤���\�����:���[��V~+���~��p�sQɇ�)�Q\��C(�/���>�d���A,��;�V��I��Hޢ�%�+�"�z���w	�ڇ��e�=�'�<��w�B}��YϞ�3>g��&�+5�?�]�g��>b�:K^���.���^u��X��5��x�yn%?|!�wum�߿A.��F�7��^u�5A�:V�Qwl/F.Q!�C�۫ګ��7���ϖ������d�m�ڻ�B�O������|̻�-��V.y�m%k|��V�n⦆��
o,B�"�A!v����n��� -�~x�7
i|W�������y7߮d��DʽUMC��3������HQi��&��y��|m�xo�gm�[d��;@L�w��<ޑe�Z��u��\:A��ӽ���u�͸k�1����]��r�}�u������O,ʅ�~�;��WE�����|�Y��1�+����k�w������KLk�-��E�I�1��.�[�<���MX�|������t[O�-�}�Gt�n��w:�κ=*-cZy�����ݼ+6��Q���6h����K�����j��%��	߹4��!�G�S�b�je7�V�g�X���\�ߚb�z.�\>�����>�\���KѦ^�>�s�Ͱ�.K7UIg��m.�3��H8�m���UH�F���!S�vD�ie�|ׂ�$й�����)�,����}h�c�[6���-a��8�%�^�5�w��g�1���ʲ��j�������V~�$(�Z#���*X��G�R��Q�*k��=ܫ�}4���d-����(��zvײ߾hc��=���9D?�v���=�*��c�|&��R�m߮ûo\"�od}�"y����1x���-�c���G�;����M���3d]�$�w[
����QM�*�!��$��2���HS�K0�9��2�
�]�w�wc����3�Ż�ib�?�/�]�oQr�r�G��R���� ߋ~���P�ߝ�{��w�.����s��䝽�55�h�>ǲ��&ѯ�;%�u(�)t��y�B��|�~י��ͨ=�{",�G�5�{���1m������e�~Y:Һ+I��w�1�A���E���;����ӓ��~m]j�˵�ж���+��?�U�+���	�eX~/��o��˔�/圭�g͖�r�9��8W֚j纁����C��j�vׇr�!��C7��i�[���uw˻�ث��q8u��x���2C?�<f��{��{�.�~緷~�T�^pC�8���`���<�#ek��s�����
4��a���5��p�*�3�����ڒsߪ��S�H8E�S板Pg�wA��3�y�k�T���c5=!��W�B|?�.�h��	���)�Q��@.B�)�Nݣ�&�ާ�X�7��YW�-X��R�O��)yqJ�캦�T�\g����!�	R�Lo��_�u�c�-�����В��n��cj�J[}}SX��nA�]o��ϰ֒U�U�������q�c�]��7,��c���oqǞ�æa��H7}�^>���|�P�oݩq�����z�MqcSڍ��(�i
��Q�ť����&5Z>&�#P��A#ꄹWt�2dQ��ޒ�7z��Rg����jM�^�b��k�G��sd��j;A/���Q������P=_�o/D�C���{��Z���� @��:_��h�O�����e��x�ƭ�H�TG�a��|���x����N���z����1�Qv��o���j��k��v�A6�n�{|��G�#:��Pk�q�e�m8uzu�1.U��/���GCyK�� �T�_�|�#�I~G�Y��� �T�a�,?0����o�����;�݁H�J�U.\�����������Q�SW��m��h�0�����'��������u�*߽y�k�q�ʲ�][�׏7�0�j�~�Վ˧Lʘm�i��oڙ�H?tl�)�̚�G��Ҧ��(S��h?�d��q�)3�(S�21~�D��Siѓj���W��vZ�e\uv;���~�ڧ��:�.���i?i�X?����Lo�_(�	��W5�5�J��b�E�n����>T���"��sc���}�8ҁ:�Or�����-�W{��&�E������;�_4���1��z�C���+������	� <��;�(�����Y��}R�7饭����m�D��o���y_��y?��y�w�x��w�xg���xώ��xG�w#���e^k���U�%��w��}�E��Vu6:��E��+���N�i���r��1��,���OUzc��ĩs���Z���=X!�^D<N�k��~G�X�-L�;��a�n���,`:�[���C4>�w&4���B�' o�x6�V�g�h<�v�'ߪ�D��5��<�͚*����|�<�[~�rXӢ�"D����w�dƒ�6��]���e��6��hKFx'���)\�兲V�1��z�����\:��k�7D���x��o��+L_(��9M�W�$�]S�?�/�Ө˸���~��=�D?��F�t?�QF~�O��y�9_���h�~����F�u�Gy�1�S}�Q���I>�Ե�等����2e(V~T�{ޞ���0����!���k�v��̀�晗%S�-|��^o�{#��M�Z?���u����o�}޿��|�Í�6���CF��F;�v����ݭ��=7�����=�i���>~�s߷�>X}�z3��lU�9�G$���������g�>Ǟݢt���H{��Z'@���z��h��	�-������,��8׾�x5�@�«�4εܪ�b��S'l�x	��Ƌ�4^�^㫀��x�:�SϬ�8uK��k���x%��T%C3������B?rs�u�d�W�ɷ��䙲��'?��/�ɯ�Y����*�zOvVt�1�)��>���?s]���O0�Wy�������\�Y7t�_��2�=WeG~�O�v��u��S��i��Rٷl���g\7}�U��߇������z	��Pߡ��D:L4�D���MMn��r��Z엻{l��q���˻��7�c"�J�Y��!����Jj�*y�K}�o�l�_�r�+���=V��v/o�(����x�;0���aB
w���g������H7p�=�g���wv�ƁӶ�{����5}�&�z�?u����t�.��.����t�֧n��|ք���V}����4r>>E�$�}����P~_J�G���C��������\4ht>�����Uy������Ç;��s�`�K���Vs�l��vW�I��C���&�=��|o�Y���}����������>#<ϴ��[��VD�?�4Ω��ַ��=�:����o�Lk���Ѱ#3�|G[��w|/Uەrؕ=�#'®Tj�N��+ro:3��5�����k���|���	ڦ`c���b��g��>d��,�8mM��fk�>j��Ϝa���#l�2q��s&��}�8���Č�}�h�������?�����?{��?#�3��?����B�_���x�w��h�^K\w�y��7���:�z�O뚉~l�e/�f���2ӇL<���V�5��d?�����4m���\�c�|��J;n�Uj�d��Q��t���)2lM�ek����G�ڥ��}��i�zޒ��l��]\w�{���7�_[��6e�^�NkV��������Z'v?�>�.�l�Z�Yz��+*�Go%��B��Rշ%���7,]����1�4S_]�}����F6�o��9�ϯ4��J��{ڏ=ج����g,����a����Y=W�w�Q��~_U�����E��w���%u{ֽޓ�3�Mn~/��~���2�[��ciW���|h���~�g��}W��ûo�������e���w�]��qo���I�S=��۝o���/(�g�|�y1���P��]�ez���O���������|�6>��~�/��{���v5��{���g|o�sg|S|Ɨ������c��Z?�{����_����3����c����#�W��Ws��j:Rі5�����O�x&��5O��xf��w�1�����qD�GK�z�WsXt������o��k��+҆ҿ����
����Ж����o��w��@��+�:�0�0���&��q{L��9�������D����5�߃`�.���y��[�m�����mw�=�����1���=��jl����������c�3�f�������_5Xc1����;O7�֬�.�3�ϛ�>�g��ضP�2��s��>���1�=���;���������8�8r�[5o�t���o�V�˱[��ϸ1Ɲ�g�=/�mr�9�x)��~�n��p�/uL��#ǺI󺾋�2x��X���S�1�{�1���C��E�)3����{J��~�~C��ϱ=��w�������3D���Z�ԟ>�i����A��H�����G������SX��RYC�r轖(Y�qT>�	A�=�&��׻�𛏟6�����>���������:�m�������}��A;�w����ݟzzt�>�?��'{�'��	�_��(�m����^��N���h:w /���֌r��>��袟�o�x��=���]�E�m^�
�oc���R�T�k��VY�z�˴}�mykwa\�v�϶�G`Ҳ�T��p0�Zg�F����A�NX�ڋX����n�oI#e�w���z�2$�S��X��p�j�E�[ՠl��hP��wY�v���n��HI'�
2X*e���v�̺v%����}���c�h�� Mo,�뚴��w��F#]���䳴;�mⰦ����!�p��g���z����4@�J�9Ħ�M]��ۊ}9���o��C��Q��n�/ޜ�Re�H��:b���	���SΗ��|��/<�oX�Kg�t�y�s�=On��C:�S`|��>Ox|E7�f�Ů��������8��DA��6�%�|��/lpD.T�)�8����~����=u�C�P�#�Y�]y�[��|���G��}�i<�Q:����#����!��^y@t�D���ÕnwQ�=����?N�ߋT�0�n�����K�>�;�{�u��)ܧ��g��{�%���Z��,=�:�s��c}�6��W��@�;������:�����{
�Ӥš�2����5�y~L�+��Q��e�]D���$�间�~�0
e���G��;�m���?}.�C��+��b�Q�5�q�ޕ\�~�g�1?����2E���A�i�\D��j��}�K[��g����=~�f������}��L8�;Ɲ8���+�}�F�; {l΋�]эߍ�����..i���!�x�F~�R�a�!!��D^E����F���6E�i�`W`[�X��4��B9ac�H9��r���yߋ秜�bZCP|i�.�Z�k}?�����.��}[�}�=�Z�#���i+�����߹t���5��}xTյ�<H!�A�"5���BT��N��$�d�3�G�-UiSAK-ִ���ms}Tn�m(��
5� �dc�b��ki���k��{�yd������5�9��\{���OA��8J��h_��w�(��Bg~&{�s�8�����\�s!�ǽ�i,v����|d6�6-���@S��Vl������z��=A~A{D�b�F]��8�� z���9�ū�9�����?~��i�����M��u�D��t���Gi�J�? s����܏\��V�8H�W�J��t�o���v�"���_���uW�y��پ�Q�X��=ѵ�ϲ����ޓ��5�l�������ZwsL�#�}:�^1~�XO�fٺ�R7óY����;��7��	�c�d��ǵ��x9,��H�u\g$��WB���H|��A�%�������kø�!�fۚ����Hfe'�G��9gY���D��;�c�o�`��
g /��z�z
���pf=֟��B�q������7�Vn��%�mJ���75�o�b��Z�v����퍎��1~e��X�oz���r�����JzL���}G��(U쿮w��<�m��86��w�o��6���z�?��6Y��L��U��|7�=<��_�1-���~��?�n�`wϱ{9�/���]�f��5ޗp���q~����4C�둑�Q��#�6�no�#�t������������c�>K�!���?W}$rU��եG"`�D�Ή��;'b��G,��#i��#��#�ۡ��#�ۡ�mg�´���VI?tm����@�΃zl6ۍ����}]���V��y���8�q}2���s�����	��0J��(�Qvg��@<� ��[dI���P��33��������E�D�,k�?޳�ony+������l6:3���6��it	�g6�m��(���#��x�<��Wy�ˑ߁F�f>�<�Yh��Y���`��A\6?�x��U�g�?�mU��Q�ߖn;Vl>�6j��*��}&C;��|3�s1��h�[����o�6h�m��۠��A;o�v�`�ɲo�r���䧳k;ص�)ڵo��ۮ;*���f�v$�k+�ص>"m��wR�kW!�v���ή�Ǳk�C��w$}~|���Z�ɮ}Y���#�۵eGȮ����w�p��nz!���Y�	h�ʻƆ���Q�s��`kUC�p�L�bӊ�C��ݠ�T����^�`e3�`-�`�����d��M����%��p�ڸh;�?�wg��]�����w�Q�gB<�q|K�~9< �0W<�[]�;\�CN�F^ڻ.rƲ;�1�����݉��߂�y�\7��fw��U���S�l��ϤAܫ��.�u�;��:`����e���M�=;��F�ƈ�*�B�>3p7;/��>�ι��{Z^�r��NO�o �&nS�����LC9���y>�q�ɶ|���}�+���/����_�Y�Gh\g�	�/��^�tO���~��DU&~�5��/��[�zb��;6�����8��>l�oߓ]���T�&��`�����c��Kh�oj���<��-�z�m_	�Bx\����w�M�6*i�9�.�=
8h�����7�1�c��� �rq�úHK�������9�;Q�C��t|x
x��F}�7r��@[��;g�m�/��+�hm�^��~h�J��{���l��񻩭�m�k*��5?�	&f`�vl�����;�C~Dѻ�Ə8s	��3)�V�a1�C|�����`����ջl/#��{�.�]N���f��ho��o���V�A:BXzh�Ѫ�9:Q�s[rbO��m��LΗ���[������4��>{������q�vv&��u�6�\��-b=Q����H���V���;Lu��;�\m�_���`Z;�_c�v�/��!߷l��hۀc�
������ˏ������6�������aikO����m�u~�s[[ׅ͇I���������8��k�?�Rv��d������6����uf��Ot��=d@�+LtX��`�t@�� �6�w�xF�CN����?:,y����*=�	z�?�M�3�M9;E��ñ6�3=�f�>��M�3�M9;�M���Ҧz�p�6��CdS�^:��(�My�P,}�)��?|q6e�ɦ�B���p�6�Oߜ}'v������0V:!�X��8c��p�����B�5���}�m;� ��ec�����v������]G�U������qѯ��g�q�_�}+�qQ�!9.��C��N��Gbi��ijMa\���+�qQ�'�����Z����˖�<[�ih������y�9��y@W�����Pּl�ћ�����x��6*h6����a9�x(v���1���h�}��./�\���%�]N�h�d�l!;��z���sv�Q�	?���Ʈu*;,�:9�`����Lg�Vh�����Q�S��\O��P�^}�HA]�⬧����X�������Kz��c�b'=,�P:-�U�!H��A�~b¡��-?H����O��������`�������LM/�'ы�I��7J�t�`�z񚃤^:�h��'ġϗ�,<xqz�fҋ�*�������n⛞�F&�^B�ԛ�L2�S�&*[Y۲�[�Y�_���(����w��QCI?�Pw�~Ի��&.:�G}��?*�-�����m�,��Gm��~���Quݱ~��J?������绥u��?j��s]�s~T�ɏ��`b?j|w���A�GUv_��y�g��ݿ��N��O�/v$��)�cb�a�A)�t��/v$��I�Šn)/�u��/�;@����K�/
��oš�ߺ%}~{���E�I_�u@�pw��b	盗�\z?j���U�)��i���n�Gy�s~��ҏjP���D�W;�w���K�G}�_�Q��~T�������~Ը�Ư9@~T�ۗ�f9~	m��)�,���R펯���>< �������v�4�9п���ҏ��Nݏ�[A��G}a����G�ݟ��~������ߏ*�O�m�O��&Ћ�RԋW쏕�_: ������ŭI��$zq�~)���?u�ص��b�[�N/�ы������>���Ӌ&����������g��lx��Ȥ�K(�zR�I��ˤ��d�����Jk>�i�Ö��a��)��e�*��K��7�"�H{�S��-�iZ[�5��2���f紝F9���'�W��][���rmYӾ${ =�#��Ic�>Z[�>٠'^8�u��>�x��� ����.�%;�Ovμ��9�N	�죌���9�����S�Gk����֥c_��+�~��>��}����@���LI�m�>U����_�r˚��{��b��
��1�����#�+�#��|��=w�ake�=/wa�����z	u��.�W�=���_��G�1x�[i}C�K��G�D��6��3\���YW}V��>�t������zCWj��+�>�J�Ͼ�%�ygW����E�,�7�N���g���g�B�����g�&}�9�����g}���vl��{���y�zoAէ�[�F�����'}��;���_픾��N�v��~������ho��N������΋�[��N�>�)}������]���%��Φh{��ܙ���j{���;#�� ����s�( ��q[໿9���1z��w��,(mgU>� �ۂ�:�Z��5�LHk�Ҳ?�tl�S�V�\�,�7��ΖrZ���5WR8�n��줕�'a�e/����������a�w$��p�n�~o�sm����Mb>I6��)��d�C�r�$p�^i�M6`��d>�W؀�.�����v�T�����E�C�1Hڂ����p;��s]�i�_�Ev��/@��i����_���p��8��̮��������h�v_���il^�K�%1ҹ�T���g)����E�#�k��D��<���Hd"�f7�m6	l�S�_������~h�"��W��4��5��=ͭ�y��u���x|;���l�_p�1�eU8��[ss�6�˹Gw��6�����.n=�����~�����̭��@�' ��{�ì �U/���w�khA��Nt�����Jy��K�'�,~ ۱��܂������xw�Mv�	��Fh������-(���7����^��۩�:9�f>���+X�}�.����d
��Th�iP��B��t�#�}�ǵ<��t6mw�vq�6�{bm��Ni�ݓ�M۝Ħ]�Ħ��#툱{S�i��!����KgӖıi�q�k���7�\�M[b�i7)�gO�6�{Ȧ=����+���}��`��W��C�+�m��W�������C�+��#���C���/=�^��\ľ�ϙ�̾�}%���+�� ]�}>9b�����������)�w��?�#�<����;�� h[mN��m�$��wP\l�';�ނ���:^�4~ĹK�G�Kя�7�hg�%�u,�_����������;p�̚���c��z�:o��It���:����cf>6���5#�[	+SKd�:G��o��s4g�<n&��W��7��n�}ui��?�`]��9��z8 �0��4C�f�����{힉|g�W�g�n����U<�g���`v��3t���u[f�-;X���t��}&�q��#xdC���2��	�ǅ�D��={_�C����so�`�ڧc�m�O�{��A�x|��jL���Y�����3f�J��g�\�'�yhg<�l��2�q�o"x�ʯ�����H><xOR��g�O�
=����.�e�}�a������"s���6և��~���)��h���nٵF�{x�K���_xd�x6����P�،��t�rC�nٖ�#~ኬ����e�Ƕ<q��lK��9o�ٖ5'�����~�ַ�Ά���g��7�_��,��?f��D�?=�M���;��7��Ѷ��w�1(�m�{�2��6����w�k�g�5R�k��y�\k�qrS��w/���g�g��~�Cqn�+,������p*qղ���+�'���9;N��f�8]�mr�|�s�q
y>�9cN%�'s��S��d�'^}&�X�c��xv%�Ֆ:���	�O3�����R�[�)�~���"��O����tB�~�TҨ4�Q�Й�u9m�S�[e��p��;�wq��6�d�]���]��<�>M᳌�"����F����ގ'���7N0#N8�<���(��;qov޵��A������i�(2�vxv£��
��Y�����0ޓ`�� C(ov5ԩk7�����-���z��>�����*�V�����v' 3��x9�_�)����l*��]M��P�1�7O ��߳�>�G{����g�0��N���w�Ey�R�Y����yg߅���h'}�i����>�����o$	���8��9�΃>1���ʲm?&h�=����@Z8���s���z���Oz_���^�N�`�
��o8��R�z�b�&+��U�H&�F����Ncy��ze�C6��2��-h�>՛fk�5���mEuʍ���hZx�%��u����鈼<�� �>�a�z�|d>�e ��|�.V^��x]�x9�{�dL��ޮ�d���4�ׅʜ�G�S�\�^���S?�􄍒J���5�~���b�e���+�ʃoy��%I�c���'���QneC��$U9����v�Y^aY�<Q&��c�����M��/���.{�'�D	�;�J�$كwWZ���=��2�$�;6�e�5�\E����Mrrp{kؾ���rۘ���Xy��S���Si�ןJ�y*���2��<5`��SYS:Oe�]j���S9��?5��S��?5���SCZj�C����}��Ci�z�:v���u蝯���1�項�O��j<sbhok8�cq�{f��ͷQ{g�Ц��lG��oooL�6Øb����g���x�{�Ç_k�񻈱=��w���ţṜ�g����d2İm�{eٷ6[g8��n�5�<�znu�7�e� �a��f����n�\nC���Y9��|�.F9�鬎$ӫ8��۷by�b��@<��]�q�_�+�/5�1�A@��c�y:Ho�#����S�>0�[v����lݭ�K2)�����Ɵf�4�x��> Ҍ�t��ul�	�Y �1�J�V���Og��t~���ΊwHc-�/܍k�).�f��K��C���n�p�צ�ݤ�ݠ��*�]��b%���S�#��R�+��;P���4lG��i�ս�'�^
����U�_���}��s�/�K�˿c�Gs���`>k/��G
�mO3��8�s�^�嶳��H�P��嶀�����ٯZv'��V�C�K������ ��T�S�|Õ��<g�i��ϫ���)�g啱}G�}�J�'��3���0��ķb�]��g�����V�}_��}�<������S�V�{�8���#X[���q��ç�uޠ�Y>L#���mJC�).�!���\G���#w���~/������
x�Y8ϰ6d����[�&�?�r�Z&��u(�7,l0+�j���f��e�{28��?`�r�?�NI�M�/����n_�k�>���vd&�<&��� ����6�=���9|�Ӕ��n����c�+<�����|h5��<���Is[�4��~q���T�0��|��U����N���nagE�^x7h�U�᧼)yZ܁�_�o�����=�b�o(e�/�i�������SK�.h���s0�x�Z�dicG�<�7���O�gL&����ˆ����A�P���ү�����ƞ�c��28�75��\nb݋����w��q=4}Ϸ�>�|@��u�B�Nn4[F=d�Lh=�y3�~���%g|��v��y�+���0��\ۼ��6�C��-��y����3?�^"�)�o�{��m�������e��2��7��_���u~v��pl*죫p?�W�Ѻ��<n+c9̺"�<C�����>(�%��bT���siư�����} �g�^i������
>��UC+�i����Zj��w��¿��������;����\�=��w��Ŀ�����r�����-�j �>��w����߳�;����,�=��w���������2��L���-�*�π�������t���-�*�O�����,����w��2�w��w���9^���>5|���Ҷ�ϞF867n��b6��}��l���^���|����+�ދa��6࿆�����Ɖ����8���G���|xxon6�A���O��:=� ;����p�]�4�$���kZ��\���/���y�8-9N#߿���.{�ԀeN�v��ӳ��r�:����۬�3O�n���-S.;�n4��ߙ����� �i���J�FkL:(o��B�d�v^x�e�
<�i���|���ks���ߗ:k��<������m����+��Fq�	U�PPc>&��59�6���rl!�R/��rz�n�[��B�n[�;T�sE��|�HDF�n+��z��)�-uۖ��]��P=����˩��� �r�܍!���z��y}�g�A=(��k���wWT��j��`0Z�q������!�	09J�S��Ӹ�W�y �q�=��f
�yM��h�= J0�sۊ��/�h�s��F����ƅM�!O�{���32�Z���[������xj�B�2ވwN�r���t��M�B��N�����h�B]w�2���lg���'�(iBܦ@���NG(�^�r���jB�p��N����y25��Fk|ƴ��D[b�lnx��`�C��~_ y>��|J���"�JϪ��o���@-
AU���Qt�=Ԡ��tc�E�Vĉ6՘�i�n7��k�[����m5M� �|�=�Qn��P&�`���s7�"�@ݍK!�n\�y�]e k߃ub�k��-�5��^[a
;Ӕߪ�i�L��7S��
���}���q0s�; ߀j�HP�9F��P<�T5.˂����YTMj��zѵ���Ej�T�� �R�_�i�Q4C��aԼf�|^�����ޔ��gݧťZ}���1й�x���Eej�h8S�gy}ΐQ��G�:�(���eaL��}M�K���(rѵ�FQ���M�ڙq������M:?T��Ҿ�c���Z�����[�3��F���x�з�;S�za>H���J7���Jq��\ ?�)JQy8��(�BG��,m.��|є�c#U�a�t�de0ޜ9j�(�����e���
3�0L�{��J0|y	C�[L�Y%��:����Z/�2�V4��}����q���\nC�+u�N��P��|�
^�����B��Ǹj��D��;k=n��v��*�:�4t��������alX���w6���GJ����x�1A�t�@�"��Oyd��� �MM�o�	�v���6��1� �M'�D��0?�� �/U��O�?'I��	R&�#̘������
[��p\n�{��4N�(���4��+���L�VZjkA���8a=���F<ᛴ���	r��E�d�0������he3�>H-IZ�@�*������Y�����*�MA|��#(QB��"��k��� P%�P�^p�����M,��	�t���
b�!�8~�L��M��)`�����A��q9���%�#1��[�k�'� *8l!��p���N_8�m��*[���Ι��;�����B�s�Ϲ~�Lւ�\(�t�۞ZOͼ��gBtz�KU�������8�A<�l�q�B9X�P�ɷ9&��^gDW����p�̅,�b�z����F[(:����)��H��&�N��2���	����3r3����Y�W۸w����P72�b�l|�6�7��/$?5*����}r���FlRC��h+E���>��X�\fW��D�w�d�YM�5��M�:�Ãk[��C
Κ7�2����y�=':�PR�NM�����Mu���52>kj��h �(jj\��[��>�<.��/z�!x�����Z��zW���������_�A���l�6q@no-ċ�����n���T�./�C���l��R�[���w�2�\���0��h�a1.�ߪ�c���h�p��9�G���[;�02���������O㯐.�+<��TvZ�4�����w<����{+���Z4~���ǅ�j�~~1��-Zd���P#��꽖��ǿ�=�o?�����[s�b�\k1�ਫ਼d1���b�
�qx2�ɻ�bL��h��8���-�'j����l���ܽ��l�O�u��7L.�>��L���x!J� �'A:N�s�ǰ�k�ƀٖ�����y���Q����ic�,cӠ��@Ǆ�K�7��z�
�=���i��&��u��e0���7&�����
f9f� \���p�����I�n�r����V� ��r���$w��6�?�p�)�x�&��u6��?��IPԥ�~O��5��1i��y��!0_�6��cN�u\<�_��S��3��M�9w�?-9/�"���\_�n��\�p%�G�:���)�tug)�1�X|P��?�u��'QG�sk��7�?w�W�u+>�J�Dx<�7���t���@ݠ�C]���^?n9/+�hk����_T�E�a��G�p;���|@�QU¡m���\4ߵ<�#a���E	W��#6�s�1��Ж�J�������Z� ��<_��-I�u^W�vO5�;cP��pX�v%=��*Y��==|~��C���^�s�o�t1�	w�UZb�u����peJz��������-ƍ�p�7��)��p��	'�L�m��Ű�J��M��oM��Xo1>)�M/�_�M��Ea�e���y��:v�����<��b_%8���Fa�h�{d�[Ρ�Da*��:SOľA�`���C�/�:�d}W����.�����(L�:
���:��~���~ODaN(C�w�	�g�_rE�0�pR�[���bQꏞ����~�� ���bl_��c~�
���	�Ʉ�l�7�Ϙ��_����z>d�o2�7��'M�s&��E����z>d�o2�7��'M�s&��������&�#&�f�%��	�񴎟���/6�M��L�WM��&|�zo[��+L�*�%~�	܄�i�'M�W>��_|F��0�;L�%��x�:~�	��7u������t|�K:~�	�Ä�i��X��X�W��U&��)~�	�˄������D�{M��&�~�	o}Y�������&|�	��	��US�Wu|�k:������3_�3�u������-:�Մ����:�m��u���m��E�t��&�ot<3�|�[:��m��a*�ߵGǿ��T��:~m���Щ�gw���._�O����xc����M�&�҄?g�������:�uH����U�u�밎o���O����Gt|��}T����F����:�>��Ca�R���ҧ㫏��w\�/��xoD�oyW��xWǷ���/������������u���u|�)�wJǟ=��t��t�y����?qF��Pǟ�Pǟ��)�����:��������/�H�7���XǷ�U�o������:~����Ot|�':��o:~��t|�y_y^Ǘ�]Ǘ�]���������/��sA�O�z_�~
��G,:~�EǇ�t|s��ߙ���u���������-t|U�������u|k��j���8P�o���[st|� �c������'su|�o��]Cu���_b���V�c�����G���:~k��o�3�g�)��:>��/������r_2ZǗ����1:~�_}���^��+���K���fxק�̸�␆��-��3�����?���(����%�.��uK�2�'��n�ؚ������|Q�R`�~��g�'���X����9^��������7��{�#a&<:~�:��S�e���L��^_Ԩá;d��2N��M�O(0�W&|�_�W�u|�u|�u�I��	&�û��GM[���M�7%���
�'~qȔH�΄_Ҥ��t|�r?q���O��	�)O�)�ڕ�K��V��s���Xǻ�]����hDx���O��Y�_'^��טҫX��_�Z�w���&�u���Z�㻔�L�S�MʯYq�U
��D�3�0Τ���M&�f�ۄ�5�]W���U:��{?'��S�M��WKxE��%W�꣤���"�,N��k%�Y�8��`��q�u�q�o ��"�v�qN���8���v����LE�^�q�����P'r�#�qnu��0γ�R?�U�Հ4���nP��'��U=I��I�Lz�5şx���A�6��&�'�v_®�/o����c����L�M�ӳK���Z�L����R���|gn��ui�,��9��o��	����[%���M¿��>�TU��5E���!M����a����&�Yu���a*�I7�,���i���1碩2�	�$�(�k�^���8�ۦ��+�&��:�T����+o7�	�`�wޮ�ϸC�[���M��
l�'�}�P����� ��q�~n,O���Gө����S�_��+�@�;&��M�_I�����t����o��NZ�|J����ɻ�D?��_҉~"=�`R��!�,�? �o��(C/�-z�wd��0�w��b�ڠA�?��g�ɠ�\���k|�s���a`?�A�����e�������`���!�f�5��ߓA��l�pk���73I��px4�Ei��/�����V_�I�'x|w&����L�Z9�#%=l��..��8��L��q�x&������5 g[�@�N6Ǐ��f�¥Ⱦ�[8�����c�^�/�r�,ϗ ^�qx3��J��~$D��Q�����!;/�,�W%<�T�C㉿��E�c�}*n��n ��į�.����_�Dz�����9�{�h����d���d�x���x����l�Y��g�R�LQ6����[��A�,���4�(�sC��� �������&�M���C)ߐ�:~�@�D����Od��4��x��-�i~D��W >s@�i �B�	�������]J�� |^���@�_����9������=�����6��v���s9�o}�g�r�ws���
�%���m�_�{����2��(9(�{(��
��x�+F�g \���t~���
=��q9��`�D�V��%��y�u�g���U%�� ޢ��@4F��� )�B������Q$�s{.��V��| ���n��W ~�}��\�����m
=���T��璿+��c���.᱃i>Z�c�%J�?pw�l�;V�K��Í�����~Aȿe �W�u0������`�����]��{��_����^��Wy���9 ���R����yj�w�p�Z!��m��(�_��!M�����s��+���Ch~H�w�PZ�!ҷ�W�ODX��-Ci�\ȫ�Ci����\�������q(�������� OV��W�;3��_!��R-P��+����Ǖ�;٪ӻ�J��o
_k�4� ��	�Q��]+�_	��͔�~+͇��� �9S곂a4_/���a4��a7�+��V ��s�<����A�?���r.?� ��R�7t8�w��6�֗}u-� ��e��y�N�#B=>��+,��� ^�����i>@�o�pZ�"�;�Z%���8�*��4�Y����c���Pi�{ޥ���^%=�OZ��� OT�O��6��3��E�n�X�o�o�wt�?����,�{U�O������E������o \�8��-y�?����-�2~��	~#������\���h>���?x�B�ܑ��~,�^��K$�nx�A�Yџ >����HZ�$���HY^�Ѻ�4�.��F��D��+#i�R���z}O �U�/�2�f�D��(�7)����h�A;���c��� �`Dᕗ���Џ/ll|�� �R���WH� �����0��*��5�������*Q�/���A�e ���0���(���� ���B�l�H�ߛG�z7��1��ޒ�:0
�G��8�;2-Q{ �I������BQ��|��8���zy��@�_�O��D|o>������~J	��)�������7��i}��?��x��_��п����87�)�?�rZ�$����i=�h��\��p�R�5����W.��N�^���sh-3+/�{��i|Z����@�i���\���2��g�}y?�;�����q�|��4�*�ϷG����_-�<��Ѵ^B��x��.��돏F�|�������o��z�o���ctz>��C���޺Έ��� �/��~h���_�!�lo<�z��Fԟ� C�C�_���}RV���0<��+��M �+�8[�'�|����$G��h��h��h>���c�.����D�c3 �{]� ~q�����
ZO ��- �^�>��8C��{ �U���g|�X��k�X=�������_��oI{� �*��wV�ݱ�~���7�����C�7+���L�����#]<��+u|��`���ĳ�q=��?x�1η�����+�I��x�R�?^I���m4U�Ï��z����=J�*�׀��"�W�R�y�g;��\��ɒ��/���F�g����KJ~[1�Ҟ<n���B��[$�:���nIp�Ӕ�n�Y��G��D��q����C W��`�R��q4�R����7������G�B��@XIo?��
�7�ֻ��x��֫���^���+p	�����_E����]�����7�/*��#*��N��]�H���J%�?_E��N��j��g g+���M�/����p����	�_��֋
��{�'��ۮ���B>���	���`]��g�E�? ������Յ 7I���BZ//�_���^������� W+��G!�g{y��\���zw�� O+���)���?d��j���x<�G����>\��d������T����
������i}���^��KT_oO�̈́}���W�~Ⱥ�E_������>{�쟨oʯ��MX��_C�!O��kh=�h�g���B�~���O=����m�}_#��7r���?��?��ԟWN����4��_	�r�ZO&�w�Z�'�ŷ����o6�����@�G&��U���A��zb ܦğ��C�?�<��$?���u)�W��ya�=S���'E��B��"ZO'ʳ���"Zo%�c:<�Q��kt��c�B�1w��I5FM 5��A�ܲ���9�� \>G�׷��u�B�@��lZi���^w��t˭7�?�Cn�u�C�����jjhx�(�C��AMVB���~	��d���'�#6d��G`:�gVU}�1���eUs�w8&�o�"L��H!�q+�й���E'G�tU����b'�����FFu�ߣ@��rL�U����@���o���k��mRƃ6C�h������g�;Z~�HI��_��"�Ǝ$�_:^�`'��p,u�P�-��_�M��遺`4�rw4/U��o줐4����ɒ���`G�8n-f�
_��^x9�5Z�����eU�M��A�Cn ��❝C@Y�bGñ7:�%�ޛ�� ۵]^&�����X4���^_�c�J�4���Y���.���nw��A<��S�Z8}�L����aoﵞ��Z���@�a�MH��>���}(
�njR /�/v���WN��b@�M�A�'a<����ϛS���#�E� ��;+̘^�X0k֢�U���3*f:��b	鈗2<\��o�U��(��»��V��AC�WZzgŜe��&�O3	������~� A��4<+����xqX���n�t:v� N����]PP�-t�^��	���ԉ�\��z2��/{똌�7>�����o�׍G@c'$�l �&"ŉ�t�a���t6�G�O�Y�s�hU>��@N������OLT-tךS��.�bA�c2널���O�t�,��|XG�f�i�t�s����Z�N���X�Yp��� +P�9&�����G�J'�2�!w?���D''�c���� gH��b��b!NO��[�����Ǒ�q9�^'ۀZ*�f���͝���쬧��F쨒I�X<vrm*��<$+d>���X�� RZ�q�����.8�D��,I�۲*�����\���^05������1oSb�*�
��ݾ<�U��TVʃ�x�q,jZ���0^�t����qk�g<�k���������I�\�@M0z�*���r�Q�Έ&�U7+z�0O2A!ʄ���x6h,���I:�-�F�x=��g�����|�=ة��&5�u)��	�S�ӎJO^z�12�|�Ɛ4?}9N,��{��ew2�6����9W�~������Xl_t��YQF�NE�ɕ$
(j�{u��G͛T���c�茢��A��DW�CqF���(NbMJ�#����$�M�@��bb+�ଭ��3�E/AMĵr���&�@�iM�0����8Y�����Lݘ�����x��3�؉�g0��q�K��l������o����Qb}�����{��za�������:j�-��J��":��Nq�65�4����5���NF%�g���������c��d�R����E?�&O�ᢴK�d�ɞc]	��70U�vɺC���X�N��u<'�Ǽ�L6[��)�D���=>:+�%�G9��	z�V��x}���7h�������Idh��ʍ���ɄIFM(�%J��HK�)��s��G�r#:����`)���Nqr��$*1~p�qz�������+�ǨL@�xh�r;0N:K�X���(AS#	��X��}�d'0�RHz$#/�^�B`vRO}�~�9�\i�$�Sz��S�%BTP�Xd'������Lȓ3�+U�$�?A6y�w�d6g]G�8�����ƋT�J������Ģq���y	ۓ�,���8F��_����y���PP��䱫_X��u�·���H��'`וJ}L�_���>	Xt!��A'2�8��,�^�t��Te�5�2��p��Us���L��8T��s�<x'���AՉ�5����朞����`�M3?������*�Վ�&:�@�x�p��C5�qՀm�R�gJ�~X��Iy��6���\!9\��1���iY�FtAz�}>��f"`�K�x>4��Z$W6Q�X�N�F�W��)�%V62���zV"��![��8S�,�f�٠�U�;h�9��x�]�b%JTQPPÄ��m qڜR����8���DU�����x�Q�u$�Ր����	k�Y-q��(���p���@Je�^x��%���H
]��y�u`?^Nl�j��g2Y/;#>���Ғ����fi���[���؇�S}���53�@D�$,f��4PA8 ���sA�+c�I�)�K�p;j�,)�)^M�uE���s�#nz�ڼI�Ƴ��D��ˋ�	'�jq��#b|(4��DS�I$3�S�L����)K�:����Q�
�\�t�����.����e�
�+L�{�j��ڼ�e��(�@��mN�� ^GџM����aI�d�u�2y��|��N�l���E%��Bo0�N��_�&w�����פ4~��m�I+e�:�b��d��T�~1pLj%�0�.6K'W�X�|o��St�O�>;4׏7�:O^0�h�Q>	&�c~rHK�!Y���s�;��X����1z_��Yѩ��æ4![�_4D�IJ֟h��17��JK��Q�3��B���y��b��Ŵn'MZ���z�䎥jI'��HܑP�)·n'�qO����z�nm�3_�j#.��}>j�x^Ρ&ʇ+(�0���,���],��`�!��)�8�uq ���ɍ/u�6�l�/�U���1f��Q>�Lj�?��
�<�h(����3���.��!�c���or����;urL+:��e��˿��LJ�b/�`9��OHt�Dsj�q��R�l@^Ol6�?�-�J�=��b��Tg?�!:)��$[�@�����g�>��#�,���{Zw���[yQ��vtkZ�L��:M"�+j;$��U�����\kv���+�:��2��+������&��`ۙf��i"K�.��Z�^��PK
    +Q�H
t�  � #  org/bridj/lib/linux_x64/libbridj.so  �     t�      �}@T���*Y��N��FEVFj�(�R� ���,jjEźad�kIeefEe�T�e��fVJfzW|A͗L噙3ww��������P�{�s��9sΜ9s�=����}}52���MH�MSt$��+�<��SS�����66�����Fg�)��E�	��kK:{��\�y�0y�����>dyv�8W1����n?>63n<�<�~|N�˖���g*F�y�5&��~�#p_��������W/�\��Y�U���	��d�7h�������q�&..c��ś��Ϻ�����q	�;��9��,'�q���)p~� ��9�7�p�������ȃ#��&�����_��)8`�|=�y��1��3~+Qp������,��K��x8J ����X��N��'�hGG��s)��ǿp<t9��z6��:����W�X�,8�絢�������oq�:	�A�}���p���Ƿp��c���H/�떍T��ù3�:��L�~�!p��^8F }έ9�3p�qz 9����p��h���@���^��pĲ�<8v����p��m��+�}���Fʧfz>�u� };�p�±��p��y���D8Z��η��2�K�X��c���;8���G8Fޅ�z����8�2������|�
�pX�^�p}6aߝ�z������p���y2 ��+p��p��c��x���'8��\���
�t8^���xe�9�ƾ�eH�s(��@��#���y����H8��r��h���#O�u��c(�Gcp���/���z'=���3���w�o��-pݓ����\׾ط�x�c��K��t<��h�����p<xA#O�q���{�g�����"8n�c�����p/��)�F'~���M:�����6���
G��1��Hj��iO���|�<� ���� O�s�!��v������8����8fp��w���@W��(�s�x�"��[��������p|G����p���r8�^,ӛ�����<����p>s�z2+8�x��kqݖyob��_�˸�������=�����qp�+���:��7���N���=�p��#@`�����:<i�6����:�%�
8F��c+�^�b/ĵ�!��pt|$��1>�{����]������W�z \?�L�^W���Ap΅�E\c8<�<���2��^�T{�3��/�Y>�؍|������gp����u>���4��>�z�1	���0��6���H����(��"�ƩA&�&�ܧ,&��_�ϣI� ������:��V^�28�)����hU���r��AU���q[�EQ�-���<XXf��䫷�O��5�$4Zjz,��v�[BM%׆���E/���5���ʄʢǋ�5�#��鯚��{~ʰ����wvҥ�V�����^���EL7�tI��xMd�_���^��_P\�癗6�d*�9����S�ވ\��ϋ�RKZ���_��Ŕ�--G�bo��i��K�]C�6��Nh�bY�&�z�ñF�/���������T��#����a<�� �M�z{�Ԙ����c���H>G�T��m�c#������8P�+�h��1��8�
�7{��x��n���8�c��0�@�:�i�П��#�1�w�'�mb�c�󜆶[`R�����2ƒ؇����s�Oq\��c��8�>c�����e���G��y��~�Ҥ�w���c�-^xq��cƉ3a�#��1�/�w1��}K��1��X�Џ���S|>�g��09/�\�3����4���ׄ�h���8�c���8��ǝvs��!���dCq��s��p^��;��n�]�?�1��y����x���>�ø
�i}�Ƙ�5���Ή0}T���p��8G�xcb��q�k�1o,߃�S6_�9�q^0N�]���s\�c<�se�!u���!�\���|���|�c8�a�3��1�����q���|͇^_��ᑟ��|^=���EM�j;+�|ۆ�kf��ϼtAZ�����s�5ot(_ZX��Y���8s�����/y��f�y�[�V�ڑ|͌����p���fn�R���#���yx��)+����ٔ����br�/~�>�'9���a>�����v�Q���Mfǚ����|�šS-��݈�M]�|��N��9}����K�e������թ'�Bz����M�o|�����M�o�?�����k�vO_1���N}տ��Q_���z�*�����|ƿu����9{dl��O�u[���}s��6�_?2�X�Y7�_|pk�����}��!�Bn����>2�T���I	�?����O��l|�m�=;��~����R���������^�o���ݡk���C���1��A���Lm�֮��'�p�%��|��/uz�r�s]�z�R��g��Q�O?5w�pmǪͯ��;.���"kU`�ԙ�}��ߙ�ewU~��}���ZZ2���>����ٗw��≀��]s�&��H:��Ė�?���Qk�/���/��:pa��S:�e�/s�n^��k��?�eO�x��\��}���ճp}�g�;z���>?����%4�����l�cL�&E=���|��0���sz�e��c�Q������s�Y�cc�Ю���3�kM��W��>k�m���pf˳���ł��G��dz�wD^y�(����5�=4���������'�ğߍ�:~hmރ����/���o��9�y׾������2�]��Y�c��߿��/ZB�����t��V�i����Iڽ��,�O��'�sޅ�_���Ң���,j2e�ڹ�?���W�-�>����k&������k3�7���١3�ռ?��K�����yD�����7V�qn�������]'[�~�_�ܘ���?|�Q�5��q����Imz�|zȏ���>ֽ�s�g������ה<[���M���}�gM��V��jQ�����~�U�ku���\��gv���ufu��g��E�;u�_��/��{��}����{l\�f��ˋ
�%��|������}��W�VT]������[6+LX�Mv蟃~ifm�=������"�v^t�P���7;3��ѓ�8;�Be���S�.y�ܼ<x�/��x�b�N_���-�|?�>���v��Uë�}�ݧw�q������\�p�<S;j?_q����w.���OKNO�n�������7I+�{e�ٗ{,�}��/��[<��$��u�#�w�<c�����w��s��M�zث�O��,��w�Y659�b¯_��+c��oW���َg{�T�hǑ��g�򫈻�r�>ߦ�NO��_Ow_ӫ��c6�X������G������_n��z���W��=��	ŉϧ�|��?�̹��Ԧ�⻗׎ڿsk�u���m��c�[�_��LjAb���W|{k׶��?�����_�2��/��r�v�s:�p�K�UOӺˏv�Y����n�a�?_�m��s�sVT��C�M���~ +�Gs�w^�x��/M�ێ��6����~��ӕO�^�9��V�g���Ԧ/}��G~�1�ߵ���w�s�<eZ��o�Y���53����=�㦙G�,��{ʤ���-fu������t�[�=��Đa�]8���m��ՇEO�0o��?�|M�L�BO�6j.i�;��;�w�\A����Ώ1|�<����|�����)��������g;{��G~ec�����OA=�|��w<�����_y�1,��'�M�ԛ���y���id�^����yo����7�{��~�գ/�K���/֣W�z��7{/?Ι�x����é~�3�5Dt�ZA��
���{$�*�����{1��:Ӑa��[}�|E�k���8]��s��f�Fh��3��Z�^�/�I���x8@��Q�>Wy��i�S��_���F�6Q�5�=�O6V�cy(�q?.g�A�.O��ߙ�ך*�����5R��+�V�39���d��%'͐o�����{��>��@���]��HŨ?���W��Gs�r^�z._�W���9A�oD����G�a\��/��ߋ�q�\Q���\����	
�ׂ>���i�_4a9\����v�X�Y�Ɲ��E���G����v����p�;�}�X?`��F{5��|�����yG�}x��(ۭ���~a��l�7����D�{7�K��S�j�Ǳ�	��=�Y����n���I�	�^�Wx/�����f�?)�^��?	4���{������Zq;��l�S��	����3ޅ�]�����X�C��>�����-��5�*����-��;�o3���g��~v�?������"�@���~�WM�g��|���?��i�r��9�mX>?����B������3�Ǒ�C�}���~&�P?s����(��o�R���?�g99ú ��T���+?�_�<ǩ��ne���ٮ�R�,�?G:��tV���T%�K�E�f�^l��lo����󐁞vە��Z������߆z��[XN�G������e���������ӹ��+����2��pyt��U��<�'ˉa�r=��S�����n����$�������ܝ�K ��~�qd����wVx0�?'�e�1��Z����"��d�{�q�C?��������^��{�~�v)�p��S4��*^t�������줢�~��g�A߿�Y(�����3~7�_�7{��}ܯ�x���u�yP���V��I���7��}��R��\���?�?����7�	�[S=,P���G��M�=ǅ�<~��z=����T��������~U~�yFm�������롂$���Jn��O9-�q�n�r=/�x�f���0�>�	<~�����K(on����*q��8�q����i��J^xן)���S�~�]�����E1�a�
绯�'ގ�rC�:���v��y�O�a\n��I��g��p?�E}�{�E�/�����N�G3��6z|;���~��d�ɳ_�b�S�����n���,x�'Y��ǳ��>!j/~H�?�0q9{Gy��������`<����P�w�>�9�&��9�4��#\��>��l'+�!�������������K�_:�~���g=<�qT����c}s8���N3^����}^q�^��*f��1�Os�>� z{evQ��&�A������.��*�w����?��?��\�$Cy3^f��a�����r��s<�x?.�;�89��O(o���og�pI�z����9����vr{U�Y����q�nof}݀7��{��~��7}t��>��Z� :����o�t�������g��݄���ƫ�q=�����z=���g�X��_�|���O2����/��}�a	�˴�����C���/}YN��~�
Os�_�vX�C��Gϻ�]��{�]O��^��#}/Q4��}8.Mg�S�7�㺛߫��.���)����$��s�ao��������{�������ǟg�� �|!σ��s����Y�'ٯ�<��i����+!��>���p��g��Z���j�f�s{}d����>#y����T��5�)��,S�$�e��d�o��.~�q�~}\�8D��d�v�i�_N/x����C*�㺻���7	����'0��gc��+��A�k�6��䬢�e��I��w^��i��7���5�?����p�6Er��3�Ϸܾ���پ��|�]-d��y��?2��ز��������֞�����]��x��7
���^��U/�vO�|k؟t`;�d<٠�i���m���}��~��n`�y�g<�6�QI����x��wn`9p�1��G<��q��p7x�)c���=�x��K�a���k�s��a?�����v��95=�r륗���7��&�XNo���Ӈש��s�g��<�m�U��������7�0�3�m<�����r�>kn��/�u�4�+oe{��v�����ۅ�[�Y���z�q��8�?��)����,��7�����O�N���E<^�����oZ�v���Z��u,�� >�ϊ&�����?�x�Lo�o�>�����H�0�[����|Y��-u��ゾ��Sw��gy���E����<m<�Xn߄�<ǵ&\��ܯ}y�ځ��_}�+�����=���Ƿ<��=[����m-U=T��_iX�������.�p�/3�s-�n7�K�'��=��\9���q�vC9{1>� ���-�`o[x�K2ș��{�o��H��C;x}����P����,�d����c2��L��|����^��4�����c��6�w˟c��e�*߯�lW��T���r�U܏�`|?�[�A��8�*C�<�ϛ�(Z�|+Zy��R�ס9]��4<O���j8p�dZ��Ks����on�
C�lR�O�����(��J���~a�&ø���S���\�	\�z���.��П���$۳ŀ�p��4����W�vێ�]����g�Nry���	���a�>����\�U�z�ه���w�g+o��Z�^�f�xg�W��8���.�O%����1\������63�[2�	i����5�y���޳��~��0����o���!�3/��o�x5קf\���7��[r����I��m�?ϲ^��]E�e=N����i����rhs%__�X��W���K<���cw����q��s�����x�{+x}F��r=h��e�����/}��T�!N���w�{KN)|�O�c�q�w��ݏ�Y߁��q!����e�xW�/���o���Y���q|��S�Iߖq���¹~v���.+Zow���<����2�|'�G��c�}��u���S�qZ��u!��m��q�����ϵM��c2���lɹ��DS����tSb�Ё���\��<�5w����,���QV��=%1eB2
H�H�d�q���/:#9/Ϛg���?y\rtrF�%9+5Ú�8$�)5e`v�NQ�c�ӳ�S
����J��gg�Ϛe�MOqa�)��--7{|�k%�����j��g�l���m��ج�����9C��@��L�yV���SN.�bKNyRS���krV~��0ؚg�ε�wRI����k�NH����G����f�J�����y�̈́���h/���J�.�.7�R�f���M��G�sm������Ծ�ٙC����N�4c���32��C��%24p�^���2�O��ύOγ�JML���fe'fd�$S�C{�S���e��Q}��qbv��Q��c]	��c�K�MWv��8!g��\+�暆e�Op��˦�����\k�m�5�le�-7?�f��2�
�P�!le(ڎ^^��cʵ�)/}L��q �m�,_�@T����{�{I�]O7�Q�Lc�������e3�ɞ�'���N&H](0&;��|��x�<0��
�NK�E�ϳ6�sHZv.IUP�}3��<���OR�����$&%ךl�;�w���^�i���އ�e�R*�!�J_UFc��gz�����P)D�*�@�KRO]egc*�k��U��\����2�����\rU�du�����T���V���P�P�J�-����A�0�1���SS��x����M��D�s�rr�Y�ʿ���d��T.�������K��A"ݨ�*�ec뗪���K��(�^�.c�K�K՚x��X�F����fʵB~yVc�Q��><Z��n��&��rc:Bve�rc:Um�����+���c�\��`��\}���7����oRՎ�5�!��10�1Q�n` C����N�%>���,�h�ɷA�G���Z���{�ge%�LiLU��5	L����d�=��e��֍ɇ�Х�Y� �� ]�yD�c8� w!X$�\�'�*�K�A��
�˂X1"!7�2g�4�Y�+a ���[3RE�a ct�KM��Hh�ϵ���/`޳���3%g
,�����L*�'c�nz֔�d�����I�M�̣*�l�U��Z�8Y�w�����ɹ��T}Pq��S�R\V�uB���G�F�Q�AXG��1�[�Bt����kM�I�脌�<<$��-=ET0N���R���G�ZS���!��y"4s� ��7;k�J�`\���l�
���#�$u�pn_���~C"�M" D�&�� ������Q	ɶ4L������R3�f�ǅ&�ݗj�������&�>�ȋS	x����_�eA����h�IEg�ѧ�Q��)�h���ZG�V=�[r�u|���Qj(���
Ò���, �1k��W!�A6�����У1Iq"��yW=�L�O���p��W������n{�k�G3Z�M �mt���f�+����L�k!����IâҳR��������`�?�����zL�kFoU�^��F���p�����w�U�S��k�1уɥ�7��P��dh6����f.8~ҬzP\�\>pCʡ��=��8��l]��~ݳr�.�b���JA�n���
�Q�bbv�l�À�W��Vϥ�����b`׫�b�dR;*59�e���9C�gӂ@}��w���	�.O�����n��I��2E��=��K~&TFvʠ��kjC�Q� [Nv^��= �����K���=�S��IA���b�L�y��s�st�;_f��zE�y57L��:�A
F7�dd�34�S� ,�z't��0`�R��sq�ks�|^��*ҮV~bXrnn����k�� ��L��7v��(d�ͰfB�ղy�z5�T^\纪�A�z�h0�h�	�1ʹ�F��q��m���2����j�8���*R�>���!�:���9��p���W� W�L��}����DםU]<8��U�x�l)iɹWe �Xo�L��,��x�r����~|> �W�Wūl��굏�����Y�lhi�骍�*٩��q窱�8�U�*R�>��j�!�:�������Q	�_m�\3�;�K���k�
]U���QC�� W]YW�0��8�%��m���v�^�O�><�@8'�ձ�:|��̫��\^Ì9����ѣ���[��b�Z�<A-FL��I�8h/��D�<���51�q/N��h�0?�izvjX}��� ܌�/�$�0�V�{e?��84#o��YS���ħ�������XS�G����<�����%�$ےM���ny��B�c(t��j���A�)5�>�R�����Z���8
���9S���GvJΰ���q�'P�F�eb޳y�Lcʸk���7>=Kgp������?P��\)��d��!�M�8�E��{��ڨ6b��ӳ\7ed�npJA�����Sf~�R3�SSs92�Q���r��~�=��ҵ�Ȑq�0��s�nx�3^��x����Ys��,���(R�z඄<�d��T�NL�����f��':�{����]��t�M>��ܗ�|M~D���+���+�×h}�:�6�����������wV�qO^~��k���YO�1��ܲ]��~�3�)~���)�>�~�ƀ0^��'�ӕ<�la���v>���+ؽʀ'0�������_0�����~���7�G�?���>��@��� �z-U8�����x�6�|��/�y���Gn�V��o&�.��(�O$�0��\~�=T���?B�V�)�l�ox��Ox�������.�ٝ&�g�#���	_&��S�%�ߴ.������r���~X�W�V��R���/*^ ��O�\�>�^������M��	����� ���>v�w�_��� ������� ��rB���x���xi�w�&���7�~V�x;�'	<Y�I�C��|��'����G�%�A�e�G�s.'�\�Sڿ��oU<��V
|��x7��Y�e���K���BN��S�	�e��\�����(p�'n�o��Xڿ��(p��� ���/�K�?T�����BN��G
�"��ܰ)A���x������&�X��#���Cn�T ��_"p��Ce���*�r�?,�_�v�_!�_)�i�D���K�xo!��ox���r4�'�k���/|��C8�Bѯ	<�<�<��R�P>�<�<�<�<�B��{I���m����@
�r�8%p�)��"p_�� p?���BN��_x����m��T�S��x�����\��g���
|���\�~�b�?&�)�Ǻa�J�
�J���f�Or��J�{.s�J�G�	\�\��w
����﬘>u��D���%��-�.g.H��w�B~R��
\�.T���G�#._�|��>Z�S���������Gڿ���>H�o'�<N�	�������S.��X���aS����J�K�������v�7�^��x����&p��k���/��(��37.�_�������R�A�<D�x���!�)��n����	Rڿ��o8&	\�vn�����o��wx���
�D��w[�^ �9_(�r���b��zU\��V
�3�W
���7|���\�&�^���L��v�k_-���!���s7$����x���b.�0H�"�*�E�����H����_�o	<A��7��w7lJ��M�4��x��˅�	�/���ߍ.�/�_�#���<Z��.'�B�Q_)�!��|��.w����N����x��5��$��_���ܴLؿ��>N��K�?�_�Aׄ��7��Ox���o�F
�_7l�����^���F�I�!�4��x��cD9'\�np��}d�#�n/�OB��ϒ��O	���E�OrV
�i����6����.�<��W�}^%��k/�k�*�/�f���p�c�/p�����1(�x��"�'��o��/�[����E�� p�2\�;�$p���.?�#�w��K����x���
�L����9ϓ�`�1��q�;:�,ŕ��ڐ�����5�W>��Φ�[f���"�
i������n��4Jvn'z
Ҹ�$z"Ҹ�� :i\bp�=i��;ˈ�4.9�~i,�3���H��֙Dt�qj�L ��8rF�i��8C��4N=�ADwE�� �� �S���H�T�Ys�VH��D7C�%�O�ҭH�/B��&��>�tҟ�H�%��>�t;ҟ�}H�'��މt �O�V��'�����?�_"}�O�gHw$��^�t'ҟ跑���'z�7������t�O�T�;��DOA��O�D�o&���E:��'z,ҷ��D�B�Vҟ�'����'z0�!�?������'��]I�{"}�Otw��$����]�?�]��F���I�K��H���D7C:��'���?��}�O�i��%��>�t8�O�A�{��D�C�>ҟ�HG��DoE�~ҟ�o��I��%ҽH�?C�7�O�� ��~�I��!���/�?ґ�?�S��"����tҟ�HG��D�"C�=�Xҟ�QH�%��~�~�?у����D�G:��'���I�{"=��'�;��?�]�H���A�?��~���H�t�Ot3�!���Az0�O��ہB�}顤?�G�F�}�GI��!��O�N����DoE�qҟ�o�~��'�K�G��D����?�K�I��6�O��D�C:������$ҟ�H'��DOAz�O�D�SH�s�N%������'zңI��@z�O�`��H��#�N��鱤?�=�~��'�;��?�]��$���t�Ot��I���H��D7C�ҟh�sI�/� �G�}i�O�Q��I�"=��'z��I�w"=��'z+�ϒ�D��Dҟ�/��D��ғI�� ��O��H?O�=�H����H��DOE�Eҟ�)HO!����t!�Ot.�E�?�c�.&����K�?�O �2�O�`�KH��#m'����Tҟ�H;H��#�
�OtW�KI�� =��'�ү�����.#��n��k�?�>HO'���xЯ��D�Fz�O�Q�g��DDz�O�>�g��D�Dz�O�V���D��<ҟ�/��O���H�� ��O��H�I�=酤�Yj��I��"��O���&�����;�?ѹH/"������?ѣ�~��'�	��'����bҟ��H@���%�?�=����'�;�KI��"��Ot�?&����'�����HW��@�U�+��|��4��Rڸ
,�`;��~�b��Rx��x��� ���QܧG�Va<�(���������G�4�n�o�츒O��}%�߉���H��L��Y
Xi ����:���[;����iiP�Gc�3�F㟫�p[�p��&(܊�T�Z��Ld�n�|8�?�����*�=#X��/��S�k⁸ Ӊ��!��Lع8�Oq�mZ.DO��I�M�"�F�ő��L�V�5�#o8�AD��M�&%���wD'�۝����~�����d0���w�F�o����K�s�eG���cq���t�����h�>��G�����gA]�MP����������.ʝ��3Ȫ�V	ui�� 3�P��hm/��pe)����b��c���'�c�PHpL�8����h|�� �d�iyq>U�|�E�`�o�{C,��"��|Hq�}JL��ůQm��x�Am��<WI��I�����sm�hx�}��F���,�M�����Km^��� r�:�M&W�\�P1�s�7� �%w��Bew�X\�A�	��g���G��y�'��^�70���4����l<T�nw.���E,|n�����D�-wn��1. Z�ƭ��4d�ͣ�Ϡvp�}���t�I��l~�^��s�]�����A���.k=a�Py뙺�Ud}�?J[�o=����z���z�������o�s�﫷�e?�_�������9wU�����`?�'�����=g�~�}c�}���j�x�����w�����iVj�8{%�il�jV�y�?�,ؘ�>���Y�vb�B�?�j��$�؈'ګF����s��3�F�N��3H��ފ��Xj�Ư��5~W��D��a�sY�5���G�C��)�_��*?�����}7V(}1��}Xm�m�i��������s�i�v�_?��#=�*��f'��D%�w�����-<z7�Q�N��o3^\Ɂ�F����ΕXL�Lf=���?�Tȥ�8�Wo��lG}��=U�=i�{О`0�LZ�������P������+U�8����k�
{���6��OBW���|[�Ʃ��4�P���xP8Ùzm,��x,A�9������ƥ<�d\�cI��,Z�IJ7m��ЋY�~�ZȊ����a?OF�m�b�U�	��pi�I�y��x����~Z�	Wq���e�Z�tv���?�1ޟퟺV冥q�e�aP~�i���	�D���2i��H7��~;�_�/����=w�[�[q��G���n��}tL����?���G���*����U��06��ږ�Ԏ�0����n8yţ޼"8B�H~��[��i�����*�n��:���������V���~����(�ߐV����Q��Μ�?��ͣ�
��kc�����\�N�o�����a�
�\c�PJ�x>ؗ}w��g����Ə[��.X+��GhXeT�ke�@��w��u��E�m�,�����f$��i�X{�8��� &=���R[�َ�%��ly��2�yL��|l�,/�G:��|���~x�_�I{��V	�ff��o̔C�j�"��Ti��^(�
������Ü}���q2�|�A{�0�j��	��vj(�{��6�n�b|�Wߠ��B6�eAMM��J[�r�z2u�`�_�T��.m��Kl��X���0��w$��&���;xkW�������s~�����~6JɁd����X{���Ѵ<�)�'4`*m�T�D�,� ��Q��e�E�����ξG�~�i����˫ZSS��.�@���|2[�;ӯ�6c-Ў(�@1Kg�!��7������Ǐ��@�5
��>���&삏��q����GL�6�^\�e1���
�\�N*����9� *�<a �����
��� ��OVP��0�΁��q~~F����??#��e�?��`���yC�+�`:>�{�1;�vI.8�<��AQ���'�xLΏ ����Qqj��.}r��ɖM�W��$&��6IS1��x��By��r��4'Oj.��/��.��@$�A x�1���ۮSs��</�ld_jؼ<��-�<��p����/Z���J�0"y���c�%-�5k*����˹o;��8�����`
1��Pg�������jw=��0�y	⛨Ǣ�/�]�԰(�0�v|��'B�c�
q]'�����؏}ö���ݪ�,	
�~
d�6��Ԗ�nW�����(� ��zdԓQ#���J\�Z?�r�ǥ��ߨ�����d�<|��6ξɽ���Š�RX
7P�U[�C�:����y,�����\��p*0�*U�Q�q�3�C����3�(�G�VM�q���%�=}�_*��1���!}�J�h�M�ܣ�'��S��kj��?Tzk��Q�o��F�tX���"�o��%�Q��^�Sqn�"֫��]�^�������]����!�}C���i�>��>��� ������0�� Ί/�����jT��Wp"Q[�����e�����-�o�Jq���%i��1���o��|M�g~DTᥖ�:�޷L�aJM�:��hic;��OiSni�MO叞���s����x�eo��1�d�o�֟:I����G�Y����k��f��0�:����\t��݈ٙ��Sm��?�'.܅�V��;;g�	mw4PNܖ���:�ԊyS۹���xx-�.�=ٝ7�Ǯ�߻��sfk���+�i���g`1tY��R��p����>�w��+�l���0��{=��g��o�/�z�r��b�O����-�8�^������g(}�+=�r �ۙ���l,����i�U�h� �y�(������:��"yi�v��JD�O��@��܂!C�*9���?���ξ��~���_hߠ��;h{G�kY��v�a��G�gn���]�����}�cߠ�߈�+-�c���<���\�ݗ�;k��� ���G���v=�^�W#�=:�*�6�[���#W?��G��갟��ﶤ����mRC��9D�cM�� �Ih�ǆ%!T,;~(h!����YR6�������x��h5--�k���K9��c��cMկ������1b.���ٲ��GPz�~.g	&���WT�W���8��>L�)��b=�\��-rT�z��rP������D����S���=��Ȃ���7b���U!��}t *��~���GK��f�&��2�օ�u�Z�`3Q ��o��*c|1�6�]�u6q�G�r4�{�}�|_"׻���qL��,�yHvN��Y[�v�W��Y��X�D�ת�t�l4)��2�߮�j�_��*W��{7�|��������������T�/8�9{_�Fn��a)B��}]Џv �� �Y|��O��c�/���Oz�Cn��S
=R��NI�H�,R�H�"��{�T�{n�H��
��ݞ.�F��6�x'�Zg�ř�p{��h��b_���/7X��=�n��^U�p�m�/7�Y&[c��w�صz�^���C��q��8&�k�`��?������c�w���VӁ �}?��;����W :c���*
� �<�mc��*��}ͯ�
Ș�`8�`���} �U�����`痨�'�g�Dp^"�-�r���mX
L)~S�=F�b L�X-���\<c�]���x0��P��ڿXU���{���/�G�U�ׄ$A�c�q���Y0�=�*��������>�����\C�#�������*�Ns�H����.��y�/��2�=���� 0ۋ�8W���7a�ذCڦ�)^U����l8�l�v�b��"���}]��e��x1o��2���h���e,���F*��''Q��f.*�Ū�5���\Jý��ll��h�ض���ĥn�!ƃ;�K5=JkT�?w����ҙ.���������5�������>~T.۵���x
<rY�?4�����`0���|��ars�'`\s��|d/�Һ�L�u�����rN�,ʽ�1����s梞��m*���D�v�4���_i��&M��eW��b�F叁���ӯ��m�6���	E��z�ד1� ۧ�&T$���@%��T3��/ɘ,��W��o��8�p����%���Ԭ= sJ؍��A��o���#�sj	�\�3�,>�=�u�w����+�n^����L��T٫8����;
���|���l�AX���ڮ� ���{m��� �vg��6w�N%;�/�r���s�	z��G{������va��w�I}�"�rͽT��}��������;ȏ&:W\���_~��h�H}z��Q|Զi}%0���,Li�ݏ5���k#vIc۶ϛ�����ՒA=��hI��w�P뗷<�{>���2f-36��;$}a�E���yk�������|�����$��{�w�,~����д�>����OR٣��r����烙/,i�-��?�|0�~X���C�� ���v���� ���=�gX�C@l�q�K�0q���B;q�.��i��C����5�������u���W�~L��J�[����%?Rxw�B�_��
�����B�Ҏ��5��+�����S0�*듋�H��TC���և���8���j�G��*�޼����΀ G��������ڿ�
��ԳL=c�U���?���,����8�e���~�GK0��8��1L��e�?T	*��}��u������0��Fn�����d����(�����Y�]��2zrs*�Q@���:W�>��=5��[��()'?����VY��L��wA�7�\��V�kP�+.y[���wy)?��=����?�-Q��nXߡ����p��>�U��Q�.�aR���%�H=��y������W^��w�k�E��y7�*����(y?{-�y�w�U�%�ѾÕ�W����|�f�ķ],���R��tƛ�Ӟ���˫��>yە�1u��D�b?���M�xX��ִ6!�G��������DgD9y��2���8�CB���P�6E�Cx"��oSA@P��o�d|��A�nLw��{C=�u\�1@���U�3�P����si�uq��._��ba=E}!u�g�z����9JKߚ^
�F�V�d�w��/S���<��l{�J?��OP��@�V`�&�`���*ճz��F��z����ӄ���~�o[h�}�+���Aja���{f]��U~�M�}����g�Qm>{�2�a�X�ƹ 4���Ut7�>qhD^T��4���\26��&U��x�o�t߁sT�k����=E|9���-��m.@�e%d�m�*���{E��J�k�7߬��wK�|/�!��G�o�`�kT��ޠ|g�Q���o�u�"󽍊^�FC�������{��{N�M��o3�煉��������d�������A������"߅T-�7��Ǫ�������)���u�� ��V�����|=A�S�n�W_n�O����|��}$.���m��xY�[To�WT�r���U�{^��`��|�|-��;M�����y"��*ߛ��)�G3�o�z�}��_'ߞ2�۔=��P�����M�)����˷������~;W���qվ�{���Xg�5����d�9<�����9�x�]����q%2�~���R�=s_��(�`���)�q�7��n]�_0�VX���m������B�����*�Z�����Ľ��7!��ͫ��j#��d�o�;�(��򑷓��.m���K�v�U���[H|�o�1��7<�^����-�R1��	m�m�{�17��-M���B����zf>B�s���ڠ�C��;���y�|K�
>���/�}�T�u�wxv]>3���B�]�ķf6u��s]�l�:�-I`�sn�������\w����� t[.�7��_ϭS�_��5j�� �a��c.J�3���xWi�\7������:���.�E����R�I3���hn��.�����:�ۅ���*�u�*�����W�����G��9.������Y)��t�����Ϩ�_#��|u��d]���n�E.�7���9�?��?Q�˟$����?R�GϪ�"���q�����E߿��3\��L/�����@=���.�(�u.�x]�����R������\�E���u����?E�[����K&�?V����O;��_��E�<�n{��m�7�1����ڲ2z��v5�0V�C<m�]��Rb���Ǜ��O{��G8�U���_�5km��U�	k���b�Z�>R��v�K��U����~�ƌm@l��V�aZ��4�Y{�`�]Ϙ�*��A	Z>b�cɈWX'�"�Fak����G�́�0vb�(�z�Z"fQ؆9
��
0?�=Ø�JUW�ۍ�d���:]�X�c�#���H���E�Ba�g)������3��\������s�<�&��^d1�U���>����jӺ�4��)��o���o���߻��� �5�������� ��R��-�����|]a����Y�����Ѓ�U�z�zq�B�����H\�v0W�UV����w���vZ�,	R{��\���*���?\�)=�C�W�̣���z��z6�;���ѳ�k����߽�v�zF۽Z��㯿Q�+1���4�QX���bd�hl�9ޡ@�mi�=!B�Z�vQ�7i3��1�!څ/�m�8�K�O-5)5V�¯����\kOCx��qu�,+�No���m�؏��WE0	7��80�M1��Tpa�/�A�+ͯ�ҧ��ǵ.��Z����k!�������5T/��n.���P�U-���"{�۩�MV���Jޗ��ϐ�^���[X� ��C�����$�x$&r%�H� ���.�{T�5a|�؄�Z��`f�e�.5�1&r%Xt�	�U綾�sT��F1�l�~�I1�s�xJV㣜��D0���V�י@�H󌍖Fϼg�Z~Z�p�6o�2��X:_ ���,~���	�����Ϛ ����Q����"�ؤ5�d�V+��V;�<�tGb��K~�pX���r�k=�W(}�~W�BH����/���ߍ_;����žݐ�ٟ����y�~o���Кn�	B�<�W���kϬ�x>@��Z�y@ӫ�?������Z������C^�7y"=�n�?v�ǏذCj�X�e4ݦ��+�S�}iQ+�}���q�Vk=z�WQ������,��n�J2�K8=���u�2hץ\���V��_S/B������Z�������`�����-Z�#R�`z���H�	v��ߧ�N4�2�ףW@��&���	�o���N�:�C�89�����ϐ����e�
�}/����ek�gQ�}]�V�_aj(�otLǗL�~��+�>�� v�p������[!C��
n4x�,��������{=C-��L8��Z �-K����r� g����_y<��Ǧ�J�y�!��h�������T+�(���}��b=u��O��5���:�S�l�Ftr������(�_,��
�iG~=Ѿq��A����=�Gc�%#�f�~I��p�wS?��T�J�6�kWV���$�t��mXe�~�~MU���B�����oP�]0�o�+��4t}v_4���0h���h�>0���Ǟ�4qᕖ��Cc�C�����v�8J���O��븟ڵ�Z�ە9:�:���V◹�?w��J��V�;n�tU����/U����0:�QX���P��	�`���ۍ�)i�SC�k? ���T|��c�[\�Q��wC<�����#~/���<�F���eQ���ϻ�H�}�D(�C��H/�Ńψq,���K��p B{W����(��
��Ō��ځ��Q}#M�\!��(�~���.�'�6�$��0"O
�?c�Ǟ�o.�Y�l��b�8���h?sQ�����v�Z��1>�d���X����f�8�_r���%HZ�e��8B_۵�֖�"����Dё�����1��6�Ew�|Z�<L	��w���Eť��7���Z������BBAϏ
;��4н߮)}���K�Kf*��3*�c@�l�sbY
74ҷj�xa9(:����&?�<�������*�rUoi?BGt��_l�³��w�rt��U���č�T���Oa�bC�E;������d<�e�hc�	������?�I�H�.�~����z��4�ѿu���hܿQ�^�G��/Q��M�jH�"7���g�i|�_]�q��������ڙ�)H�M�T�E��o�4�ϱ�>���׏�1�����~5���U�z���S?\m��E�y�oGK���z�3C������X;��<^��� Kq�����܎��S!�fq܃~�F@���ZAf�	�G+��c�@;�h�zmY��Qp�"g��7��:1>x�O�ﲼx]���)m1k�W�XpX?O;�.���H��	$�!��NL���Ξ;�"C�*�����yY��uz�JM�z/���S� �s��&U��kIL�h����1��A*1g{�)ʾ�3ON�n�,s�J��7y),ܒF��WWy�8G@m�����v�R�y�NA�B�I�1f�����U�)��Ш��ˇ�6q8�XX�W��՚�����gS3�h���A8B[�>!z�m��k�p�p|Uyt:��%�IH�)�N��жf�H@akE�mճM���p�u����xl��l�0"P_瀴	1���ap2������?�����W�O1_��c��yK��߷O�:�z��nFS�����j �z ���-Q"߉pz�?�%�W��V�Æp���!G{�#��4丆c�&�2�Rڱ���O?����;GM�I5�:<TO�Ӭ>}؂'Ćw.S�!7�*8��nC�8�B����XԗF�P��ݾ��l���@����9��p�yĢ`�t5JR\����I���4l�&���hյ���WFp��h��b�G�AoH8���Z�:�}GK��o�Au�|��؎f�*�����x��W�3���n�����ޓ?�3Y�'�;U�n>�{��	�7���[�Q�P/y������f��g���+�������*f�gnʍ�'@1�k]�,�Vޯ��ˁ��U2�e��7W��7��#��;��b.GY}�����	ܷ<�7���;m���<߭�و���,�~v��*���T���}g�p]���=���3������������kC�z/�5�4�����k/A3��<��%��nš8��H�Y��g=��YE�kwB߀����i��-��)f������0��ZύA���΂��I�1I��D��EnR=�:J�ޅ��p?���d�"V���zG���c.ʡg|0�_�А�K�w�_����6��z�V&��"��x�h�}�ɻh;�N�~��*9�{�-�W=D������ɱ�}/���[�[M���VJ}Ґ�:I�!��(xf]��a�V��z,�R��c/q�3p<�!st�R_�=�Y:�:���hc�`"�y���RO�,| � n�rk�`O>�O5�hCi%�Э�ǘ�C)c�D��j��ml���ʠoKf㧅a�]89�b�����<�ڢ&S %�j�rU�ؒ,K��F>��k�V����D_di�`z��$��s�8�/�}N�d�~MFh���Ƶ5�h��^������M���l&��+K��ռ�k,ݙ*q>�SzN�;o�)���(���Qz�sc���e�{9��jzR�`�"�G��6s��O�����2�ec��I*>�K��@s�Ut��Iڤ�����E�/п���?�ϯ��R��߱ �:��+*��\�j�+l��εM$8�2p���C�yK9�M�c�ډ��Bzuprq�y����XL������0�=2c���ڀ�|Q�����r?�g"(���T�3I�3`<Ė�@t8}���x&'�pS�G<��~z���"8Jw�3��}Mb�i�w��5�E�|wpqz�:���30Y��8�r�9a#M����䆺�m����5Cߍ��9�ٴ�<k���v��G�U)o��C]w?�N�'\`;5����)Hx��pm~_�N�oF��LY(�k�4�q#���[�&EվN�M�	�˿�K �	Rl�������X{�'�Ƣ�'���U�4xY#DM�:���Ry����s�����!OP��"��oӔ?�U>��+H�r�P��WOW�j�|����|��3My컵���t���؏R�Z-��^��?�l�K�),'�P`?�}�]~��~`�`Z��vN�i>V�u�J�ž��}_�hи�Z�E|E�Fj����}���F�׿�^s���*؄hg�7k�M��U���J�K���˓o(���`�\�C,H;1��!����i���Y�`?s�l�g�++pJ�X�*�g��[���f����?�ʟ?_�+�X��s=�_:��Hu��Ք?P{l���3��Z�7���Y�˟��,���)�g����(�ܫ*�왲���^������������M�w�*��G����0���g�.�]���e�d+�Z�ֿ[Az-�cx�P��ځ��Օ��c���q�?>�Пx�&�0�x|����Yu�㎙��ßd�e���@_	'@��gq�h�����fs��x�MQ�o��+�>���J�i���3b�w}Z{�3lNC��3_�'}��>���ץ>�'�k�O�Ч#�D���؂;R�V��J�����x]��O���%}�ٚB]��e���/�V����>��PJ�;��s,�]u���N��S�P��_I���]
�t�[:��c;�>��]��yR�wg�{�U�v	��F�z�^�Po��K����o�����?y 0�kT�#FE����!A0�d&���y@P�h ��+VT��j��ՠ�������>���X�)R/m��}��k�9�̙I�����G�a����گ��^k�}���cr��O�������+}D�F��x.�y$�d�%�����������a�>��}�r�RB�I�㯿n��[6������Q|iN|��vr�9���fw���R�ߦ+���f����V��k�:~Z���1��^%_Vs�\ �m3�l�_n;�x�y��+(z3B_7ZW�[x��'�x���:Lj�OU_Ԧ���w��G:��·2vi��O-�B犗�Y�|m���{q\��}��&93�M6����H	���kxƮ=d��?c�̤�]��|���ô������s�*�&���v��躄��h�0E8Č5b	�ٓŘv&��vIg����N񦇌Nq����C�t�*�C���]&�����OU�~t�O�^���7�9�lu�ϿQ̇����I�KS��d�
���J/���F�Y�!g�$�{�7T�������}���u�t=q]a�u����u�)��[S7�n�������uk�0��1y��k��U���(����k؀��z�?�p��)�X#�w�w�C��C7Ww�+�9;<��5*cWe�9{z��|�yR݌�p.�UO�m9gktF�#9\�\�?�o�qbR��&������,G��b�z�����h�C�w��D�!7G߂��9��r����a;O�T�~ �K0�CB/J*OM�Ґ�8;�u�,ҵY��8��&����J�ͤ���b��Y���V��~�z{�8o�Q5<]VոI�����"��0���!i��"���(�&['�?#�������	Mz-ֿT�$�`��!�y��dҚ72*&�����,��@���|���}�:��q��FyT�k�G)�U�ۣdh�<���Ո�߰^�9��?7DC0;���{�i�^�KUR	���}�V/z�4N���5����ʑ�b�2���%k�o�Q)���o�Fd욟T���U�"������#s�.ay�L=i�S��i���gx1���'�h��{s��/`Zfh�4����ᷔ����Ts���"�v&��_YC2��3VOoX5H��9�u��R:��R���=\��}륊���y��<"f&a�����-����rKּ}�"O/s�G��~��3+����r�Ћ�߈w��^�N�l�Ѿ]&a��o�����Z<����h-\'~�Gv���#�b�z}�Q������V���}�n��Kz��(�k:�D��j�>�7�|y ��5o��|?݇�%aB�j�M�0�������x�B�A�!�"̶��~ʯ �u,�"��R�yM��(_�S�qnY����~ӏ�ҩܡ�ȟ!~^$�a�=Lu��y�2���2�y���ly9��P�f:1p �-�ο-��'�����a���yc��� �㟵q⟍��������\ؼr���/�0n	�y�Gk)�Y;��g��������5��!�}Wv0�
&,�$�zJ�AS�."���0���u�C��+Jx�:��%N�i�����(ǅ1q�����֚�x�:Ӻ�6N�f5����I^�0�f�)���9�c�G�o����й�w*4�+�ɥ����������q��ח�:��'Hm�v�;�vփ�P:wu���M����Zc|*����n�>���ևһ��������z����g�_[m����e�rO�cT��\kU���˶��k�������*�z�N�������W�9�z�N{y��a��/לh�U����w�[Wmo���>�� �wl⯭C�{Ue������(�*R���!*��4Γ�h҇əI��G������!/�z1�9Hs��m�8�(���؜��m+�lkn���@ض�-����m�S��6N�i�c��?���ͺ#6n��Nc�!��@���F�붟X�����S��~�F��[���k��9���I�6@�Vc��,��
�Ik{���N6X���v
[[��'^q� a��5�rp��B?�7O�;.�k����]1��u\X�w��Xާ�0�ȵw�D�g����_Y��'�s��I����e�*���>u�m��l������O㵌����g����6��6�x���7�F�n
3��ôaE���B�����~k�x-ɼ_��6ٿ�2^R�D������:y@����)V��n���7ۍ��#&�2�-��?n3	����޺����C3����">�듲��"N�^\"4��O���.g��v_��6>�n����ͻ��ܽ�[7���k����o5ltg�ݷJ�l��3�^_)�����'�?]�����?+��?w��U�?����?]���s�s����8���_:����?�q�6S�s�U�?��g�)��u��g�}��u��j����b�ޯy����7A&�/���5[=�PU��菒�;�i�郴�~,\A=yy��W)zA��n�4�����������a�w����7ݿ<6n����%�ܒx����N$^	�)2Y����4*N�q
'2D�Z�StQ/w��iW�Z,�����Y�c�6�v���n���uq��n
[��+�����~R�WO�ĉ'2��z����r�#=cW�a���1d?���8��j��S�w�eH��B�ca�|x��D*&h��������/ƶ�o[�OS��T*6k��g���/n5����~Le����*�܏w��Vl�Wv_$�Mޒ�������������-����b`�e���jӭ�i!������������G����7���q��i�������{~f��~���D��WjO��2{�Ǟh'�>2��'[�>�p��ɂ�ALo5bEh�e7�&��`��dv9}��e���X�nN�>yI_��>�>)�����Fy��Jm�>���$��<����`�'�=4���Ko�յ�����g�>�"l\��Nl}R�7�O��2��dts\�^�`"��n�}��}��l?�)a�З�<�}�m�ž�ӭ�e>�}?��}�|��}���/mߝf�>�k/�O�Fy\�r��ݩ�|Z�Ѿ��о�-�]�l���u��S[�t%�u�O��46�~,`��?����Ӧ������;��O��?��	� �����\�<�+����r�v��'�5Z�'�-5Jl��_�>�������iq�'��7�����~���o��Wy�>Y�d�_:����x듪���Onm���e�~��b}��h��ĥ�O�����M�&�_���_�����޾�E>c�,��6��Zu+l0����A���<��+��K���f�u�'��7�ƿ�D��T��+���������/Z�������8��
�ړl:|E�3�h��O32����|�U��,�$��n�j������zf�z��.
O6��������e��om��k���IC�i�)�9}��M���W[�g����kП�:�el�7��
���Hp^u��/@�k:e�狩*ę��d��������ϩ���ХFy9뭓e��Ebb�ԙ��I�g�]ꊱ����B�2��J0���	�i'x�x�a���ǥ���䦈��p�'b9?��v	��F��bf�F��?��؜~��{~xrG"��}�e{����8�_��/���Ŷ��=���2��n��8�_뾴i��U����7�՝�i��՘��\�-�]��{�#����M��|rE�������q~��Kb�~���������~sq�z������u5��K�9���<?�k��m�Lj�e�uS�W|~x��X���6������;?�[dYO-Yb�h��z��+����?�6�l:C��U�!�8BU~�;��͓��`�H_2�&�xi�9^�n�����Ksn���kM��&�x鈊���xɵ�����
G�⥫�P���'���2n�L�����d�P��)⥼�d����Y��v�������/��sW�Q����S�G�y�I�/,(����v��|��Wnƚ���6����K�k��b����c��-�F����m�Pi=,�����u���#��ů����o�#Q|�c�َ8��q��7���7ZU.6>�m�%>�]�_o^��0��U����_:>k����������7�h|�]�/0���������\5����|�c|���^�"c���W�w�|���c��C��S����L��ϋ��~Ui�B�x�|�_o=���m=���Hﴱ�.���Z�?9_\4/v\"7ǥ`A̸�;_��:��-�o�?UF���/������8�a����gn}��nکx3�}� ���,\LoP�!�i��㣾+��'5��P�`� ��na���ø�w�O�~�������"z���oG*���,1�V�%���� v�,���#��];>�^�W"��/G�W�~�|�^��Һ5��=�O���T�� E�K�|�z���&���DBc껜���r��w3)!�̹��������L�}����>���o^	;�y�E��?��/�5�����Oz�/���V�ֹJ뻚d"_�T��z��:���Ij�3�:0��g���~�n_;�$qo���rH3e�/�'集6 ����7�!�������*z/�^gG;�s�K��F�#�N���0�o`��<4���BgF�N���|C��S]��8��Vz_����}7��qN�] �[����K/���C���2�Y�_2G�i�c_��#u��.��I)i����}+?�1O��k>�C���%��X��!j�U��������������ǥ��[�6uN��٢�3*��B�ק���l�8���0BJ�L�4Z�����oӯ�5�����-�G?�L�ߏŰ�un�����*GΘC�껣�����\�Y�1���"ǿ��Q9B5�E�ax��m�83.�ё���9IӰt8��>c�yG�3����0�oR�#���u;|?�u$c��nM���e������g�}t�����H����H}���YB��Vs�꘳��U���Ez�~ӖC���>-%�s�Q�q�3;!g���#㵄��F�܌�ۈ�D�pv����ug�K̜���ӌS���f�(��4#���?"?�s8(�~%��+(K?eqv��A�J��yl��0n�:sGU_4C�q�z�#q�OD<�'��r�mmb���	�w� ��D��X��6��-�t�|�Q�	��'��o��O�C�ڧ+K��\�IU:f�F���z�Z�ꘞ����A�Xu���x��H�d;�:7}	�_&.Φ�a�8�#�P7�S���!BR0�O�!�(a;E�z��w\Kqjso���%(�P1���� g��ŉηĀ)^C��הF"z��\��d��u�."�{8��ڏ���.(GZ�~	�pRג7m�����~l�����~�Y�h{_��c�I\��Ѣm։^n(�}%M�n�0��zg����Q]��&������x�ꨁm��0��������Tz�+�TԪ~ӯ�LBT4[)Yu��v�3T��awLP�Q���{�s���1r&�!���7Xr����7J�2k�4�,�$�Հ^aK�`��;;R��.�(qZ늣yJ! ��7Rѽ_��A7�ޕ�~� Uc���<�Ҏ����ш�4c!�%9�UN����E���g���RU)��h��b�h�s��Bb�C��ؖL9��Į�-��sJ�FKu��v�7��f|��<o�5RJ}�n�t�����IJ2����?�;ބIM§�6�������ˁ��r���y�o�T,�G;���Ls^x���wgǟ>������g"�-t�w�D�:/sGZ�X�a�S��z��=�����#T�O��?�V֙V����̞��ޙ��C����,��C���ຂ�y�EzPX�M1��#|���}�Z�E�+r�MS�<�ܡOai+�1c�Y[���X����L�v&����x�^*1�?�dc�9�����:tcx�s��K/ҴW&�!�����軺���>M�����>��\�re�Bf��q"��eD��H��)�If��ӗ4��)�?.D�2�+2s
e�YQ4��s����������M���؆���B���U�:*4,����<�� �����c3�&_�э��!�C�Bs:S���CD��ǝ��i����'˧_�>��@��=2��Ww4f���f�8g��&�������̑���|!���ƾ
��HG�o1�=_R���ʨ&�HM��A��(�N��t[�t��iQ!�)�r��'iB�I�s�]�N�1�#, ��~-t���Ia�u^��ٱ�gP���Sr)o�23�p�jBU[�Z�x���s�о�����o��U�;ʰv��ڌ�*�*%ՏuR��J:�I��"��V<`�{i�a���gRXxx$S�莯3iBq����Z�A�0��fb�IՑ��x�G����7�sg;���f�Mр������*����F��5��+�����uD��m�+6�=0�t��:&�j7敍r���c��y��׈ʏM�z�W�$�/�w���4�����s(�ts�O���E�gk��j��	�>72�fG5Z�X2����r�<"+��Q�ET�W�1?�w8_jt���cºgj�'d1�K��x����W|��q\9�m*�'L���R�B*�Rc���:dc�K�Wy����%�}{廲��;D	�R	G��K��K�3�#�R�"��B� ��䪩��dQ�ˢTԷ����	񠶤G
�/�ĕ�b?%Hq���^��$�8s����(Ǚ+�P{_���|��$^��)*mbF>>g��K�x�'�x���^�����!�iH|S�-r�$|G7˚t�9RO������5�Y�H���������Ksr�z�Je>�d7�cwS�gW"�
��i(q#�)�ҋP�W>�#��b�n���|�PϾ$9BB=�2�.�� ����^.�c!��,~�㰁��[}/��u���s�k�W?˗���kh�2ve��:��Hel[u�2t���J���'��a9��}E�T�~�1�KE���&�8A�.�A�k�j.bbf����>a<7;��IX�cɡ����'�2a�ۏ������B�.'��Q�e��/�������t/�"�8eL�*�����3C�q�p��e�����/��t�8��$����A�|U�u@ޕ�u��������p9o���p�D̨��v�H��&vl�����A�ȆZ":'��NȢ[��U� E\�0����+x�
-����^�?���uQ�sS���"lR���Sg$�� f�+��ɑ5ZL��ir�N�;F9ć][e� �| �����Yto�7:�9�+�DΥ�!�,k*"�BDw�4q�B\��q|DD����Nq��L����P�/��kdq(�6�M���K	5���F�C�	i��ڍ�吤�%SC���:;�#}���y^��><U/J#	����m�#�/�p
m���0�uA��q�_ʟ��R�t��q�Oaߢ��Y:Ӏ���JiV0��+���%=��̰ơ�0��U��՝\����zp&�zZ�i�J��#� 4OҜi�ap�)p��ZG���U�EǣEd�����6#�%'���W���;g�Sؐg��􄇒�=<Dg�;����i��4���9��
R�@J�v�j�[w�\� 6k�4���*��\(���bk+ټ����$�cf��)g	In���}�w-�:����Б�дx���Pz�i��WK����zy<��,n�uqS����+i�3����m��+��-��rF��N�/����RV�M��B�y8q
���.M��L}�M�i_���5�
��(b��M{�v+�:&R�s�}�Q�r�M�E���B�k*��KUx=��(�3,B��'Z��e?�ܪ�d�����8嶜��?������@�[�\,�������	�SRsh3�y�_
T�9����Rq̬s.f�K�HE�:2�z���>4�����Q��)ԴOP���D�y(�CgǞ�N�����2E�xwDKS{q�}Ʒ(����|���\���;oBVd�Ou������V\F��'i�0�&�*+�|���Q��z.�/��ZW�2G�/r��<��s�!����S�l.�FO���P9˛����h�7�B��#��ʲJ]M^���m���F���j��u����Y�UѼ:�.�X�iC�Z�����+�B�h�5��˖�7��
4��=���_��l�8�~��ъ�����>\ϩ*/�y]��޶1v�����!Ԅʬ�����ɷ�_�
5��1��U
�GM>����i�Y�AW�Ǒ[9�x��R�rץ^����ya_���S�Z�i�j�2�r���n�)�1ڵ�'�T7��xT�.���	'�it檫����(��.ԋCR8�3���(�D*��>=��`$Z0�?|4|zAO��P����?mv$����Hd+>ݸ>6K��p?��i�g3>��9���;s�W��z�+�6�E{��r�ѮC>|ZvUHZ�\�͟n|z�ѐ��g=���J܏����h;p!���?>���^ ?�t��6|�W�i[�G�Y�k����x=�=^G0ׅ ���'��Tz4_�kW�pԹ|>��bb��������%��?��[Z���]�JE5ֆA�V����l�W��j�.�Z���!ȶ2�#Z��t�+r��mF��)t�����Kal�Z�������K/��t��e��h6/�&j�3/,�pL�D����Vb�TZ�m�����Z�m��]e��� �Q���܊2c��ŘK/�L2��o�X���Z������,�Ř�pe��]���ss�)�����|�s�V+�9ۍ�l2ɘ��х���iu��Eƌ:�1k���j�t��J���1O�?,��Xs�K�Ul�%��CX��g�E.w�/�l VH�k���&K���oT	"�5�]�PI �h��O*�e\�&]�Y'oK���`�.�TxP3�
�nL� ]
��J�J�-+3*�^�t-�	E��{�rk{y��eP�yV��g"rq��Znl�1��Ԁ��2Kg:���@�*b��C`�g�����sy��ee3�7Df`�g�fT���ƣ�����͵~�W�G�	���֤���f.#��=]s{��jYڢ2�z��R	�Ԥ��	Z�?��p{�J{�U��ܞVuSIkn}=FH�I�8MA�C
�^T����� ��,�������|2�uF.
^�`���v���ҥj��k0��:6�E~�r����a��wA��r�d�v}��9W:�̭t̻�l�FZ[���CY�Y���=��D���^DI4��*hX<�0�UW�I���W:��[s��Zu�@��f��˭;�\���U:f���?36�<�BL����<^�c�Icǒ�4�nY����;A��H�=~~�d�R�G����/���_n&-:���y����-f!^�淚���huH~��C����hݾL;b�}!	����K�4�'�?���Uv�D���N��1~��m�2'��6^)����xy^��y��CM�Kg�)�5S��A�"�x�&Ԑ0#X`͋��o��5�7���m�0.��S���Ѹ�WTO̫��B���մ�_ɼys�]������#���?�.�Ҝ;.8?x=VT��� �?/�v����W�?��������EL�8D�nj��AǕz�yrͯۻx��*_��Cp�kF
�����}u�lM�''��[�Vy�V�g>[H�>|����������g�����n|���O>5��0��.N��_~��~*������o�"�˕�_{�4N��'�����~��u�c.�s�b�Fү4A�Ԇ���0���9��E>�ϣ�}ёh��;7�[����;G��B}ƽ�G![��O�P��c�V=#�Z�R�],Y�3V:ƍs/���H�^�tд�%W�<��R1�g\��-.���ІM��)�K�<M���Hd1>=6�[������Ч9Aڞi�C����d�{,�c��XNW]+[��h|bhD���
��ȩ���7�\�����G"����C���N{2}�"�￳O;� ��P��a��~?����R�B�
��U�������`�X@+
���)�%��Ҁ��cWD��uY�/�7��CS&y#+:��NVò�=�z5�Z惀�*��W�4��\�nr��&/�q�d���误w\�ȳM�n/%�Iע%��2}�I�vY��m;=y�{�ȶS4m�H����D�`�sr"����!s�{\$�	x�*���o��������"�J#�0g<�'�$�,�x �:RӎG���V^�l�{�^�!�!�<��d�kb$2�,N��;��ŗE"�]�t�OC�ۀn`����� �C�ע�����nn�><��*C?���G�n��LM[�����  VSgB���j`%p0�	�|�xxx�5������b�&�b7`x��Z��V�F~�f��r�3��K�`��u�Et�^��[�j�Q�N���P>0�U�r�9�J`1��W�"?p�(ppd�� g S�����y��h>A.�p'p��<�t�����VzP������?0�-�(0�khw�88X	\<
\\�=�,C�g�}��ぇ���P3�� W? ��F��(��<��Z!�l���&�����ۀGoC���
�:��3�G����v�݁��P/���މ���܅�v��r5��Y�� ~,^���B��b��nȋp���r���m�ЛsP�z�X�|�C�W����=���O��.�r�C?�Y����ɛ��� �w>���7�o4����C.���M��o���`��~��@�����&�ݏa܀�����"�J`0�	�x }��C� �ꧠ��m@:y ���4��}��~;�J��F>��� 0�Y؋�P�s� n���.�zz��v� ?p�g`��0��b��6���}��w�]���xt�<��p��hp�+���~ >`1�x ��}r�!��^G��M����
�z� ܶ|������Y���n�wC������m��}��x�ҁY3 ��ނ�s�^`1p5�(�Y��>�=�(ݿ�����h7�X	�C�{���/w�< ��	��f]�i�������7�!�Q�&`�;�� �<
�	��i '������!��	�M�N�π��g�� f]�im���W���� C���M�������(x�)0k���ԃ����J�3���M��w�}����G��?G�K5m%p2���J`�/�X	�l��@~�����=�!?bp������C<�����a�x�����[fMԴ����y��*�و�B�+�����;����?D~���I��C�d`���73!?�< |x�+`�e��W�d���D~�����&��x+� ��Q����ɚ�6p2����9�����������? �� f]�i�����>�'�x1�yZRkf��#��u!^�)�蛠�#"�'-=�4={fƈim�5gM��2�Z��Ҋ��֑t�cf����ץ�Oِ�|������?gD0��vC�Rp�;;)"�������������i��*w�f$���h�v�(7uC����Q���^Q����WN����\�;J�=;i�-7��K���B9�Q��P�������3��s���央M)G9��n�A鋑^�t���B�kev��vһ��C�m�ڡ��� �UlL�79��e#�� f�Hv�G�rw�?m�}�Hn�8Hզu`�9�A����}wؗG����׳dz�\�&9� �t���� �ў�69�`��7��52�|��w�B��?�=�7jj��ӻ�*0^E4^5r��@`��;�/�ED���z��r| ݉�qq�O�N�������|>ͪ�&��hڱ����'��Ӆ�s�s܏��sҳ�S�M�NJޔ�]`h�(/���h���ܬ��MH?��d-�G�gA�Щ{A��r��c��O���:��7�Q����BҺqd*�������{�ӳ7���;6����R���vhQ���a�{����E�y鹅�p"G!)W�$�$��P����X����Φ�b����M�#���c}��2��S�֦��e��{�7뿥����s�w�5�'Hoú�y!'*
�!�}���#����@���;� g��pJ}�I>%$�B�Oɧ@ʧ%y��
G���$��لz�".��z��!�7צ�%Wɮ��y|���((dCrIz����t��T�>����\��U��(�C�q�9���l=��i��3@ϳ�}���
�ՠ/���z��N�[m���ˆ��A��B?���a�O6��A��/���b��m�C��i�z�3����z6������� }��'�W��B��3"�}>�@��L�B�
u��E�}L���[`P0c�qS1=�4�+�?}W�� �LL����v��_�B�Y��O�$yǔ�O�?��;�eJF������g��P}1�$+;�Ov�o�s#1�kfE"[�z�X�� ���z%��f��!����_h��}�,���!�N��әD"�JϜ���;��.�
a��㕃�	�{������*�g��Mߚ��L���"q��G�`�i�?�Aa�?�]6��A_7Ǧ�\������}N���}��!�w���>b7��z��o-g��o��~��t��ԯ٤]d�+����L3�'=_�T��+�D�P@�Cqz~��ӳ���(���N\��C������#B�?��[l�O��O`t��!������z���N.?mވ"�!�΢
?�>D�O��K���ߩ��R����O�U��o2�I[8�t"�����_��8�F��]B��8��rh��:����I�+D8H~=�d�o�?��=%6r+��-)eQR� '%5�.A�ǋz2+#�?p{�����t�GNc@��]U����4�BO��M�E�)"�u)����!�qs\g7�g"fMٓl���OƄټ�l����w�^H�92.��Q;�H�F����hЎ��xҔ彊�*E"�X1���p���Ql믨���3-(�;u��smzoRʲT[=5�G���ռ>�Ӿ��,,�o���Q^f��O���՘�T?=/�@_�۟��{�Rf�$��x8rG� �)��g�}��Gy(/��I}��+�����t�03�є�Y���U�w!��r��׊�m��죔������F���d�-�D"�g{�+����.���%���	���-�F�o5�6���,��"��I����q���<7���/�/$�Ak?�y͎�h�A��So7���SDX�1E�a��6�ޛ��J�ŋ���_����tG���JF���ԥ��?si$"e\C�o}�R�?�K�E�q�'[+����r�}��S����?�ۿ,+���b� �lr�Y����`���?�~1�.4�%����r�������ۙ\*�^i��!9�������z=�i-ͣ�T�~���tG�2�h׭�[ʿ�7��q�9M����V��$9l��G��-�ȣ� ��+6$�OIn�U��c�s��������t^d���������8-{2�>1\�q
��@|,�_q��?��:-�����0_�c�yɷ	��<���i/���?NG��9<�8�B�k�G"�q��c�89c�i1��X��g�>3�Si�8m!��x����ue�8���6�/%B]t>}�ʘq�
�Ɖ�_V�����"$�&��/�V�%�[�G�*['/���?N[�����|�WE"��ӓ�q*��T,�v��\g�7�SQ�8#��;'/�m�q��\�_�~.����O�_w��w��l������;/�T,l�w%�3�_f����ߺ�X}������A��>�>�s������X�yy����i�������|�����������x �ww<N���wO�>f�{���H�z�X��k���7������U�96��C�ۼ��O�/�\�V�+e=����Fa�ߋ�^G�E$1_V!�?��o�ꛌ�8�X���^C�� ��5����]����Xw��zI�2*����:�Qs���;��G˦�ǋ·�m��g�_�&^�b��31�J����}D"��Ja,��_������y����C��c�<��G1��m�x�������|������o���/�:��e��*��Gc��b�k�}�b���z�+l����;6t:ߓoC? �T�'��Y�4~�����"B��gr4�~��$�P��4�['����ij��3�[Ur�B"�>Hr�d�G��G��w$���o}
���k�K���b�|���~��]�r1�6"̧�_��>9y�A������f$B2��'zJL�9�/����s��e�B1{����?�1�|���BHO{,9K>���R֧��������Ӷ��3�����r*:y蒑��8� ҏ<�_�/��E��H�Șg!��	�'#}�u�1�1�^I���>���M�sac��/��'('ҧ%H?@��A�$cz���H_�5��+����C���OF���W�����m��oB�S�����!=Ϙ������ ����<Az�y��a�t:wd+�[��[�G����>�J_e��y��`��7!��W�Æ�#�&��bL/7��s��G�^�8�����A���H?˘^e�?�_LоJ������Q�����_=���z��z���>�	~��]��#=�	~ު�k�G��Oį�(үHP~���v��7�����B��bjXo%ҷ �kJo��C��\��M�-��S�O�s}=�FO߉���>ϔ>[O?���H�1�W����O�߬q���yϖm�Ƚ�����@�GI�����A��O=�|ה����#��oE"�M�s��Gz=ҟ5��-��H?�=��)����G��oG"�2�?�(���ğ���>'Az%�[�N窢�D����g��iE��0����Y~�������#����.��?��?ҷ<��;U����G�#���o:o����?W�����KV��D�M;"�"c����w�>������M���?ҏ"�jc�J��Gz�|>LϿ :�H��B��c`*�^e�_�矌��t������J_h�?��B|�nB��	�w"�������t�����Ot����'#���t.���t^��D�G��D�G�݉���;_�oߏr�x���i�!������@z�i����G�_�?����/��p�>���o�^$r�1= �E�����3����߿�������������U�+1�^3=�q����0�H�w�K<����$�|��Y�:�����R��>ʒ��f�s��"����^\>��A��?C�z��:�����Y���Y�������>�0�3{�L�7���+Rg�U}_Dd���?����~���������[�������cK^���AƧw1�c|��#���ʟ#־�8�q
c)��z��kd|�q�>��?b��q���q��R������2>��4�.�}��1~���е\?�8�)�����3�e|��i�]���c���3ơws����0�2.`�g\θ��AƧw1�c|��#�������1Na,e\�Xϸ�q-ヌO3�b����G��1����1Na,e\�Xϸ�q-ヌO3�b����G��1���g�8���qc=�rƵ�2>͸�q�{�1~�8���g�8���qc=�rƵ�2>͸�q�{�1~�8t=��8�q
c)��z��kd|�q�>��?b��q���q��R������2>��4�.�}��1~���Ѝ\?�8�)�����3�e����}VEW��q	�C�]-��q�c�?b|������k$�0�䫈�_�wmQѕ�ܪڰ/�����
��'\1�K&�q��^�&W6�\��P@b����C�	����p��}I�[w��`�6��҇�C��\���tS�����"F�j�	��}B�V�_���ݮ�K��i����=Ս�@�N�v��2��^Z�p57աjH�'k�%��ڄ:�xS�W�G���U��?Ɍ9�T�==sbȯ�)
w7糮khO�3��*�Z�(t��ϯ���F��[�K���*�Z��kr��u�Bӗ���O�95����יqf�����g_�u��
;����e��j��'��T�}��j]�P��g�M~zg�D�;�:X�Zߪ?��-�[�ͨ�_�eZ�vK���f�y�>��[mɯ��
O��[����T-H2��g����ݒ���$n�4�Z�VK��I&|�b3�U����j@�S�}'ɖ�z��C~���?��op�U�c��� ���5���+����<j�D�W��c����1�2����.C~����W�(����M��[�+��En�9����T��]ce���f~��}���Y�*�Ez�O1�m���?'����D�����l�L�Ӿ���jN�S��#2���ן�/��m2�������o�驺?2Ӈ�~�L��3}����4�ޛ�'�v�L��g3}�nw����=5�O�����&z�n���L�^�����L?U�3f�i��0ӳl�1R����n�-:�M�3l��h��wf��14�e��׈�>,�T�'�_�,;��2.���c�_�t���Q~��j��:V��s9�r����Z�~�ġ�.��8�O�Ї$���y�����L��v��8�`��Du5����^gz����[��A�[�����3�ڞ�U����Ó%��B�N�/gl�}�&0�a�Ogz��>K�Gj���v`~��<]q�Mq��q��š?�,�|�ٞ[����j]��۷����W2�}��u���1]���1=-E���\���\����z��d����*���S�t��?��˙����0}�պ_�?�)��}�0�_c��P/�/�^Οġ�"��d�� _K��O/���J>L��tߴI�����g�b�HK�n�G�����b��A��2]�S�y�w[����3fI�z�LO��>�C?����5�Z>�6Ğ\��Cd;{�,���W1}�<3�$N9����Ö!�^a����6=������q�6��o��N�����t���5�wX�ġ���\����,��H�ϱг��Xܒ;��0S�����)C��-N9�C���r{Ը�š����i�=6t3�5~k��8p�P��#�q��"�oJk�l��9�z����{�w0�8�I��֭�w�{5�?�!ƿ�3�y�x����-��������~���?��w`�0ٯ4��~p����rz~-����uL�8*���m������[&Ɇ����a�g�����*�'0��kΕ�?3��4I�|G�+9_�����1��`z׳�^m�T0�����V�_��8L����Xo�`�&���JIWvkk��|^c�|�ۘ��L���'�$n?�Z�����y��Ɲ�3
��Y����$������z��'���d֓M'��e��.�?W�����;��/��y��0��ey��q�p.g�dT��;����}�Obz�(3}�p��>K��1�%��q�rU+�ҷ��>����L��=/����3/����X�p��>e��J���������yz����8�!��a_~��=,�_ez-��y�m� ӷ���0�6�;~�����s�.s;����p��;�^cz&�w���N�����{Ob�b��)�m����L�ai�%#�>|$�պ`�k�)�L�0��RYa;���8Ϭ?O0���~&��a9���L~�y>���W^+�`�1U���}!�G������'�_��n�>���r~����.��y�޵f�g�j$��|���ey�=�w�����k�s9}�r�r�I~v{�I��-�9LϵЯLg9[滓��,�3�����W3}���oN'��U��;����O���1��1y���w��`��"��1�[z��<(�ǋ穮��ΎW��.`�r��>�ez��ߐ���g)�,~���-�� �c���rv��j��%�����wX���S3�'���-�I��L�)�Y��xc�۾f�3��c�ٯݕ)ۣY�� �Z���r*^2���Lϳ���3���.�E�r��N���-��d�"�\i^�fz��h&92�w����O�o��n����8��П�z������0}+���K������Ͽ2��+�z{��鴴3�T.?Ӭ�����Q�^p�}�o>U�?Ʋ�X��Y�s�*��Ov�C\N�eܷ1�%^z���-�������2�~;�.>?t��o�-���\�wx4����C��b��y��˧�4���/�r�6�{�����O����[�6��=���w�gz>�S�ϲo�9Y���-�4�����=�e�ML�q�Y�2��=y�;ȇ��y���o1���^�����e��?P�s ���e�.�o�_S�g�۲�~�j���Dޫ���Ng;o��M�_1���U�S�{���R��L���y7���K������5�ܾ8�~O��m˺������n��|;�.����
.��y�<�k�?��� ��x�����~�ە�o�rr��*���/s9;��|7�cz7������ط�3x��t5�r�����W6�RE/0�Qә�] �*N�2=��l���3�x�d���ˣL��y��Y�ϐ�鱌�K���_��Z{���-��	ӻ-�|��.��ٲ��Z��2}��^=�:[���R�u��m�G�)�~�����#�~����l�x٣��tm��>����Y�s �^�������u�?��o��O>��e��u��L��t�~Nbz�Ps����]��z=�3��w1��g�~�X�����x��#b�C3���߸���u��x�r������߫�������1=�׃c�~�k,q�L�ղN�?�~�ne�~�3���ߪ#��V�ٿ?����G�8�~�A��Qr8ۼ~����,�O:���O�<۾��0?������ҞyqʩW�X�m?��y=��.��2�e�<�ole�N��������j�x�#�ws����DT;�ުq6J�g�E�cF���Tޫ�S�2]K6��|.��"��Q�X��l^�{��
�:t���!˯d��o�O8��<�+����/���z��7��3�n~.���ϙ?�R���_x@ޫ}�R���j^GT���HyV3�X��<^L׾%�2������O1?�_�#�R���a��2�7O2�������:_T�Y����4S;�1=��|nO'ӧ�I�T�O���W=���t������[-�����_X���2���G=��ӹ�^����j?�g��-�Ӻ5i4���pܻp4�/Y����WZ⽕�����8�������fz���+u��/L��6�ɧ;���l�}{�;��a���L�������1�������3y^���0N�?g�<ޘ����qH?Rc�#��pe��icd9�`��3}��z's9[-zR��l=�lW�):ۇY�7��د�qy��������ci�/�?�����'����rR�=����ɖ}������6|�T���[y}����L�����'�s���!0�����h������{cy}dݏ�r�/1����؎��Pϳ�e���D�S|�GY�_��;xB<�t7ӯ�j^�,cz7�7���鹳���~�7Ӳ����=����#;�u���C���m�Ϡ�oD��'�z~G����Mⷙ4�]9��-��eL�m�q9�<��=Ks���3�g��`W����X�q}�뭰Ի��9��a7�����Y��.��6���3=��%u<��L�x�|9�����-�9�|ɿ�X��]��c~����c����Y�Z-���RN����:.��o�簛����~#�Q����W��E.?�"ϟ27t*���;-���c�d�������B���Ɏ[�]�q���w1}�����~�b?���3���}�fz���g�����aS��>e��wj�N��Ǒ��z�u��ߗ�ǹ���������Y��̿��/������L_���S����v����������_�>b�y�x��]�����3ry�����sY�O��Bv�e�_c�_��yl?�y�z��sչ� �[,q�7���=�6��[�p9]�-�վ�/������C.g���az���9ӷ[���9����W��㘾��:k&�k,ql�鿲��1��bIW������1[�y��!�wX����j' ���O��������EEu��Wz�����
A������2�qr�ElO,r�:�W����^3�_���-�����<���\�E�?����̿����2�W|.�}�gzM����۸�lK���~�����sV��%�2}�e���t7D��gz/�C�/w�x��<=��-�~W�����}�|��s�&�iu�P0���eu�̢y��e�+��5�'�ih
�<��Psu����5Ru��_���׺���?�v�[�:s���'L�b�T{���o�=�P`�&���77�D�]u����Z��zk]u˜.���	��E--ћ�@ ��Ek��%����Mi�WG�Q�k=>O��n�k��RbP�b^Ie�եUs�*��Ω��0yJ�M�����>pVx]�z���\+�BM�=���
W���ER�h��._�����Z�L�x�W�si���x]��V\T��-�6���MA�!����a��)�W0�Y��2�	�>�iq���F��߈B��ʅ�!�G\5ʞ��p�_�..қ&���UT6<.w����Eo�BM^���e�E�T�V��m
��>�j��JX�ծ�&����$���j�gI�@�x<R��,�f���ɔ�}��R��{c�E��@,u~�?`��2�Ѿ�R��e�\��zm�]�o���mI(��LB���^D�q4{���&��oS�H#yd��i��3M�'�iq�N��0mR��8uL˻L#����>.�����NC���Uupes�i=i��Q}�z�u�+Z�*���[@u�LXo7Or+):{�	[��ɇ�FJpep�a�2��``P��6 1L�r����P�M�.	 �%s��)�[�>B]C��&�����Zh��7�)�]Vj��"�}m���깥��K*�+
�K�f��1(E0��p��P��0~�j�Ẇ*��C#�xV��Y0[hz����*���i�kY�/M��	�&\��E��c�jM���udD��(�pe�S��V�kj�][u���B%愽^�[L�P*ZAK������,�A�a^��sag{B�~0xB(��?�j�S�Ȯ6�VODqY����ni1
�?�x=�j� $�G�hB����Ksb-��_=Q���I_�7���*���+	���JOs����穷��<�P���.4P�*���-�s������VW{��rw����	7����-�7�\jԊ:2�CR�tM�+����RP��MA�%�����=�V�o%��J�<^w��Z����P��-ǈQ��e�����&Y��IvM��A����k�1sD&�I�^���U��>��D�&�,wCj��BUd��!)��&a�?R@��&��;]��i��+h�4��Y�h��e��q��r�{�O���`S���^	13**�7̐���ZR�B4r&���j�J1��  ���Jk9]g�Sv����+DUKˇ�֖���wu ���&L�+2�2k��+�|	�0V��Eʊb�A���<OF�#�mGM�e7�HW��EWL9Q0_�Ga���Ȫx�A5��R�7�h�,]���C���=�e׊UO"�bg�Z�k��ji����0�K�Gܺ�.o
��.8��U#�����n0��/���'�3�5����P�Yj�"5UȬ�zx�+��?:���xD�2�4��nJ��(^Q��V�S_�[���Դ"��*��xd�+��%��P��By�s� ����Ƣ�Wka�b"�
x=c�p-"4F6�L�\,��ǟ����WX���"�؀SBf�[8{)��I	���[���"�� �R�B��ͮ�X�yΕ����)#i$��Ʀ �;��E1U�b�r	�2�W��k	�^oiUeS���-!�di8�-�����:3�`̈���4u��I1�% s�V��j|��`lS��\u��<���&�E��n��'��x�A��R?�<�,�7ٶY�!DY|�ّ�h�&�9��H����Ղf��y꼮 s�����4o s%g|��C"�L��� �"����)��A{�x�Q���N���1��+�iH����i;A��ES1��9uH	DCM
�9�)�a
��-C�X|��g]�s��2煒4^���M3��P��L>1�*cb�+�j�I[��1�a�K��\)��ˠ���%�p���rP�
��ju1�)=(�(G����XX�#�=�tz��<�k!��z�u�=)����iX�ĳ�0Wq㱨g7��6�W�w���q5�^��n6І��r���<�-1-���;�	�j^誂5��7��hER]���tNf �'�^��?�!1ٴ�F��2_0����MM���4�6��������:�D̪;&����T�m�oq;Xo����U.o7b�8����1`���"%?�5a��[��P8`[;���p:^e�0|���%wBQ*�L���e"���P��ƪm;�Fq�ͣ�w�cB��2@Lr�Li�<$�j�N�����<\�l����$vN�΄TU�0�����!^xkl�
��]�Bn�3�J��prBE�;(� m|�칉���7^�i�ǰ��̣9��J�-b��7�k�"=�zi��(镱8��TǙ�(��ȺN�l�0���G~H%F�:��he���.��)L�ɣ�A̰��Hw���T��Q����;9�bSY�~��0̃[�j��[�n�$�3n�����*_ ]Q,�1&`�"G!��юZ��τ�6�&����.��'�ta�j�A�Ƭ���UO��zb^T{Į�i|��,��k�����ņ�	x���fWS���k
��^ĭ��2��j��!��O�sT�����>�	cm;�#��	�e��.G�BɽNc�+w��8��[�E�FC�p,fΐ�t�IY�v����_��R��/�f�uA)5�D��iV3�O^���b	>PLe��1n��_�
O����hi둞n!��w�������+Ί�)XT��3�]ha�=�3��+e�>��+$�re�բ���߉o�0�J���r%�[F��4?)��:�#a��i{�.��6�~����{ML)Zt3�;��МH�c֚�3�W���D�<A=�SŻ�L8lڱR��D�v��N��O �r�`\l��e��d���U3�(S�Q�ڨ4��� �kb˪K��k�Ern��#i�Glg�QW���Ϊ��_�S`�j��>�����V#�6,t��xt;�	2�!�9�exL��1ƨ�����:ψ�����ÞͲ�f�("���l�igM<a�9`�z�Z���VR����m�9=�C'���q�qc\W�hTi7�={=G�z��O�m�|L��
���)������t7�p��5I��뒍���P��D4���f��"�,r���Bj
�ٷ7��F��u!�̔M?�]4ws�v)�ku�\����y��)d�?8�y"��Id_O�t�����]>b�<��@�<bxn��"8=Z�g�F�C�]!e����������������θ�-���$h�ZR�PK
    +Q�HZc;��   #  org/bridj/lib/linux_x86/libbridj.so       ��      �}@T��?|GE#�"E�B����Pddd�(jd�h� �5��/]*t��Fj+oZR�/IEeee��ie�f��Ef9�&�k������93Ƚ��ϯ�s׬���{��^{�sxtd�(��������Z�%��wE^��tW"�����F-�%�f�+���SO�H<��R�CQ��� S(�G�iA{��7�'Ԡ=&E<j^�o���yE}{*���wP���Z����篖<��>�BQ��MP����S�x����z���Z��S��;�N�)��� �/�g�lk*=���� �K�.�	VB�~�%�$���y�~��3S'`��w��=Y��$����{���DO*�^/ӳ��-�E�IE��~O��j����q�'I7�����nJAp�LO��|������|�W�W�=���<D�Xz"�����y�~/&x�Ot<����t�-�n�߯J��u�(m;�5O������SG�i�2�(�q������	^F��~�$8�������{�����Z����GI~�A�2?��bJ�=W�}��&<��{=��s��'����=�']�O�Dt���`=7���e�az~���O�����$�3����^�m�0WΣ�M�&���\z��SC��7�c�g+=�P���Kd=/�s����F�9����:��B��������Y:���I�'z���=?��B��,h�YN��"|�29�?*�gL$<��)�{%=���7=�SNO=Oa\$W��3\�C0v!�����[!��/�ߙ��FO_')�u��~��z��s��c
��-a�����R�*����ѓ@O���}����]�%��y��Jؕ.��~��s/���[��~����*=��'Q����?�D�;���u�I�ÛD�Je���ߣ	�E�%�A�<�z2}ʆ�S��o��=�)�����ͤ�O]�bz�t��Aύ�����'�$x����~��ӆI�n�g�O�R��(�q���Ǟ�)��v��F��=!>4G�&�ަ���|�W��	���~�?���S�U��"8��"z>C]2�#�@��G������&ӻ���ջ��>EM��;Ǉ��������g����+c�S�����v���/>�]t�GJ��.�Q��]����/��p;���`4�|zd^��@���c����������yӇ��(�HOOz��<�#�[$D����M�c2�]����=�������b^N�d�ݗ�x�?���������I薐BI�I]�T~V�*<�^��[	� �KϷ�S�܋qG�]�c�<LO��/��۬����\z�mI;|m���B�!���$^K�0�Ϻ�.�o�,כ�N�v#=�鉗�*ʻ�@���.�KeY�yĲ��������=Ô��]"�����,�T"���		3
��PLs~D��{��������w7��v=�b�h%�b(TKS���()	ʹ�J��@%�4�AI�Z��.��]�\�]�]��+.3� ����C.��l)	�aJ�Ҟ㈝��i2��휄+�W��P*:IY�5G	�T���0(`���3����R���|�4`G�b�=$$�N	�Vz爊�!f���p&��ve	j���7�\%�[o2��K���G���cX�D���\����+�$%cB�����v��x����g"h�#\cu�@eX@�j%:$"�dk�C�@X0��O+��1��Hg�aUH1��簂�H�C�`T��"I�!���Fz�0L2%U�*�	�(�Y���H(�f##$�z�""1(Í��K�$1;!A�~�ON��ri��X��5b&����t�0�Ʃ6��u�jw�WᣱI���81�'�+�cu���:N�#�D��9>��W�I��t���`�����3Y$�8
>�<����A��1�
կ v�@�9[�Ǝ��@���N�KOI�1�Xs(b-��Kt|a�� b)��d:�I������0Wa~�S�Z�z?t��5!�e�҈1O�����"�u��E]W`��u���#���C���H�8��	]=K�>� � 97u�����i0��q��\���������0�"�źk	�X�a�xk_���%=���z��7��&#f@쪮��b-��k1�h����J���n��3��'q�-XG"�ź�
�< �I��9�u�1�a�=�!`]�����bw�' �V��шQ���:q+��X�c͊��`���za���B�>��X������E�j�w��͊�NL|bi�w�^�l^��Z��Lߤ�kY��|���z�п��^m�k�I�_���Ӟ�#K��xu�9tr�6}txkF����R��3_>���:���w�n.����;{�y�ļ_�+i�y�.����W��z_��ƕWl���z�%�Ώ/}2���5�y�N����_�L��s_�y���6����G������p��?�:����J�/�����y�yq��~Y�o����\um�{���w�uO<�t��z�{��.+��pQπ/������w�}�{��vE���>9q�{�c��d�𝕗�u�9!���}x����c�������9[��z��C���6����+�}6k_���B�&����g7-k�~Ujh�Ⴛ�G?�r�+�.��#p�O������l�Έ�}ʢ'BGX��|�C^:��\����.z�tݑ�o;o��;��r�k��f�U�9x������3�ƽ�(�H��k�i��{�{����b����t߬ǿy�{B��^US��9}�C�s?]�f��昝+"�]������-oO����[w.8���{�����I����U^��Ł=�߻�߿�f�������'8b��s�OJ��rqӐ`���#�w)2���E��q������-y����p�C=�7ՎVp�������g�m��������ox��M��<�٬�����{�}c�勲��=߶|c��Z\W�n��]�֜8�ǯ_��Č�֢���+H6���Wܘ�ᘄM��`����֗�*{����8�o�}��׆-a�ϼ�ӝr���MG����9�\�s�����<��_�<��Ш�O~{��a҄�5ek*w.�6��u����_��yW���x����m����Y͋7�x���#�,�><�bLi��K'_��~���9���滏,�c�7�z}��;?�4mI�֯��T��ؽ��_�#dD��[6�;t����z�ֻ*GN�����s�}ё;�Ϲ�݅W̪��~�nsF�
��OU����{�?z0�z��A�|��������1�~s�R�w3�[�E+>�Y�������K�������7�^Z��2��zӌ����c{?<���d�w_5���m=�)��븝=�}c���}h��E��Q�؛{�п�<7櫔��ܐ�ڔ��>v�ɺп�X[�x�զ[w>8)���/z�;.�%`m�?��X�8��X��_�y��[�/�9&�&�x�3��;NԞZ����?4��r˛Λ�X>��󗼱�?cg�x���8w��ǜთ�n���Ӧ�V<�B���9�I|���껟ȋJ,��;��K?Z׭߸�?'<�ӟ��2���5{m�7u;���W��j?4�m߮�诗��ۗn�g�s���tO�s��?�y��7��������v�QM3�}g畗6s��>���W��|fy�#�}�f�m���[\����'_�2�N�i�����ݷ�o-�����G�J�ҟ����_uAt��ߏ�����.������{�c�qH��3��h~"���_��m��k^�u�U�}r׳%�~���s!�ս�U�%#��vs^���ݖ<~�����L�q���Ӯ�����3o�<�}�=��$�*cw��Լ��?��t�ܧ�&<���9OV��T]����8l΍t���c_���(���9�N�<����qyc_�q����7�O��S2�䞈�����5g䇫�x��6K�)�j��Or�Iñ�룣��'Ӈ>��7~i�7����>���)�ç�$<x�7��o��_��\�M�ħ�=�q}xA�&��D�#��f���>�������ާ�!X��?�\o|�?�}�3٧?����Z��y��o�O{u]��\�J�KR����%H|���q. |L֍�ÀN򩶋�v��S�~Z���ki���S���V��<'e����;1]��8�~�9��HG_F?n��0L�ד��эZ��ԟ�a�OG���ۥ+?��?0�������'����X'!��/e�X��������E�>�ꇴ��@�W���heRG?�ʟ��7��k)?��JeD�"�b��R�AWg	/���Ϡ���8o~�[��^��
~����s�|,֐�(?e��މp����)�����F]���|v���7�GF�2��g@�o"~[�k�{�u��o��Q-��u��(���N�_���N����W�]��}3�Ӊ~��������ke�>2�h�RB����J�v�f���	�d���K���_)���bOx0�?AW���x��R��a�Ξ�&<^�����:����qiR�w�"�׋=�k���:}|C���J?����8O~�"�'~I|!�=Eo��^5����ȿ5�gG���߆e�7�|�N4����R]}={�Ϣ��U������I~�h��~���^Ǩ��ӝ���N��j��ז��0P����7�>JI�]d�H��ɚ����x���g����;֟죿&�9��a�h�=�\د�W���:4��筪�P���D��kd�kTu_��C����_���fb���Z�!T�q�&/�b��?������/��S�x�Z���z���n��:�w�������S���C����aTޭ��I�K|v���d���ЏP�K�����{����n0([%}�W�>;�P�q����&\������%�������j��M�-!V��9�߆M��^���b?��#qu�ǞNi���E�$�ﺍ�>�*?���&�gx��.�8������-��֒ \C4�i%~k��+�b��@}�Qp�A�L��*�E�]���@��@�yD��Z�V"�ҁ?D�^����7b�6?�^@�{�g���b�
8y#6j��k«u�Q�_�����ݢ��qj��wM��a��v%��تx�7����0�WH������X*�տ��5���f��Ĕӊ�>L��:�Z�W�nq�������n �_�|��c/H��!���~jo�X-^��D�*q�<��K���(�S�5��F��}�����8O �6ɿ��[^�ګ�gI���}O�[q��O��4_���#�Bk_�豏�@�3r�F�1��-'�����R�)��=\�g!�X!�P��T~����ɾ�i������jt��Ix��L����U�`�_��_�$�eݮ�+�
F�h�/�y��K�g����~��<���k��R�����2Q�P�!]|kCLl�!�/#�t]h��?�>+�^5�l�������W����;�PO�F�T7��"�������4ydҏt��)��]�h��=�×�>=����2qV |�ϔ���>���H�~F}�<�s����^cu�K�_}��]B�i��/��ߖ����H�E��i�7�c-�����:��J��5j��#}6���ǩ$���x�|�E�ģOQ�8�|k'�$����)d���C4^�t��d�u:�K�Oc���=���O����&L�G�9��]v��B>g�<~��v�����)Ҥko(��sFj�w���������?��2�u�??a߹D����\go��~�N>?"�;�x�=��o���U���� �7u�k���~���Z�8��e��%y�t�;�����}A�k���Sz*S})���
��EW~O/�q��3���=J����?/���O��#(>1��d�����R�BB5�;L�R��l�_�|?���K�M��T_���2�[n��?�O�����
�����x��̧�(����׋3B�+�~]���F��zL[PF�CQ~���!���(��͟�I�lN5�E�i|�g�k���)�7w$��D�����w8�o����Կ�h���_I�����c�G�m~�O��0L�ǩ�����}$����h����g�<ji~~>Dο^�[�r+�_J���:_}C�̤�µA��c���S6�{��7}�����c�Q�o5͏պ��'���:y,!{�^+�*Y_�Z ş��;&R�x�x�3qO����4�FI�;�7��� ��p����l������g�@Ϳu����}Η��n�����?�O�<a���$�CI�Ku���`���O�V��.����V]�_�����/i ?��OV�o��=���|��<�[W<�_�_�A[����5F�#��,]��߬�+{!����g��(]���0n ����wH	�h�����n��߲�����s2�?��ԿS���a�.��煔�YG�
ɳe;�S��sz���ڃ����Y�G�� ]�wQ}t�d���?���k<O��J�����:t�N�AO�h=��(��_+�?J�ݮ�?�ƣ�.�@�D�W�%��[�h�&w���| �{����.�' /#�U��� �N��{�����?�t� �g��eܥ[ϛ����w<��������0�۠�%ŏ�i��/�?F�o�?�:��	���
��]�J�6S�_)�m��M�_��������8�G��
ك[����#����C�>&�]��������BҿD��e���L�hѯH���])��&����#�Ѻ���ר����I�e@~ �Oi�������k��]y�W{���5,�߫�O�N'�:B��47�P<��	�E��c�/;W/_�?��W<���ĝ|��~���@�7ZgO�|����H�~<Y�O�i�Q�o���yX[��`cꤸ���K�Si��\��]����?�:��C��N�{���si�=L�)QG�v����D�g��#�8��3q/����_�
|P�n��_���e����2
miiJڴ��%mL�miY�BsvN��\�z�k~�95c��,���e��@֜�;=�NI7QTd.RF��͘�1"�j���e5��/��deޖ�e&0�0;%?'�J(�D3�8/Ӗ���H�9�\���I�ʜ�#�Y
�g���i.�̶)If�ȼ�
�ϦO�N)̷�3m�,%�0�`|N6�_���m��(�T�x[F���iV2�挼�}w��l��f�$s"������ʈ����6ې|�����Q���2l9��j��S����S�(,�R�hKMR61?'��,s
m����6K~֨���TKN�,����|�5��H��Y
�������l|arF�M5-�\X���f���`�������:Lԥd{��}� N�/�N�Z��u�'#���E��9®��fd�h)4sn�2!/g���<6e��(.,4��R͹l+�m�ř6�K6�
F(�">t��
�Q�ե�1�
mL��dg�q0��6̖/T�"����"���S�z�1N�ѠdS���8&Ϧϟ	 FY�38I�������*��dd0�#,�H>˦R���r��	{�5#{b���kO�'?Fp5����:�`�cn�٫���!���	ySE���b�_Ne�����ܤ�D� ��Y��%J	�o!#�l9Ŭ��}���^�%{F�6-#�*9��/)G6@n^�f�j:*�F���]���c�T6��:��~FV���L��z�y�2�L$�pXA�9�,�8�����N_r�Y��1'��x�.��:���ʱY(S��<sy�D���U5Iɟ�%�:�0�"ARˆUr��6��LU�}��beý}�:�4�<ԆJKSS��|��45���C��x�d�j�����ȓ��@�>D�$�0\3iU��%t�Z!!v��o��$5�U�C���)B�>d�D����C�tܘ����3�d��۔�b�}XVV���H-{gq^^��j��Ӭ2V��
�F���m��7-_�?��KD���� E3ZE^}I�*hpȰ�܉�D��.қ@0���8��2&�b�<��4"aΞ�8ͧ�d�#|ТQ9fk�.C(���J����3���Ь%ge�I,��;5�:.#W��ǽ��Ts�o�\�:�̙����}�df���Sg�u9�fb'ϓ�eL�/��Q�e�R'O�t(���2�l��a��Ӧ��x�C����u���E�0b8J�Ĭ�Bs�MO4"�Z\�G�H��-'S'`,��T9J��Og6g!�M9.҅f��+䛟7�B%�*��R�6X��%��co/�i�'XS��4WA!�9#�'!�<��s��d�,<o���Ƴ�(YV��
�G��ܐ�Ss����)�(�EUQ4Fd����<�7[E��?������̷E��l�>�G�'��<-5_�t�y�I���b*���EӒ��!	Uq�9�NTsV2,�Ɠ��j4FS)"����'��/�6�J/�	��9�Y�H�^j4�[ �lZ�٬���a�)L�/��*;�����U��e����fwp�"�Ԙ<]�<�혀�,��B�~�˳�4��deʉÿ�
�iS��@Mq'�T��������ss���'��Ǎ��>В�C�d@�8�h��?�*�˅���핣�e¡�m�B:A6�4�[݃L�i�(jwm��Ҧx�H_L��8���n��( �� � uF>o��1��p��<A�����N�T���W5{mS�[�UG��0�3�[�欳��R�Bd�E93)��<Jh����]�f�efd����mŜ�Y�׳QNn��vY�rr�Ns��x����m&c-'-�1�%i���Д���S�_��K�
P��
�y��?-&��0ï4��N�S��-��ȩvZ��H�9�/��,W��!e~���)��n�5��M�Mg��SJ�/�1�ug��)Z���NI�)��K'r;��ٔq6�65uJ�M�
@�Y�t�����ݻ�xl/�S�l�;V?D��nu��y˴dv� @�.�g��tg��Yh|�锁��8 ���S��F��Y���~���Y��d�4A�ic�$9�9{v���l�#���|+g��و���)��o
���wV'�#f��x{�S���v�S��ECgS�Y����)��W%��e�Ϊ�Ԟ�����̷O�)�`ZL{oCg�������NX`+�ʙ6�3��b>I鶌�b�ᶌ���A�b�m�<��m�B|n�+y]��GW3-��gym�Z�n5�R
l����y�\�{����sfδ�LOZ�.�׷��W�91Ö�Xs�����E�C$x?�K��D�QV&�-�:^�Iy9\��Ԧ�M%�����͙�M�H�78-�ڲ]B��T�l�\.	�}���f��]w-�L��h�jCz2�;�`��5 )-���Z�\?e��;*$���͒S$�a0�����^�i�m�+�UDZ��E[Ҭ9y�3�5����Ԣ�vJ#G�M�~2DM�$��5��@�5�Ȭ��f(��y Y֌��ByP/�y�f��9A�0A���o���=��1pq�e��Ql�i	��e�f��թ���wð�r�$)>$�Z���g�� ��3ɤSi,N(2�<C{0��(�H3g!#��Y$NM(��dR��#Ү%'�����+f�u����'������g���ݭ�2E�y�<Tj	��~]8������������K��s.�J���n\��L~Cw%9���L+�$�Fa��m����E}���n|d0Uº�6J�W��HxT��P� �Q�@	�$L�0Q�d	S$L�p��S$L�0KB��V	�%\*a�����p��k%���^��n�p��;$�%a��{%tKx@�	�JxRB����0H�	C%�0\�	MFJ%a��q�K� a���%L�0E�T	'I�.a��V	$�I8S�	K%,��B¹�IX/�	$�.�	wI�(�^	�P�Q�G�(	�%��0N�x	$L�p����JX&a��s%tI8_�.��Z¥���F�Z	WK�Fµ*�n7���%�u��34> �J:���d�2(@�h��o�� �EzL3(3�%�>`PJ�Q?��O@�A�x�AqF���㨟��"���-�q�O�m�O�)����	�jPV�N��ʠ�fP� �J=��e3�}d��@�A���#�`���7(����} �O�x��Ӡ� �I����#`�A9��#A�Ҹl%�x�A	�E���A	���'�
�x���<�?�l�	��!��d��7�&�~Av���!;oPFV�d�Y��9��(�?��2��p%�W�򏀏��+J�F�?�d�?ࣤ��d瀕��fP* /!;<�wa�d瀥e`&��z�?�+e)���� |���V�R��0���LvXH���� ���$�N$�>B�����G���"�N2({2(n�!���x��`�A9
���x�[���^h�2,"�op����Z$�,a�FCA7ʠ�I.a��&	#%��0Z�X	�$��&�*a����IX!�\	]Ηp����+�p���.�p��5�J�Z�5���'�)	��%�0H�	C%�0�N�2I�)�K�%�EB���$�)aP�A�G�fR{�3H?��H?����(1:H?���~ CI?�ϐ~ _ � ��
�,�W��h�>Ivx�W��4���xL���_��G�b���4^��x�F��;�W���d�41�24^ { �Ho.`O���׀�H��ͤ��p6�W@+�;�w��I���i��C����+�i��
x+�W�34^��xE�9�ee�e�4�F�xt��|��+�4^��x\H�؇�5 ���� �F�`�7��do�����g��� �N��	h��	���)�h�׀O����9�a�׀�I���H����D�D� �I��4� ֒}� x>��!�?�U��P�?����H����!�^@�4�|��������%�N!��D�0��5�����/$�����G��M�,&�s=e`�?`��j�?�C�����B��0�?�-��!�Z�_��|��p��"�?���o I��1�@�����ݤ��I���4��1(!����ד��R<K����?�X�����n4�������?��?`�AI �N�\C�g>H���p�p0��0�p%�7��?�T�?�������m��M��.��~�?�$� ���p ��R�?�ˤ�=4����X@��C����?�����&��q5�'4��xp�Ao?��K�a��������Z^g��Ɨ�������l�_��xS�uI���x��F*ں�S���-Hl�co�Z�M���Y"�W3���H�.��^�o*eY�N�T�8ޜ�$ Og����S�>��EoJ`E-xݸ)�q|}ݒ<�qTeA��BO�O�7)��j��IS���2�����8��Tp�ǗR,.�?�hڲ���8�\e���3V,+�����oK-��q�fY��g_���q��������,����e��q|�����g]������o��3��YNr�O���7����X�����^���?�Z����W3^���b|)�x)�+X���a�Og���<��լ�	��a��f|-�x�u��!�׳��+�of�o9|���x����v�?�����?�X���Y����������Y���("��3�����3~����g�$����)�?��q�����3���[Z���C�������GY�/���8Tm	��8�Lo	^�8To�g �j���-���)X"���_�D/e�a�^�8�<bI ��8L�2x
����%x�0�$�ьc���`�d� a_���3UM
�0-�L�-��^��g�f���3�/�[\��az�����#K5��q��e��q|q�R��g�iY��g��R��g�j���g�����g�k���g_Ƿ4r�/e�s�/c�s��`�s��������3�b�o`|>�x�X��k_��^�x5����ौ�`�/`���<��Z�?��W���'0���<����ױ���0^���0�����$��?����?�����?�;X���w�����7������e�s�w�����`�s�oa�s�?����3~����g����8�����g�����8���$�����~@S#��@���^�8��%x-���#�W3W`��b�<x)�p�8��GO ��8\�e4��c�� O`�Âς4E3<x�p%��� W�k���r��?�R�?�p5�
�?��]���z,���O^��g�Ȳ���x�Z�?�pM�5�ƭ�����UY6s��o��3�e���g�x#���R�?���2�?���
�?����W��q�x��Y���_��^��"�?�jƫY��]�/e�/e|�x�5���ײ���0���<��5��ь�e�� <�n�k��?g�i����m�{���a��b?Zi�@�+����+�'���f��|���r�c�G�������v���s��j�:]�u'��5]bؼ�d�Z���
�F%���lk�o���	RQ�]\�]������&�}�h��ӎ��a4�/�!�#�O�U�h �U���S_w�����Y5���m����V��JN�nqM�Q���w��b�%��S�{�T��&�M�;Zpvw�L�N�)�a5�9���`�(��Q��u�e�@�dD_���f�<-!�"����P���J���Gb����V(N������@j��7}�3єL0ȝI���8t�pL����7H�N�Y�`����tмV�;�Ln�cӿI�ӕJ{��8���UG��I���!��I�n�{!��h�:M�T��N0�``e�)�����s&��PF��PGJ��*��[:D�� ��@S�S���E i?5�L5E��9���#B�j�M�('����$��H��&Ss�d(N;7����H��djM���>��S�Hg L %������[U��������w��������B��ۯ!��.�5���|z��eD̄8g�GZ*K%�9�%���ᨡ�0�<�D�z��	��
���n�@��ؾ��]�d�WV��j���uؿ�P?�nK�x��KU96AZ7$}@5PK�A}IZ�BJ�kR�ft�z7E�w#^hʇ}i�����ŻG
{�����Ӓ�����N�����/�����hO����i����������Cm�	*���#̀�*½�/}�)-D��5B^q��@��4�SG�v�o�-'Hų�??��DsԴ�>j���x����ln<��z!r]{A��Pk��?��I���4}�Gv���h���������r4I�b�&��S���Gtڶ��R��4�~uT��ѓI��M��;��V~�4_I��'ҝt�I��&��C�FFA8��Þ^	�;��l!�8���95�;uU�2��m{}�do}A��O����O
M�7P��F�E��UVm�"!��pR�{�h:�y{���AQ��萃�Z�?�|W�k29���R�^ȈR�^�ݱ�|,�Df��|��r��Yo>M`�G+�a孶s���8cpv*�!���t�����b"��'{�ϑQ��D�$]��G?8��e�X���qpLNd�'"=�[n$��.ß	�*�3�H�H�|���(g��yF�'�ؼ"�(��f e�{��f�ɑ���A��)R�ߨ�~Ȁ��C�SKF�|����x���<��F��9��J��;���ۓ����cP�㷜}|�������g�����?����ￛ���G�����J�7�=�z"K��_@��TS�������ޮ���/fb�E{���>���~|��.l�C��߬�玀��n>��謾�Z�軱����M���~M�g����w�����П�C�o�h0�ouʳ	ZoD�O��SMq�d�N&j�<���`���U��z�b�{[��8O�
�+����il���|���l��}g5��X�*��u���oF����k�M�W q8Ȗa�4
[,4-8�9Z('�^�ި{�} 1�Yf�c�)��;�+�Fe�M�J!�z�ג�R� ��f��*�6"�ԧ�|�����1u�^��9E%��є�c�|�d("��%����/ǻ�����C��0�.�8z é���>l�R����p�j�t�8�1aĦ�E�c.�3Y{�N~PN�b|`��X���n+�n��I�&�ȻфI
iua�����zJ"4%�٭���*�����Ŀ+���NK,��ô9���-�"܉�P�U��'��8z��Ѡ�Uk�\f$��D
V��d��	��RVU*-60��p�<Q��j��eC�.�Su� ��'2���qu��sj�@AÀ�D�����>�qSG������]Rw_���lO8?��kM8:q�pԘpf�1�h��*X�Ӟz��5�U�۰��L8��.|V�;�$QY��!6�D&D��?��@��W�Yꝃ?X��� r�S3{#��t�0%��3H�4|��\��S��)z���]I��׉$�Pw�? �nq��"Tg,��Fܩ��1�O�}̹�O.�3�s����b��|���)��C����h��g�珛��ba$�}��~�x�f	�V�c��6ƃ������i�)چ�H0��7��;�`o�.B�C�v�ĳx=��!�#�$*cu���`kV�Y�Y��*��&\��[�I�E��_��E�G��{���d*ku��H��B7�qei��_��<�b��܂&=������e�A���U�5'q�O��f��FSM�����8^yD�<������*f�I�l�L�o�M4/���'�C�H���������ˮl�0!�����
��FQ?��Osq?Ĝ<����wI�TR�J=[�E��_2��K6�)A��!��dSl�g�>���k�]1��ǋy<�=w?�>7��^ /�U�D���+9�&v��k��Į/��mp��O�g/v94�l�_�{�ŕ��ϋ��1R�b�&ߗv/� �
g���(;Z	��&'�L�V�	$g�&9?v#�p��F�� �q��e�c�̔�ha\n�8��v �����n�
�_G\1O��D�(��1;KDb
��4�*���p�n�o������{<����Y�1����9I�S���������d�Z�����^Q��z�W�r��>
~5�-ا�>�Ȥ�Q�U������t��V�>Z�.H�=|Ƈ梁6"�?#���H���8{��1<P�j�ϼ!�Y�=�H�bZ�w���(nE�!b�������X.�9Cݪ���鬟yP���h;�����U�����ݼt� �M�β��� ]1u���$�h��q�3��꺻j&�Ѝ�����[]�
�c#����F�/����
t`��9"���4��T���i��q\�qe�Z�]���ݽ�'Z!��mO��Kd�7� 8��X��_/UX�����vi&s�WQ�Zۣ�}�.ǉ�H�x��j%k�z�i�o>�wy�;�06]����-{EÜ��S7��5?����a���O�|
�ڂT�e��ط'�֞��U)�|TH>_<�ݎ�g��Gd����@ӼӾ�����xUv{q�iMر?j¶��Mwj�',�TiϔC��>�y��gr�x����%�6V`46C��{y�7��a4v"���xb�&"�Hfc��meu6O�b�[���]CDd8Ϭw4Ѐq�-��^����'�'�3�Ϳ�����
�do�� 1T�qz�� ���Īq��9�&��r��51��{bB��Q�/��*��_P��v��03z�c���`��h)9S��F��Z�9mT�0Չ!�%.�d���S�S������B�����u�ڈc�1�{���N��\.�����q��H�D����6��C�C"�G����4�ד����h�p�zѦ�TpY0��;e{[�h�=���ӫ��Ϩ������^��4�� Z^vF7O��'z�[A�� �qƳ�����v�(�6��z�H��T[2/����������1�Է�������;Â�j@��F�����������?�o�X�-��[h��}��11�7��X/��VGz�Ǐx�ߍ�V�J�iU����M�<�W϶����K�o�t<�GO��=|���9�HR�W�"�vx��$��ݓU����g5�9�Տ�\����g�nO��t�Þ �H��BS?�he*X�u/��-�0�*��B��B�2�xS>�.�3s��v��X�w�b�z7�ɘϚ���wM������.�Շr���(s}(�h���o��v){��rr���� D���~T�:��|�k7|��+8�4Y�j{�f�T�f�Oݓ�kS�q۝�	���Ǆ�d��YU/wn��u��9N�N2�_���;�弃��^��E�����b���n~s��"�g�%}����U��侎���ã{](�VBa��|6�.��S������](v�rޚN/��|���>X�z{c�}���%�Ȉ�\�V���N��W��>�{�U�VM�~�c��)p�B����ɦTZ��羭^-��&�M��x��,�,�����;5��ʹ��[��5u��+C�X�D?����Ss��+��'7��c�?�"��o2H,��
��r���\Mp#�E#��pY���KXgo?qi�������]��k?�єባ����Q��s{N{W�sNĮtykp�e]y�8HUA�6yH1q���[��+̀�I{,��:ZS�ݲS�)l�KFQc���D�k�HX��l��t�O�|�viX�����)G��*ݔ����A��ss�J�e?�_v����%�,߆��<�J�_A[���Uow��蝚�m��=a��D���l���]���K|:��-򚏹?v��T��-�ߔԪ����mDD�bG�X܆��(����E}�vU���������ܮ���I��#i�L0����K瑁rW�=�+�%U�d���7x/���ʒ�9���\�S�[|�$��/r�M��:��.�5���yX~��wCm�k�z�N�J޲�	��K����T-h��nT�mTdAS�Sz=�<7���G�G��c緿޴�S�Is+���Z����S�U�{�S�\�Jތ:rCM�:~��w�H�' ��������7���NxAe��)��c{�s��+mci��5Ҩ�+ )��;q�әgصr,� �����]�UOׯ�?��t�W���5��������+������N�?�����#׵��j�e6�P�z�NL�x&Q������C�n�n�[�ų�gZ����bYՔ}�g}������B,9QQk�aDc�w�,�mrGw��c����������H���-��z���&�DF�"-�Nd\����"�?.CUM�u2t�F�o���t��9�@�	�{O�B��s��>��<C�Z��<v;�����1��"��{�ٯ�#�p؆�{�gs�{������6q�S1�yw�jJp���x�"��	w>l� $�v��	����з�P���M6Sx�odj�F�+r�����(0h�c�]l�DQMdJ��n-�"q��������%|;��ʇH!�0z��7�z8�­�Ñ�s
����7�w�����|��8��t.j��r��u�](�-�u繂�hw5�T���:G$v��1��
��V>�����D^���>ۆ=1�ǻ�r�c��[}��/֭pMJx;���#�]��߫[Q�z�W���5�_�x�P����N�דk���_���w�ߺ�T׿}�������s���k��������������;��Q������x��_����y�w�?k���c��(W�h�v�[������*��*o�V��ou�h���?�����%^�!��I�<-�ɩ�WB[��+����\��a^�$��g�~������yO�O�~�w�OO���7?;��SӖ��8'2_�ް��AٙhJt�,1
~/�4�ݠid�QΪ�T�N�)��S�A꽐)⎈Q�O��&����+���%��kW��]��\J��n���v��혿Ϸ�������?w����)�]�5�RM��y%ZYU��/jE�)2��j�Hwl�ˡA�U�D
��9��1WV}(��_���H.�4L嵅 /?��\�2&^��cS�$�����&5;�EU����r��F��5^~��P�^�}�n�>�d{q�U��4^F��aSp��V��^�'�*������|�	�U:w-����0��֪�������M�V������IE���P��at��;���5FŠl��1q�r�����Pq�F�Xhu\Yb
w�}J�|'e�cFZ����wb���}J���M�	/��m���zY�=���cԏ��+w3�jP�)9��~ �;�ȭ�W�Q�_ �����a�f�����# �G�K�l�䪺S=��^]����lt�T+�T����T���*g-��ɆJ�e`�����5?]�K;DL���/~�)�� P�0
�Zb�<�Ņ� n9٤nQ( ���N�g��q�ٝlW�گ��F��o���v���L�"S��J��/x���h��aU�| ��t��Z=r��Z����3R:9l��R���B�[�ֹj[�1p9Rᾒ?������FX��Pi7�(���ᑞK��D�՞����~ˈU*�"_�j9�E�-�n->K�q�c;h9��<Ż�t�-'˖s���$O��:hy;�����E�[�![^v���<-�A�S�寽[���%R�?��壞��t�r,�l\��r�b�-�dˡ�;n9���U����.Ր����o_ܡ�^5��2d/�#����C �~�A�����;�"���N,�IƎ��D��%/��@��#'!�)���Si_��=[������U�\̾���� )P��5K��"�hL��2�=g�p���0�ߥ18oSd������t� 8�IK��!���9���}U(j��T�[���U�tZ+�w�A}9ѐ�e�x���ʿp«҅��%��'U�b��F��m��.���*��y�r���d��Y��Ӫ�2��P��={��؉�~����yߌ�����F�.�����b��v[�O|���Ep)a$�&��mB��X��ju��w|�rՎj	�*�6���毫}<��]e?����i~&�E���f�e�8)���c�T���@����=�G��~/H�G	�C^�R�-�xF-���w��ZO;�2�/i��^e�B���]�����al#��~]���
���Ņ�B���E<�O+<�]#�AEUV=��Ɓ`�"�v~�vw,�2�L^�1����]�|���O�����9]�JO-���"s=E։�P��U?u���fx����VJ4�zZ9�q+O�_ޭ�n����"�1��t{��V�z�����/��J��HWO+Wt܊�#�y����>K��f9?d��%V�}�|��Ƿ_ĕ���"��[�і
oT`�tOzO�Z��.��7y���)GR��Zr6��w�G�S�<��u�7"��Ҿy��<��s�K�|�S89U�|��Yq���Kލ�|?�q���)�9�Z��F�z�j��%/@�O���H�<��8y�+Z��HN�䥺��� 'g��A��I�|�8y�R-��M�\�K>�%�����@�܈乜�K�ɣ8��N�o!�8����%/D2�t��'���K;�SL��E�c�bQ�7	s�L��.���yb��V���S��_���{8wJ��^%�x2'N�s+����kAY�y�c��:[_���MW�W�d�A^�\x���x}��֗=�O8�r/y�U���L^G��o�:3����݋�p������Pb"����������Af�������s>S���u��=�[�Y������C��Zy��(���|��#}���d\����q���jB���Aη�:{�����������m��\��T9�wyc���O����}L��u�W��7W����Ow����n����N��%���E��)|���,�V#/��w?ϙ�+,�J{����x'��������;��,.��xƍI����{�-~��</r-�Cӊ�p�*��-�
�n�.�y��;WޝY*q֘����f��{f�~Or/zC��̂ZD�����8D��|�����c�x@��T�L�`�J9��(]������Vi��{d.xq��g��O6S\�s�Jp1�eVT�$����_VR�)Q}���O�$?���i��*��?���T�����V��<|�<6O�X�;�C��8v�q��
\�;\�]�/�8��n�:<���M�!Y��5��C.���/i��-yx��G�{�SW�j�+���6VQ}fG��g͔���,��MA?)ЃA߅)��$Z�+r�%�W��'�o�RUh\�v�Fv��S�N����q�U��8Y��U�R�l�����pxŻtHZ����؀#�l���P/O�A�
yq�ζĉ�t�Z����Nݵ������K��q%{�8f��)��s���4_��#*�j�L�r[�cD�p䪴���}����7{�.�+Jo�D?��2c�6�?��ɧ�5n�NE�����ނ�������ϟ����_��qG��K1uT5��ٻ͙�)Lj�6*s��|7�ﵑ�{���CGЪ�?��z�$�Q�_o�~�3)����������.�C���i �8��oB,��#^u�7b</˨~���ea1���������/bô����f4"�61��j�촿�V��<�~��^�!^�qpë䯷�\~�������T��pq��8��ޕ�3ܽoU��4�O	��^3րe<r_����o��������__�r��z���ū���\1�x��0v�k��7��w���9���D�q�7����Ӥ���2�>W�)�/uxli�NK����
��J!��y�<1����1�q�d��GE��2�{.ko�a׎
#m�rf/�xS�3D�I�A,Gu��_ulu��w����8����s>=_}CW��-�~����lk�m�����Nz���Nj�D�[�/�6V�;��"N�����)\�{�
̡/����X�HR}��W�2&$_A� ?�s���t�8"���Hu=�j0��-n}a����������Y�S(p���N�������6���@���C�	�����gm!��ߍ���9��wly��[�f}A��A��K��#�+�v�A;;�s;�)����M�q����N���i+n{�{«�ul��C����U�:�~��g���&��!p�;�17&>��|v��g�x2��z�-�Z|4%���+�cz�?u�^��B@�K-��\�~�v$׻v��N����J��eؒЉZ�w��5�\�N�'{O���'��ڪw���[3]]h8��������5��:]���5���]k��u��\�ZSX�Z�	�T~_'A~_'�}�U�u�({�8���x�7vbm��\��"����C�N�m�V�y��d�r|bT�k R��-/�Eu��=�����/�GGwq5�A`�`_�K��gD�{�t�,��>�Q�I��&,:�M+!��#�6҉���:2əd`��-�}�v	/����S�X�W���	�R�BAnm�<��m�3��r$�%�����e��HR�����qW�d�8L�̓�4�5�������o�)��x�7���`�!@�0�c�3[hPU�a���2�q$A����_7�m1�&W����;����U#�IBƈЏ��(�=����%����=1�>��cV�wo�G�B%��{�O�F��Cƕ�n�v��|�!��g��,�MFL�Jp�~,���4�������)>
��'�4}̟�ؔ��kzE��Yi|M�����IA�wCHO��� �W8Z�Ea8$68�}���2���{����?|A�e��!��J�~q*�� �[A#����ټ����8n*6�����_�p�x�W�q��y���&��v�w;���tW�t�/M��M�?dq�����e����<����E>�H�'-��n+m�<�u�<��v�<��w�<��r�<��s��W���_y�'��
:yW�Nx���C
��E;���	v&�ʀ3��_��F��&(�O��X$�9	9������T��w�<��I4,�
"�
��WϏսz)��c��;k؛����|X��=���e�cu�e ��^�� ����f7�{a��h��6��J�V��v�N���R�c�f�U�G�d�zN|��U$���B;�'��9�����f[Ԏ%��|�Y�x����K��>�#Ϊt��I>�*D�'f�)�)dt���1��q�Ȫ,�a~<F��7�?O�x7,��n�W�D(�޷�U�f>2L��Ǝ���d�#c�y={n��؋|2%9�+8����h��㉻H9�F��/�t�N��p���)��	u��0�"���E��/V�{r�6>����+:M�j��	��3!L[߫/{���������HC]}�ą�\�C��3pGO>�Џ����36�@u�e��y�Ǉ��6�J<Ђ��0;�g��ا4�9[I�ދXK��m�O~����'�S�����nNZ ���i��8B�,>��>�,&�0�u����v�^�K���7��H�"_o̒L�L�L��$58���Q3��t�Y�Q݊L��n;�	�b	�e�Ď^2y!7/�x�S8��b�!;����z���6���N;;�@m�0���nSZ�.��N{��O~����D�}���.���g�-/�'9�[ڭ��|��v�ܚ�Qo:��o�bf9�V�����i��[�xkẊ�#7?�t%����Ә���J��l���/�φ���i��V{}I�6q��Y���/w����>�� ���{$1���H�i.�FQ���(�м�Z[)M)v;�'������R�7�>��۝��g��!Z-��)|�r�i�6D��!
7e���YC�ĝ���ml�lx��.�w	�$���Q������Pb0��+B,$�H�r M�I�*=�P�~癶�F))1���EX��O����{<��<�zk)U?���"��7?Q�/��Ì�ro��y�W����,��l�~���Ѿ��8W��w)�;����ug�ZG�o"�D�1�7�'~'��i���?��o�ߌ���Z�8V�ň�y\�p!:�9OsRV��r0��\UU�|������h�d���T ��^���"(�����Тr���&Ǭ�rf̨������>�Fgt�i�n��C3�1��y�k�}���~	Z��{��km�]{�����k���>����N�?xK��4#R"��G:fD�e��D�S���B6텣Q����Ͷ-(bwC��7��ΚmTњ�v�ȵ(�,7L��K�,R��55�"�*U�GM�R�nS%�9����
���P�P^���?���y��Mu]b.\!<!������9�T���K��������O�����GS��o���f?�ʹ��F]���A{�GdSyt?��xq�E�� ȋ=��Bk��&{��x�� �\}۪;�=X��$�)D�r��IF��@,��)��D:a"�[3�c5Ld3���{��?���V����� �w~d�7��mg���<��w�f��{C_lǚK��a������޻���}0R�ȳ�v��o�oۇ^���n���ttf݁x����o�Y���7Y�,'��&�r3�75��>�#ݽ�%���f�9����4'Ǜw�Gw^�=��d��d���,r08%�H�7�5yK��q?fu���k�������BF�{%Gh�3���ԙ^�[��Ynd��JV4��l4?��)z#��Y�G�Δ�RKՠ�B��#�/�2ȪE7��df�T����82]#������*e6Ѫ*����0{"�I�Ͳ=ز����GvrA���?:�h���(�G��u�V33I����P���.�l�M�-���b�XVV��^�HvA7��ك���0���ڕCv������J��!��x���	*��[q��M�D�ȫF&���#��q/�7��P��e�ɞ�E�N=�O���#N��OVʢTv�p�b�O�\�$��}�"�����S���<M\�lz���ȟ�A*�v��l]���n`O@�@R!=�z��	���eɮ�g_���z����)�����ߏ���X�����뽵�Qs�|��m��o������������X��p��_����ۿ���o�������^�����{��Co����Y��94����ڿ���un�����ul2��q��\�����UZ�=k�A�W������Ծ����C9HZ�ft��Fq�6��&2�M�TO�a�:S���_y��v�m0����|��j;�ǟ�F�oE��3I��yʡZ�}O��謹OxI�S\�a��8z����Zo���΋<��L�ع���^k�㻵��(\w����<md��;�]�O�՗#'��5y�#�d��P�@y;���'�ט�f2��W�����K�$�t�Dn�҄\Z��v�.��,�����t^���`�2_?2�:��|�F�%�GF�e����/y��䕣�k�a1���L�m`�?s�W��4y%h���G���:&*C��6��"��Mr*�MN��u���Џ9\�\H�w?�D��v�w+׫(^��ʥ���#��,��M�����'Z)D��������M��H����xZ[�e<�4��S���D_H�����E�1�^\�9�����t<e��x���~�wY@�r?L�	�����Pd{��O�2��u��_��2�_��V��sr���}���~'�������R�涘s1$�(7Uq��U����c���̊�c�_y��W{_d<J^�7^NU����ݕA��y$�����[�V��х�v?�x/� �d�����hd��Oe�w�Ԏ]��X"����4u<�����acT�?c΅��&Ti_����P˾������汝�{�9jzg�w^���W�F��[�k��}�(������/d�����{8d�dK��VzN��ϡ}��<�o�8/P��S�s��Wɫ���H��,���{ y!���m͏��V{*�_�y�=��ޤ�5���|>�7,bqA
��*�c0�#<���L&	t�M�5y%��x{z��+��lhϗ��V�\W�g�??��Qu�!�E�_�|�~�wJ�k+�dG2�Mʡ��d\FD�8i�:�-{���`%0�a��ആ	��0!�g��d�A�
/r~��$�Еnr&?����x��ԍG�&����E��t;:�A؏����r�}RO��䷆>}��v*(d����!9�ު8jxy���{;��~ڷ�"*9�`J]�"�^��RU��W��4����C&ٜ}�,�#=m���<C��[Vx�r�J!�&�٘��@rD�F�<چ�ǑZ��B,\�>$
}H4�a�,ײ�$�e҄�����G[s���j��~�5�� #�2-���/�mt�,��Ln�d�N��;�y��1kL�nX�^��a�Lǖ�*iZ�m��x�
=�r�XoĜ�Ȩ�o)l�庾��{�o|����*�daN7��YA#��o���4�6G1I��~��cA�9��j����q�%����r�����\x�=\�]ʼ�~�/װ��>�J��t,��N귅Կ�ŐÌ�U��P�������\�bf��e�K ����5�8m���me-u��`�l��C5AtGu���vĒ� ��"���%�U`ZnS�V��O'�������vU����G�*&�H�W�����Y��oN��M�`R}c3?@C��C�ۗ���w�2�Y�ː-��e�gz��ֲ��O�=�m��p�5����C�M��i��s!�<����>0'&��b4��b���ۣ�B��I)���>M"jE��Y��B��U#�=U���9�ƺ���7�1�%��xt{����JUM��,�9/�[���*��������\�����G/�k����������brg}��R�^9��[j�����P��� -�jSog�F�Z5���q��i��W��$���g�����,ܟ0R���l���3t)���������x[��Nc:����f�xO�ߧʝ�8��3+���Cl9�ۃ\%"�JCv��8���٬�<ս�}����b?��������������8dwuoD�RD6���۠F��SA}�����CP�&?�-�FV���o��i��bu��O~���ru�p�����6�-7��n~X����V�Jϭ�IU�[�b�5��3+��K�=�G)x@�/���}�&���
�S��BNQ��R�]V!�t��G�Ų/�p�%�mk���I�}�1f:)���0�E��H�~�$�O~����M�(��^�o�-��>~��r/�����_Gp�qm�f�;*<}�Wj�3�{�C��xf����-��̃~l9I����q��s����<moŇ��Z$�:Zv��T=H�8N�cCv;#�kǍ��1N�D��c� �w#�>Y�=,&�"�z��8�qz`�ʺ�vXD��Y�6�G�V�1�G���?�Ӣ��ʙ죍o5����5�Ϋ��&ÖR��^��r!��?�^�5��Vԉ�n�9}=1L$3��a|~�i���(�3Q�g���D���B?�~&��j`��3��b������o�?o���_�m��ʼ�_��_����v�9����9�P~9���͟������{�磽��J���f�I��K.ӟ��D��O���]�??g�ɟ���}���{��W���v�������m�*D�|�9d�R�,S����{�=�L��D�ae4{�٧���9�p��A��Ձ�3:���je��`�M��mR'���K�׳<���d+���F��fz�F[l]�UaZ�]�8v�~�n��3�nc���~�^��=�Wq}�k+�_vMt��?�����j7_P�}��3Ak�X�6�"��؅�AԻ-�AZ��I�H����.F��G	M�)��N�h��n�����U�M� ��
���̄�&�KO7�7w5:��wX�E���坌5�Ss��ő"��łr��bG���������8��m}�b������k��b}����E����/E��x�t��_��T��;��v�������ƾ�ɟ��~�/���s;�u�f?�3��Ћ]�Xj��-��o��n����B���by�[�O�~������^�`����ۤn�;�I&w�)dBO�L������p�
�Nws�;�
W�ܥi�����;�ocO��ڶ�Ezn(��,��~Yb�o\���v��4bҩ^���ㅞ����ڳʞ�������Y��(#Y��X��7m)�
W3dVH[��w��7
��~u���w�	gs�bMzh"w6�<r�߽b�ރ
���d�����*����F�VO.�8�Z�C7I�$wj�^�Oy�z���<�PQa3f�7��$�x������i���3y^�m�"����J^��4�y;����t\���)W�w痰�?�����H����\/r���$�ڼ��w#%��*�Sd7\��[�c�wo[L"��5�ߍ����~��c��LZ^�q�Usi�snc	� ؾ�-dwX9]�E3�z�s�AtW����W%��(�z����W���p��04,��G���k�8!������З��½�YbTv����_�b�(��\���n(����t��?}���{�W��?�>����j��7�v�6����o��aqi�ҍ�AS��tߗ��\O����H����,l,�v�_��r}Z��'n���OUh��k����a=ڇ������lO?��Wϸ���]?���d�������_��o��T�f��:���^�.0٫�����8�j~���=�����|!���=�l;�����Bv��N�y$������u���A�}~k���>�ojoG��_�;��o�0P�����/ܯ�ݞ��g���>o��r���W{����H��5���W�y�kA7�U��$��_���wY�_�����������|�����k������M����e�+�R��25����?�����T<�ף����^_>����/���_^���:k�������_f7����w����������Y_��g}����o_�����n��������loϿ�3?��ӝ��ȹ���g3/u}}2�m}�|6���/s}�z[wV�?���
�t�yO�����,���2�g�k�l��u���[_o������O��������Χɾ�����۵L�V�э��_��Χ���.�sr���˙Ocgj��wY���m��|�}>M��E���g��m�eΧ��f���;�8���aZ_Z��?����V���F���s���:�{��]v��uR�i}�i�宯?�~g���z�,�������������������#���u�t���'sL67�~y��in��Yv��5��^_��!�Ó=���������O{���4՛�?���O�����i�~��e���Ӎ��������.o}�5���g�y�sj7����iw'N�����)��Is��������S ޗ?�b�9��e�Sfz7�U���K�����?�z9�@�d��k���ߓ?0Ȼ?;���3��L�L`�$��)�"{5���si?����a?���~��J�k�Uw�'3��/���Z����2�Ղ�cWXk�	�<Ϛ�F\p�o����t���7�s�ɞ�oDS��f����D/�m.����m���n�"u�1ZϤˊ��j�M�IdW�:{�Iɔ���1����W>�.?�o�qnNE���֬�������"P��c���[�-�.㌪V&�W������3���U��Ư}��|Aj��y�6,wL�\��O�����R|��u���������[)n�o�%�$��T�2�ߪHV��o�z��75Q����s���t�������7����-=��?��|����w����S�Ͽ��1�����8C~�����w�e=���?��ʞ?�=�Ǳ>�O���M6�I�9��Ͽ��<�N���߉�����������S��Ͽ��z+��o�Mp;�Y�f:��i��y͞��ue���[j��9��I��o�0���¦��e�����ߊ�A��*��m]��TӺ>=�}]߳��6�㶮0�s]�e����ʳ?�z���i���[��-�+*�T/�q�?��ߪ�`�n�7�V��Kt��C��-����͚a�3rH�p,=bЉd�B���[w��ߴ����'��╏��wOx��g���K�M��ỽ��'��{B���x������w���w�x�n~*���U(?�Q��תr����	�RS�p�y�F~�!�uN��}�$���;ZZd����o���_����@��7�{:s�=��'�#����ԝ��Pj\���Q�����~�����EH�B���/e%Ȟ�ĪU��d{wFL�_Ț���5��t���z��%����I�ٵC��Ŭ�d*� ���U-��_@� ����m,�{�n'+�\� d��y��^V2{/ˇ�[�q<S�������c�j��a�M�:̉꧹�#%rN0��L�w�~�|�w/�ce�����c�/���f�c�r��4f�뒨������hO��L_�yz����{M�!rl7�sU��gJ�f�XOg��.�??;Z���L$���=��q����1��?�c>�4�2��8IdW�y�l��K���e���'���?|Y�c�?�>Vf���
��Ϳ>��ߟ��ݿ���X��~�Ǻv���_7F��>�����6t�߷XL����>��6�xy'+�]�y]:�P�U�ڇ��#�g�\��ױ�~��͌�MHm�'�*��Bwf�����zV��zV��7k뇨Q��?�3��c��{{�~V�H����X���w����~��CWO��b��[&��~�x+d*o��q�*�Ӷ�T�,ע����z��Z�qB�?c��bk�j�2���e�b���xvp���ty}��.�xc8]2}0�����L7,��������VJ�
�2��)��㲹����a�61���B�����?ݮls=�R<���iq���mV0�2a$�z��TIm�Pu�n������,��k���҇�����o_˿�[��eX���;���x��.��c)��:�n�`�#���5��d��H'׾��z�y}�+Ty�oX��>��a=�#�Q�\���G��dd�����H;�v�qr���ɬ���D�XY� W��_훬�!)�z��,��:��e�+���e?�Ng��0�ȍu�_6�c_�ֱƭ��O���ee��!��X� ת;��t(�}-�PB8�{�M��m(�,{V���̙7k��̈c�?zH��:��;��[������6���N_�=^'�`�����]]c(�5�Ҫ���ёi!�ImQ�
[C��ʴi7$��f���n����i����MFBBF���U$���c7U�g�/��� "�"�}57���l��SI��؊����r;$O'o��{���3���A�ML��n���~�#�=i�}��ٍ_�j�5)M	�M��S���}r��=:!�iv0U�`��Ȧ������)4���g}p6�la!�xe��
�_�A��Ҙ�ٔ���fkBʢ�|��Տ��#(%i"'�;Ä�)�X���Z���G7�e�����矜���쟜柜�l�O��O��O�j�F�?"&΄������b����J�.�\�V�qM����|A���5� ���H�)(µٌ�,ap][8���;�Б�T�Ƈ�iL@��C	l��h���P&���G,`�A�a�b�u1��/��&�0�B�)�S�7���s8/�o�V��I�ȄUj��<� �d����7��<B˜k;�C�����s�'C�N9��Vkf�P?��L��kqq-�u�ɞ�`�nL�`�{��X�:�V͎�V��R�²�j�Er}�$V��1������w��c,���hZ��k�ÒΑ��~¤սZ�.ݪ��G�fN溆��F�g������\��������w�����"K��r��v���y��V0��,�;M�j	A>F������%�uYV��{@D�Y�vX-�RIV��n!Ŵ���g_�v��Sѽ�3���g�E�O�E��`�0׿G�x�]#�V�����և��ÚF�["��ʒ��i��V��M�O�����;���m�R�#�b����{G�0攥�6Os7(�X�^�L��A:E�Tw/����6������(���.�l��Is�<���4�v�r>�?��uY�3�gu��������1u]δ��@缯�h���X�+o����^~�{�z����	��}�@����5�&�t�.hZ�,~�kZ�*~NkZ(~&5���8#�Mk���V��MkjC0�O��zJp�ivWc����I(�U���`M��o��@F�����s�6U7M��R���Ʃ�Î4~����� Gh���g�$5���u�
�L�{����g�%uӜ���Au_���֔���&{PSypS��7���/�Z���h��7��t+�v�G��ɣ�m
��3W����ΐ�6)����N�����PҊ!���l�s�驤��u9��ND�Bv��j==���	)l=}/՜���i0r'+�S��!N�s���Y�Ol�硇:�feoF�h����l������d�a�%�uI%w5;s`�;g�L��3��V�e͙���p#㺱�mѪ���[I7��%\[/7�l�L�F�ma��J�4{C㄰�)[�*}܏X�4�KI��74���oB8r`��|ʅ
��6?�[E֡,��oq޾�n���L�h;xc]�	�X7h7��F�tX�mwK��-�="ٛR2�g�Gܒe�duz�Ɣf�ގ�e3�ܦC)Ը��'��nhl��H<����	���l&,!�,�غ��UsY����$�5{s#�^��-M3#g�}�D�m�Z!���7��$׉$���0F:�|�Ҭe��1�CU��_O�y�m|JCȣtK%�_��4GҴcCI����a�VZ	���f�`��	a��=�a��e;�2H��C�TN�f���}'��F>�Qѫ�V+5W��q���V�tc8({?��7)��V�g��-�`�G�yK��
�����������>Cؖ���S��z5�t��������.�w�kM�{3E����e���AU�Q[��6���X'�k"�m�͌�f��~���r�Tg��r��3X�=Xv3���?��<�X�0X*<X�K����a�2��ˊ�Yng,�,/ʊ(t(tc�ci����b�HxЬ�F�Sbfa��&�0Lp+�!�|���Ɣ3�Rμg���r�.�,O�t�����||qG}�X៾RL�֍���Mli��$7�%��̒��6N�0�����,�3�� �j����*8:�{+w1���)��>)^Xס��l����m�kB]W���`���5�dZ�u)�O��� ؕ���JCʷ�+�m�K鲬m�ڇ�ip���N	��_R	W�B��J�b�Ѣ��Q�?DA1���WDA+�[V�FA���"�������D�
�e�G���
��
��d�c�R��R�
�pOV�aIw^�K��K�\Ǌ�`E݄T��`�@�V����hu`��-4@�.��|v(�{�7���8<T��5�]5�2�)���:#�<��Ϋ�R���FDe�`$����?zя��A��� ���y�u+�z��g�KN�b� �U;�JO�M3s���C8���U'\?7�i��<�PbbxTfHd�&�v���C���ټ,{�f�+�4�t
O�F���ײ����g����hS��3*{E�M��W���ɷ.�N{����|-��������ܕ�~��׻��A|�`_�̜�qj��<��ϋ�EJ��u';��A3g�U{h�y�`���gl��ѴD��v�_��/t�/q��Ow4Y�5Y�f�;f�wª�O)��ͭL��%$��7���=�}#V���DU�-bU���#BiuDN��i��D�o<�IS�S��SW��>�c%��rܝ�-������&V�7��?2�9�;�A�����y#��u���B*8h�>E��Q���t��Yf��-)���J� �w^n�b[qi�3�4�a���ʜ6GM�#�IIr�p9*�u�Q]\��-����:6gn^	�'5���Q@e.t8m�"�m��YTV��V�-a�ZF�D[������J�-�a�+�*-�--v�V�V�[�kYX\�܊�UK�N[Y�͹��a+)�%	m�|"]Y)~O����
�/ɭ���u�����+c�%�B�u�P�F+�K���s��(�e�h��X��K�$P\ɫ�!Iee�B�-2cz��aʢ���;KrK�9���Y�đR��(�b�I�չ%���V9�nQ&:J����>I�hZniA���rD�R���}�-2��9�>,z��HU�������څ��7��).�u��6�-���.Z@�W�/��^P3{A�I�]�f�m�w �!d"� � L=\@�
�JJʖR��4�T���!��jBB+BBЧ�_�"���]3�&�9��z�q�����Ќ�5����CBB�_P�#]�	�I��m�/T��G���V鬨�wB���Jt��?�x|�2�����elP��LCF�qj�́��P$�O��U��eN��2~����&j	%E�(�([J��D���W@wg9!׌��|�K��:^AÒr�*J|qi��)��y�`\̚\��/�Xxg^Eq��;g/wd ��
��9TE%r�t7��
���B)iE�3�/1%�#[7&7^��$҅�
Tc��F�ZL�,X�Tz��(�eV���R*��x�����i&,s��'(y�!RL�S�)AYY�#�i�+y��H6ߔ���IE��Z'ky��L$L��\r�Ԓ�\jY�RH�D�T9c��$�Uq�JV
�O�*YNř�.����%��*H)�Z"Eڹ��b�2L�eRia��5]�Hϭt�TT�U(U�\����k2�uuMŴ6��aw�d�
0�+�'��?�L#DN�$+�^�x���4�9lA�{}�@���J�c�$1Qtr�J�g�1���
Ga	��t�c���-�l5X��_���`jY�y�.,�-5�4i2�:�Ls,Ud�v�p�Q��`Vq(����eK��J��.q(�L~I4-+|�dѾ+,�d�z�R���NE��LRʡ�K*��d��U*|��#�²����M{��<���Q�!d����X��٦�R�AR��4����+��W&�K�*)��,2��
z��Y9NF,p�4����~j�`r�4� _����jL�$�U����G�Ԛ�q�27q�q�i�3lɉ3�N����f�+�YWf+��E���	wD��;�G�e�����8�'7?��H
��lI|J�ubj)��WUT�3y�T��[�&�HI�������o��IH����{�Ŏ�ۭ&m��&H��@�|��t�{Jo~�Hk�_I}��O��5�����=Og֖��w�>r��m��Xf�梧�����Jƨ��WO��0v=#�i�ܹ)�y{%���25[�S9�M{���1�P�n3G�e�9����0����c���r��9yڤـ����N�/���A�����YQ�Y���������b$�Ԙ�H�ns*3&;&:�^����]�M��̜9}�8����--r�ڜ��	�O�T�t6n�m�����b�7Dx�����l���ӐJ��`��J��Qu����ِJ�8�>���u;�k�7������5���&Q'�V��%�_>>dnEy����#�J��:�D����� xZE�Q�r���؉��w(�MУ}�GE(
U�Z�W��PB��' ��U��:��!w�T��B�E�ϯ(�$�W��ˁ��������ҲR�RUj���#�J��--e���`�R����5ZP��()��(峀�qOyJIavJQA��8��0��G{61^9ʋ�
m�آ�R+ujA	�'�!�d=��z	2-��B?�/F�y���+ߝ�m��d�~<��I1�̳������n���d/A������'��h2Ͻ���n����'U��?RշT�?Zn� K7Ѣ(��/�Y���[U�R�� �_��}Uu ن����jPE	�|�-�Y���i�[	<X3PU�ߕ��(EW�j`C��� n� �v���x�����V\00�ZUMlt����m���S�3�P``���X4HUs �n�}�~���������a��a�M�]�� [G�jp(�7JUc[��cU�0p'��vvR�]�sQ_�h�.@;`�h��x�f���;)~�� vR<`�('�� ���� ���"=`ীG�R�8��X�9Fnl<�9��|�$y�4��0`3`�t���N|�g� ïF�z X�	�X�����5�����9��	�� �l�H�J� �9�z�� �`�(.�,�l̈́�B�<�>_UÁF� �q O��f��,ȅ�}�/[���u��4��\�Y�iy�7`�r�|�Q�]�v��b�G�G �Jџ7 =`:�a����N��
��vFVB!=`,A����\V�~�,�\j0NnD�2U� <�\U�}��V@�)~%�nB�U��Q�@�j�3`����!�݌�:�0��lY�| # �� 5"�À[]cm�|03g>�v�>�r ]���G�nEy�S�q�K;� ��<�5�}
� ��c���i�x�� ��r��,�9`�O@l �,ڢ��C������'��y��e+�x0p(��3�`�6����ܾ��=��y�����z��D�����_E� [w�\��_b\��
vk�	����p�k(е���B��#��7��7�߀�{��ނ��#�۠,lx��۠��]{!�(��< ��^�5!���;P����(�&��`\���S�8@`�y�L���;`````:``�a�Z��#�#��0`+�y�����\{�
X�� ��C�����t�gE+J�v��0p�
�2�̀O�|�8ী�{��1�20��X��G��w���8�����G*J4`<�t�,�R��7� ���q�.��� �(�0�	��݀k�n��S�p�p>`P��<	�S�4�� K #��p1�.�m�GO���3�w)�,�d�Z�"�6���� ��;����ǀ��e/`4��퀖����# 7>�
�6�Q�/ � �8}�(w �N�|��u�̀����=��R��8E�
���/���倛����'�^�G��x�8�m,�|�`	`	�Z��_� ��3�8�00t��|��&��`��9�p0``*` �ŀ�� �_,�p�?[���8��0<^Q� � f���v���
��(�� � ˾@����q�Ӿ�^�\xp;���\�<	|��Wh/`�XsY��T,+�,7�1X:�Bg�w}skM��: xrHg`�r���oq+]�����?ԛ�QҀ���iu��L��Z��8tp߀���
]�_����5�x��&��6�n=�o@p�A�N�O{��&����E�\�7J��.Y'��� Z�[yS����a����yG'����C���,_�~�kU�E�u�$dw���GYOh�"�m��,���l�"�'_d�P[I���ʛ\���zԇ�;s}�u�!G�oxV��]/��Q�j�8�Ѿ����&�/�w�^� +t���<I���u��z;���9��tAL��^8}]����ټȤ�V�V&��k�?��&�L_g�%VV�͠o��m��4�.`�:�uJ?� �O\�b��'�ɖ!���Ft�|xVi�`���>`2tt6-�@��{H�70�n@,�|To��p�SqrV�"�/��x�ZX��,�Ѝ�����?�	�o4�d���&�Y��EA��O�kc����.�Q;>E�ĭ���3Q���~�_l���E���Bx��3H7��X>m�<�T���_���au�����o@XҾ��jp�!$?�:{#�ݢ'���A�i���x �^�������}O��Nw'����A�[2S����,ƖCc<�X����۬�CEz~%�A�e ��_�T	�������b]�U��Sq�~�1"�� _֭�%��9�TI�N��A-�$�D�i"���Z�Ux/[��=?B�ú�Q�ߡ�LխE\��g��us��Y�ާ�{Cm�������XJ����� �h��A�}�<yۉ^����/��7���'�Nz�(�w��T���;A��>���'}4�m��o���C��t�D�In�7���'�N�k��o���I�	z��=�A�
����G���z���4��A�*�/�F�u�>_R����O�@?~�<��'�6�y������ a7�R)�}�ZH���{\�6 '��<ӑ��9T��9��E��_�u�����"fa��s���PeÓ���$,��$09t �豪:Uجt6ǖ2}a׵����y�f���[1ei.V��3E���h,m�y-�'\�����G�A��~�L/5���r�3L�]����<;�3E��hk����s��=]nԣ���X3Hy������!�sƀ�$QO�;���]��i���h�W� Ϧ �}�l	�x�>槒*l�����j�S�q;w�G{����%���qIr*�6��$�	�:�Ж�=Z
�\�`��lacb|���.��3�e�>��"]�HG�ű���&�>����#_�� � �H����wt'���^׫�:�_�P�BO�������ï���c��E���I?S>	��N��ٔA?���)	�C�0����������60����<AU��ڽ> ��R��f���pߤ�����e�L2�1�C�笳��K4�mD2_F@��u�v�;&D�c��	Je�K���[��%�귺m!yc�`��'�>����ab�+=JV��O���y�թl}ԅ�����W�}me��m����22���=~�M&=�HC�|�{�u�g��n�����n$��
^w��<E�G�G�U�'���� .Sﻀ4��Z��I��H�<�}������v�)�4U���v��ހ�����@i���zYm�r�g8ѳT��_����̂B>�Jq6���2�W$�X�e!n�_�����7�Q�����YG�Cz��>ǰ�l!��}�!}�~
��¿�>*l�u�A�N?K��K��y����ߺZRf⏸0����?����?2OU���Sj�}���������"�/7�W��ւ��]�~��<$�������,�'
�d�OUCe~)�z����t�[}V�6Һ�ؾ`��������b�n�.<�����ukB�f�=�J>=�<��;"GU�m�bQ{�y\ 
��q������"�Z��>��w<�~9�E�¾�{R���gJ�b=V�e�@��<��~�B#�g
o��<�tY��z������'�M�ԋ���	�՘/T5J�+�$]H��gR�N��������a}׋C�-^�y�(T�5��,���K�C��<c�Nt!O�BU���3�q�x�68ɗ���,/R���,�8z���]���{�ȡT����o�T��W˺b���z�������o��.p��V��{����P�'���?�M[���D��$�u$��@ʥ���B9�t̫���E!���1��^ߺ����i����=W�T�=?���ϱn���<�"�媺׏>����M�H��¡S\\��Y}m��>5гzħȶ�>݆�l�.��p�=�ܬ�4Ͷ��m�Dٲ>-Ӎ�5�����<��
8Uu�I'�ǘӰ�w��vsե���m���RU��g^�b}۟��1?רj�?��+��>�O�t-���l_�r���\Z߀�?�>�}�<��%�s]t��A����c�!F�g�7@���>�@�A+��g$��Ŀ������<��~��Yս�CgS:V�|�D±l]}ic�ν��=v���ࡴ[��mͥ��q�=�P��N����~�N��\���:����r|��y����߱��c��e����� ���K�f�Mh���i#��/.�?�9v��1��N�Jy�$�c'
�M汓����0�G��M���n���{���3^�\Z��%��d�o�~}��Y�����A������݂u���&
��o����sȚ~��uhϷ������&�۳��;���I��z���%�������~a��$H����i	Ee*��t��K���vGK��g-�����q�"���RՏ���6oyN������]�/�?��Ƭ?��T����g7�)|�q�g���7!.q����tf�-n������wR�G����Z�q�hd,�gb��dC\�3b/_{� ��L��8�W����^��d��$��SDg8�w�dgmY<ڋn ���Y�y�f[��<� ͮg|?�9.�Qr���i�}?�/u��>`] �
1v�yYt�4�Y�p9/�!�4Ћ@Uϋ��σ�s����r�u>+���ύ���q͠�~��'9�N�0�����J�Ig�X��{�ኦ���q 8P��8��_+�g����q����A��~�������gг@��'��%F�7�+@��O��A��}�P޾�2�Tj?��I�?��8�������g�������7~ү ��_�A���o~��A��_�/�>:�|�_�A��z�_�k?����~п��^,�����������'�A6�H�@�c@Zg�K$.�S��[�3P�g>ga�$���-�mc<����x�<*�<���Űe�'�h�vA�5��>y��l�����>򧸠�9}�[W�:Ox����x���p�|��y�"���� x�x�J<{���7� O������'��s��O�s��!��'�9�z@��G�^�oy&��x�?�[v
�/=h}�s����F?�ӻ��-��d���/�����O=Z�W;[A��O;�������.B�w&�~�L_f�!�~?�/�,���ݫϝ��
�)�9��~�Cm:b9x\2����G0���[-x��l����8Ϫ��;�Mu�g�V�y<y��ϫ[�� O�<����V��%��<��3�*�L�o\��ݩ(�lS�I��N0t6��O����J�s���u�:����>��6��N���/��ޑ����:л3��;A����
g|���&<���[�ē	��/�C���_�gx�_�g?x�]���e�'8�}��.<�퇇�?��姟Z@������$�����w=
z*�Cdz�d�@�z�L������/�F�0�q��|��\G�L�k_�O4z�A�}�ƹ}>V����B�T�������w��R��w����Z�V�]��
���G3-&�`�(�^T�Jw��Ȱg���%�c�����o_��ڗ��]�1.����"�zd�8�v�<$���?x:^2��i��J���Ƹ��I<�[8L�2чy:)�j���iQ���eQn ��'�>H��)��Z��t�&u�}��pv�Tٌ|�sKl�͢��.���O�@����o�R�+ۃ0��1��Z�x��v�T�� ���������޲过.��EHE��P�P���I�m�"|�p
�B�E�a(�h�T�9����D؆�� �g��!�^��CF#�"�A(D�FX��$�6��>C8�p�w)�#E���0��a�����!�B8�л��"�FHE��P�P���I�m�"|�p
�Bo8�� E���0��a�v#D���9�� =�P���s
��!<��a7�A��N!�C�]��CF#�"�A(D�FX��$�6��>C8�p�7�5CF#�"�A(D�FX��$�6��>C8�p�7��5CF#�"�A(D�FX��$�6��>C8�p�w�#E���0��a�v#D��Bۻ?ڭ(M,�+8O�$�2a&B;�>��g�A�%?�^�o�ߚ��MN�(�C�=��H5�,��Հ֝����-�n�Cz�Y��4#�!i����u����=r�iQF!܏P7ӌ�����OLJg���WUꬺ3��4���;b̈Qw�T�ȘaW��˖8s� �i�J˜�K�F�U��Q\�0�(��HQ��)9tVpJ5�̈́d�V�(!>���ĩ�`w��p:j�He��\e��(��"w�#�����x��܊��e<��{Q~�D��|ׄ��Rx�y��ʈ��%ty���/zG�|�0]s�h/���#���(�Q�u�9�K��F!=ؓ�����?G��z^�E�_��pߎ�����y�Q?M��Ç#��BV�Q�U��
��X;�x(�ڦ�ӻJ}E���o��A�����L
���i|բ�俒La�9? �.档��*xWH|�U<�?7�ѿ�$>�)�lz����x(�\c�i�5K|]���y�������Bh�'�v�
�cZ�n�i2�|�N����&�%�L�e��; dB|�f��S�z��Q�}(���EI��ޣ�����G�e���c��w\��������	��(�� �k��[���K�_��~��.��"�@�T����x{e>J�V
~mQ��Z�}�㲯[~�_X����l&��+N�y�a��K�	�p�j��u<S��S�,�o�m�q�A%6F9ޗ��E�9t���U7[�Kȴ�
^?� �	��0H��q>��oi�@3t�J3u�*�t��\�C�_�+֦�|�j~a [�r������:S?*߰��}_�	f-tI8�谄�:�U��\�����p��8*�1��!���g���>z�o���K8�6H�t��C'{�)�왝ğ����mN�=Z�i?'A)t����ߢv���Z	����H8�y��{��D��'����M�_��I8�#H�pz��.���V��������b��}��{:V����p���	�����۝pe���o�{���i��,�x�`<Ԙl�7��n�Sn�7��n�;n�	�	,�M���9��7��x��_��m4p+LT����#���^	��`�a��$�:�[$�&�>����"�GK�d2�|$��G|��G<�N	O$\�O��J��O�S}��f�����$<�ʗ��5^�E�K�O�ʯ��e$zp�T���9����q�N��*���O8�G��S4H8�G��StI8�G�&��/�O/�p���E~X·Q�N�5S���$��N�	x���Ŀ�����$����2��P{%�����W��D���/H�R��4>$��	�-�[��C�y���l���x�3�K*�j�5���B�1�Otç��s�p�^M��`=L�
ٳ� �n,��Nk�[�*ݻ|����M�N����	��ܑ�h��#pZ�O��&��F�	�z!pZ�k�Ձ|O#A�� �=��{��~K�����b����Ѿ�V�ۀ��V�t�oH����I�S�i�E��׽�^�F� N�2Z��������p�W���=2C$�8���-�紃���^w�o��M�ʇn�?��_��]���X��H���>f������N{#��7�<8�u����I�>8틌xp�#���̭����ϲ0O��'�[��	����J�o���F�.�3,�Z����p�!/���I8ٿ�N�G���6K��6O��>�-�d��K8��ۤ�ɞ�H8��{%���X	Ē�ǳ�/�$| pU¯n������ ���
2��XA��i���:-HQ�$|���p�[�
����	o�k5�-����t+���UU�����[���	?	<u���o�'K��'Jx_,��K����$���f�Ÿ���j2�i?���Pef_������z(�k�T%�uP��\&�?�F��k��,XOm�k��h'�ɾ����?���4�������>~�t[�\	�8�C�FW������ѻ�oQr�Z%���٦�uѯ��=��'<x(y���9�C���;�('�0�C|���o�:h�/߂��_A�����9K�7U6ɢ�!� ��j6���A�.���tve���r�N�tࡷX�(�%𶷌��o^�(7
��DoQ��$�%�9�,l'���Ry��%����*���H��&Xغ���|��I�߂%���d൐�*��lQ�E}���'[�ʛ�g�s)�������Wt7�$��`C>6�3������_�yǿ���������I�{_�[�{'�ϸ����sB,�)A���ޅ2p�7�\��n� �g�o��wT��+z}���ܟ | ��3�~�t��&�$ੰ���	|�T~� s�����)�5|?���x�;|��n��I�? O8�e������+B�̱��uc�9����,����9���������3�?�1$�x�z~/)ᇁ��eQ���Kw����� j����t��>�m~7�/�D����J���w�	w�a����oL0���;�+z���tϖ1�5�_(��2�<`ثp��^���m|����܉�X$���;%�����/�W|�D����%|�$��E[l����[��yl���Nӽ)�,J�("��/��^;���Q���m�G&�x�x�^�y�A�cD��� ��dÞ��Js}�Ɵ����-�P�}A���&k�{�����N�?�*c?�J�
ep��2O�O���_J���}�D�]eQR�[�OÿZ 迹��"0��7��{v#����x�)�7x�VE�/�'�o5ڟA�,��O�q^$������c�'�p���ہ�~���� ����?�o H�?��ߝ���П3��5W�]\��w/���`2p����t�!�Z��O���N�����"��!�x'�W�>�R���<ΰ�QJ�O��������k�.!���ϐ�E�~��s�����#N���������Џ/���^�bb�����"<�]��g1O�� �q�!���|DQ��/�w ok��{ʿN�����.p�����pb�	�w�������_{5#��7��D�����> <�V�~��o���J�F���V	���=������g�u_����J�.��m!���?�U��%�}���[<�!������G�OI1�ً�����ڷ����'��<`a�F��p�~E����A��Q��鎉W�#��Ɇ}�q�Y��ۇ[��r��$_��&ᒿ���t�2Q����;|g;~J�s�OJ��u�Ij�5���l��EwJ�S�?0Ű���%�R�����%�)�mg��{�p��}�9������No��Q?ZLnB}4$������!���T�;�[t*x�4�W o��?e�2�zI�2�L�/ �	4族����s
x����|c��c�0�Y �o����|[
�߉����i>�D�E�}�Fs����n�K�^0���=~�Ο��Y��z߄6K�ɕ��f�n �vg
ѥ���q��T �/�=�Pi~{�I?���\���G/�=���Y��ρwJ��i*����A�бR��QG�`K\�����1���;��~�K��ß�������[����s���1��*�w�X�|��T�/����)\9��͌_�y?3��=p�`�����7c=��6����<t�E￟?.�GwS~���\iȋ^<�U�7�ޢ({���7w�d��q���~��lQ��<��o�`yP�?,�N<N����?�n{v����'��(	�
�}�E��1��:��L�m6�'5�~j�O4_+�����J�|;�-�k�.��C�0�'�`y����N��&1��"\ҏI�#%�D��7_e��~���`~^ @໨!7����f�~���|g��?�c!��L����	�����c�a�������)�	����Ծ��^�'�J��
�I���p��چ`~Ch����)~A�ץ�OJ�?|��=�f����g��� �K�ۇ���?T��7��L'��Ѣ?���pA�|�2E�B�WF���狘�_!���~���O(�s���oA�<d��#�,��k�����y��o�K}��_t�����3��I����n����%k��a/D��.�Z���k}����S~���[�Ӄ����~q6���x���	܆�Z�s"��"-!�;�wIx-���=������Iߨ2��,��Q}o6��x���|�H��1��������4c��|���N�l�a_�� �_��+�eQ�Z�R����a����o�ח�{��f� ��%{8xοa3D�〗H�g ���]�x{��7�?�?�(��{�4�裰ך=�)��=M���N����+��<l��X�	)�x1��%��H�x���3�<���Cc?�xg����'񓾝 �.�	|�����N��i���(��R�Ch#�̃��I����)����,��DC� ���UE����+�$���7�d��C����Ͽ��`?���Qp�C?o�o�I��>H���.�v�[��I5�:��mn?��g��_J�w�wF[�/�_�0��l�7D�cȣ�:*iQ�j�i#��=x�F��OX�(�^
��Jw?��H�aO_a��R��|�5.��������?ʰ�W�I�����G4p�5��4x�Z~��5��J��#z��i�f�_�4����`��}����w�i}���T�[���(�	�$���;3�\����1����1=�]�������A����)��M���H7����~�w����o�;���8�:jT�KiG�F��,&v$�;���e�h�wK������b�w���<��9��9:��ey�fy�fy���W8+�U�������I3��'����V
��ŕNGE�sIv~IY��R���]P����,/�$��YVQ��[U��-)/q8#FS�2e���Ίe
%��jɒeH"a��{�������8�}-��O*/7���J��}X�����DG���8����c%�}fJFƼ���Ӓ2&M���="v�]$@���NB�N�!Yǐ�cH�1�C�1��z�u�U��/��9�2�����L�0��hUM*[�����!�CyŰ1�d
�����L�+��Ō��g��#YF�&�����#Yڑ,�(���-fo�(E��=�53w�\gq�#��binE�&k�2�������f;�KH��JQ��[^,a����+���KK�k�FK1��[T����t�˭X8��K䄲��ؤ��
��YEe^�H/+]�=�;%��,�K6�eUy%�MA�����Ơ�����ť�Ff�V:�I�;��D�^R�]4�x4A�����I�?I�ؼ4mai������qL^[���yL>��53���Nv^n��mD�(S�<�(=�ڑ+����Ư��eK|��Qca���[��dGanU�3�fA���G�](�"�YT\ɘY�h	O&�[�����GniU����l�d�8�K�*�ޢY�Lk<H�By'��a��ƒ)��,�]d��Q[%��NN�(�*]�]���$BT�O%��ܨE�E;qۙ�cm'�xǙ�Ͷ�4d�.�����		,a�Lwb;F\�ǹ���ׯIy��f�����U��`�oл��V���q��Qɖ�(�;(|�F�le�_�
��r�.үؘ�Y����J���ǁ�����_��t�ډ��eY���D��z�o����-f!�5쮃��/9 X��v�H�*S�`�D�����f��O��Ҭq��]��v�z��E<_<�	ߒ�)��Ho�(j�*Af��m��R�UR�����Wmߪ]}"��S���Ů-�x"6�ۢ���\ �p~��SORtC�]{ �=�Rf�,��L�M#�,2h�,����XU	�����[_�,���<W����"����y�8�5���������b)~�rX�[���])�O4�����5f��Ů5�6CDČ��{��cڭ�����eq�D#���,�����Y<��xu�N�ֶ{1:����B���',��߄�B�A��r]=�6�z�)6�Y�)�gB����B̲B�-R�����Ęٹ:/�E}¼��U!�l�	�MQ�˺z���m�:�������ǘI>�Z	�Q��0�!���T&tQT�s{5-X���R���9c7K�UP�\�hǏC��B��t!�,�fҐ���󐑒���8XS��a�v�ưGX��̕efx�@�ߥk2Z5څ.��'.{�,��q�� ��B~>%�[�tٽ|��Lz#�_6���)m\#�/� �� �D�(~��G�En�G9�ۘ1��6���L�]F/�-�D!�U�,`�dL�nv/_�a���=ʖ����铄�R�"���z�V^����j&q0�.���4�Oa#,�INܳ6IӀ����%"$q�էB
��͛ة�f�{�v� 1���T7U������/L�$���������z�ce�(G���'�3:Ŗ�֥|ę+�d�۟BK� ������~��"Saاt����Q��G|t͸�3gn:�b�S~�^ul x#_Q�KiPþ�v0�rF�j_��I ¶D5��@P�z�'�*kX$��VgU�.w�a	cF^,,�0��n���a�D#/m���-Ǟ��c�a߲���-�������?C'���4L�����q�e:���Θ�r(��`P���@��}�%�	����;�U������p ���`��Dɫ�5"z9��7m�bP0T-8yn����l�����%�閇�c�yX�}q=���B��K')!V�<g_~ǆ�S�%�Եhk8��K�L�ܣb��� ����4?��<E�ǽ+w�� �����u,����+Y5�3�a�|�uk�"�g�)=��V��.5
��3᦬��a����Ɣ��i�,X�D�(���͇Mþ�ʋ?�}N�&����(Sh��:L�� tT��Zѭ9B�Mx
a��D�� �T��������c���3n��0��a����`�u(|���ĝ�F"�՝z�#���$_W"(�i���)�)4� �EͱS��A��(�gY+�����<�~A�ݦ�<
nk�C!�dr�Ea� 7�a��l	�8=��(}�����ĬR=��"�}���N��(�M_e��kF�3bL��v���`&i�Ow�Z�C�C�v���V~��8�r��X<W��"���JN��[/
by�@,�A<���JU���U�)H��!t�7�Lt8$��|�5b�@t��OON)�"��Pj1! b���.��~ջ���y�pꁒ����tS�����lh��̓�,�*`{h� �㚲V�-��xT9Z;�;�c�� �����?"��� ��!�;e�gԛT������o!d�V5�i�`:� ��]���U�A���jz�:��KzbI�r"vW�K�Bpx�q��"��� �|v�7���z�ԙ1�B�s��k��ߚR��tM�����p�\7^^�F�7[�h�{�	@��{\�A��g�uH�s���
�Ñ�'�e|>���� �(vJq�_�~#f�ٍ�/���toV��r�f��4�>J|H��y��Г����<k��di��z�����9����
������7&�$�jy�X�{"m�uz+J�����B�L��y�4  /?�&����9�vKž��`��	����]%E��}��H�F �/�F�ž8����<��̮t?�A8,q��8��<n��l%��SyT��:���u�l�90i�s3Fأ���{q�4Fn�NF9��\��hW�!���tt���p��=�"�
UĹl�;���p��?�h&?�(j�>c�a�fΆh��]<����`,G}L��t����r�:�g�u6%� XO�W�N��^���٫��TB?Ų�K��Xr��&����]H�*swP����E�م^�0M���,(\�5δ4$�VB�0]�r�<��J�v�C�@u�[-�O�\��g �}Ǟ��,ӽq,��.�RD���H�=�ȓtL���I�����,	��G���4It���
,����9�X��q�ā+A��D曮͊=����dO�T�J�S�^A�GWe�F��-���.{��G&П�:�5��
ƺL�$-:S����w9B� ��1���#!w�4�c�`-�2r?ˠ��JN�J)�0���ۨ�8�3��e��L��T��?�^ex �}@Q�*m~N�y`To�1�8�%��7��Y����"m] �	�)�>;�P�u�ċr�e��g�Q��4�}M��(�A�PK
    +Q�HG<	9�  �� #  org/bridj/lib/sunos_x64/libbridj.so  ��     9�      �}`T���"D�&h����m��Cm�b����|X�AĊ�H���l 4��f��FA���iK���Ɗ���HT�y4jj�n�X)�"y�3s����l�����^�����93s��{���>����z���'��y<c@�U�O�'�3��5P;�����u� �ī�$	���H�x��x�������i\�Ni�^�����J���8[��_���ʸ�d;��������PЦ=�c��p�g�4��P����2o��+=��@[����U�}ϡ�����=�~P���5���ܣ$���չPݏ)��=)�K�t��Uݿϑ��֏BN�@x�����?�iCΟ�X�����q�?ݎd}O^���t?�֘�%O9�,��+}'_Nv�!�#�f���+�Nw����u\�����L\�p��st�Msq}Wߏq��=��<}?NS��GF�<\pM4�&i
Q�L�5U�5���"\k\誷ȸ��OpA�<sp]�Ë=�ؿy�Jq��������rM����T�pU�F����U��b\Kp]������q݄�f\A\��n�in��e�Z��v#��4m�u'�ߥ��5��/����~��׸�3�j��[W�~��~W�\��'\��3���js�{��g�y�z\pm��(�ǌ�a\O��b���ڦ���y\;p��H����\/�ډk�{E�Wq�v�͸����������F�nM��4������ڋ�F�5���#\�������?��9�/p��o'4֓!\�q�u�����+�pv艸2q���4>�+�N�8�k���+�:�Lг��٠���6�\\��5��p}�h���p����z�����y�o�O�M�j�O���q��W�K��"���5�e�r��s4�BSlq�\W����|П���P�q���u�Z\�t���t)�p݈�^��ڀ��-:,��r�f\�k�3��Mw�~��w����݈�׽�~��Օ�w��qݏ�:n-�Sn�������I��0�N�t��_5��*相�0�Y����PC<����6�|Ǹ?W��a?�u����������i��X�|#� �\���i���u)��qʾKp]'�����V�Ig�4]d�]��:/���8�\�I�ی�fW�;����ޭ�*M����7��j\�����tm�2�:H����6�zד����]���U�o��l��^t�5�_W��3AYo����G��4퉓�����߸�Ը?�,/ր$�$kj2)�z��V���]�G�I�N�5Bǝg���+����q?ʸ�܏��-#,Ǹ���?7��v~���:|"�$}?ٕ�B�������-4�/u�q��5�����p��U�î6�*]e��θ_��k5�^�e��7it��
ܤ�n��+�D�
W�ρW�_��҈�5����7��5�~�� ]����'}�� �0��=���.��´��oP8	;�����p�׹��.�҅���[\�Y�����.|�7����	�P�N�����e`�t&��)SyS�qm>W�L<^��s�:��R�����x�'ј�28F���C���m��S5�bz(��k�����4����e}F��̏I>K����d�a�������n�2�Z་��j����b�����C�@A��L.u�J^��ˉ1���U������j�<#������>�,�������ۀ�����?p�C.���Ï���y�w�Q����9��ۢt����������`��4D�r��'��G|'��Ug(��`q�$~�z����e��w=��d��ݸ4I΅�Cܭ7�t�����S6�_ܶI�]��uP�C?	ܾ�)o+�cC����;�����q�P�7����Fu>����]�y���|�%N�.ny���b��F��1��k�R���7��P��.�Eb��l�;��`��R�xp��gi�	�2��_6�H�����gzJl���>Pv<���WlV�U����q;�R��݌G�������>��~�}���������өG#�ێ�L�e��J�>��1�Fރ��(�o����_�x�W燧y�j�w3�C����{8�g~���Pb����	\��:�$AF�~����}�:e}? n�>I��#׌cb��1�|]\�r�����[�?��>E�gY���,��=���<�>�Gk�9ؘÁ�Z<��t��n2�>p�ϩo2�Z��_�g.p�Pg=���W�s=�/7��
6��ސ�6�6c�w�`�W��w׷�3boj,?S�������n0��W=c`�����X <�Ot~�\������g��������6��N6�{���!��*�q��Ƴ��soVgG�\o俀�|�+�|�6��p������o:����gÇdx6�nQ�ی����:�����Lp��m�%F�0��r���c�������;x�lg����Y1�%�}���b�b����y?�O��9M� p�1on{H��|�2����A�{I�8ň��x��f��.�i(���'sxG=# ��}�|]\���߫���U������o�3�������6�ۋ����腿�9:�ip��zqYz����?04_��o6�)_M,�>u��{������+�S�|֧�qo^c��eWy�1�������R�I�i�k��}m�zF�)�i�3��oR��L�������a����b��+�n�h�����x>�ޥ���C?�ǫӿ����e�Vg��7�v#>�n1�2�vuf������3~Na���]Zʀ���--��	���_X)�:��/Y}/��B�~�8k�W��o��bک�?X�;���x�NyY������[��ݞ�z:�m�W����,�:�G��3���M'���9�sNⷀW��o�MN�A�d�Ӏ�"�~18��<��1�-���x.p�}����	�.c?�-p��������~�p�7��:<�h�	'A����z��
p���N�����`p�	�z���)G߼����֟����8p�Deo�~����w��!�7��['��\�\=~��+�;����v��_ ��A��?h����]�=C<[�ײ�����pG�����=u�1ܩ<p�����v��j�op�Z���.0��A������k�kO���눯��z���^�o��)p�S���X�چ8�kpG�W�܉gdƖ?x.��t|1p�yi�2�w3��N��>���ɧ��,g=�p�1>����Ny?.�f���O���8��[���,�����/w��ߝ�<S�Uv-p�Ց:�,?E|��/���lP�͈�`��m�op����*��3t����ݙ�Ӂ;f:���Sc�/9��Ƽ���70�ǽ������0�g���	��y�����jw��l������Ɛ�T(B�=���]���^�ǚe�9y��x� \`���͜_��I�|����s��~� p��L��E��	���x����0�}U��bo W��$�T��Y�]��X=R������=���}�]�?�{C=�'^�������]�̟��[���9�����ӿO��u�;Yk�w,p��{q
p���]�s��~[�݈�2��0�,�QG���r��O��Vg���*��I'���s��W����~��<��g �����w���n�5�]��gI�_bc>]��m�W������_8���ӑ>���w�[g8���I�#F�?�h�_X�Z���<I�:�G���?�? g�=���p�[�w`����/3�Q��l�ao|<�\?��o��_cďn��د�K���
#}9���7*O˲b�8o�}�p��bz��Q���ot������s�o�R������b{�9��(0&����.�q���0?:f8��e_�B��Ӝ�x=pkP�'D|'p�y~�e���n٧�5�� �3���3�~��?�w-������9�5
x�Q_p�w��k������ov��#���g�>?�0��$��_�y���pk�zo��4$g���u��O ���]o��:�����	��s^�ʎ���sp�G����{_� 8�9��8%;v|N�2���W��w.p������ħc��Z������ay���������P��[����y�J�ov��
�c��8�/���w��mg�R���},���{-뛱�98����Ψ�G�ᵎ�Q��_�����E|�Ӟu���8����9'9���L?�/��f���p���}�����5��K����u�M���Z~b���<�������3b��r����d�6�s.p���/7��l�VC>�����6�MF��0}tV��m��F�~��G�mo��/��h��:��7�[~����y�g����YF���/v��"��w����w�;�wkX�J�L��[�����+,�lg�K����gg��2�����<��Ӝ��)p������r%�>#�������u�wtY^�7��k��#��c�q��R�?�O��~�;������G�7�O.��߹�_zv,�� �2��*�snQ�n��V�_uUMy�Oϩ��̫	��S�YTRQWV���%��cPm�n�|��V/�������4PUS[\R��3��daYqi��z&�TT\U2��%��e5�3�������͒yeՁ�J��u��x亂RVYVS>�E%��޾�X�paU%.�h�-�(	̯�Y��KJ_T(_T6��fqIM�]�
�5e%�ӫ�T �+Xd鵕�(.�.7�Y��J���⚲ڲ@�ߋV�����)�_R0�KjL�t�/��;l����I
��+e5��1�����+�JܭE���J���F��}�_S�Z��A��3�U5qZ=�_����*)b��~Q3Md7o�Dvk��f��!^��i����(^��i�5�ibfJ�U%�e��YT6��
�$�:wŵ�.��w5��/����;����D������JbiO�Uٌ���o�u�&�U5�x��*7/��a���8�jIa�²Bpg<�\:��U���fA����X���*�,epa�D{驍�n֍�ydniymUMiYMYi���g�˯�)��6^�²����VLoO����T-#f[L./�(�VZ���&PWR1���l	:?�^敖ͫ�Wb�Ӕ��.���"1��2u,�ho��������?.��#�u55e�c��T(э�UU���xᔊ����LO��5X��{��8M~��Q ��,��~�i��H�H�4���H1qd�jς�,nw�����
�`E|�|;d�x�Ċ��Z�d�5�-��������b2x�8���(���)��WQ���L�,��7��X�ƪ��-�*!��."�
������Mc�(��4��fn��P�%l��D Ŏ�G)�XXe��ι�T`o�F�sW�w�5�+�U��r�#^j�*ʰ�q5,+����U1+�V9�J�PT�.��󫰌,f��V�%5��
����_WV��H�`�M�D�P;-A�8(���щ�FZ�+Z����Jp�P�X�+cs��WՖz��A�8)�2{BI@G.�ʧ�M)Ֆ��<tu�˱�5��3�V�"��\3Â��]D����\r�Dߤ�K|�ӧ]���S|Ņ�'L�'Z���y(ZՍΓ��Ŭ ���6O�����f�~O�xIY��������[���xj5��fPA�#ƺ��3���D��8�ȉ�^TWQQV:��|A%�N�W]YJ1�e���\=Ev�K���]�����\tEB?j���Q���j�O�NAYY���h�@	l�K��B�#�JR�-_P���p�� 8�]�h�+Ou@v iZuټ����-�nPS�PoF����X�z�w��v��x��'��^|���3}���U^e+%w�����U�e�ն��6b�Ɨ�T#�̫˫W�$���-��,2�l�{l�\�4�TV;��\L:��G��J�%J�e���'Q�0ۃ��h6���̉�谘��:����������`��}l�E(�O�b�x~q�b�����@ƅ,���Uں��0�h�U�bC��Ճ�Sd��)Z��,�z'�>�Fg0��@Iii�V^�RZ1����̃��~-�[����U@吕ɣVG%��\`L���0J㤙YV1_�L&�������X!�� ]��*��מA���`��y�Tm�:r8�`�S���	�m��ئ���u��@��L���sI]ee	 ��
kJ�EF���nA36�8�7��}�j16�%�A�$��L����;��"�p�q�}�xAy-ou�U%N,�Z�^M�_SM���*���!6�J+� $��>G±xi*��n�1˥���~l�#� �Q۪��l�E�͔Ԟ��a:	�?�ޘG��RYZ	�n?��O��?��fbIuɼ�@\����Y]J�/��s�ث�=�mU�ul��B���Z��s�w+Y���.���>l;��尋Ju���|>W��j* �E��K�G���,�pQ�%z
�:\fn��b7����Ųl���ڜ���~uٵZ/�,\XRml��֛P^0G��a���ʰ*C#Dr��#��m���G�'6� IWcE����G� �/5�p�k�>�fJA�w/��x^-�^/�jl�~V69�ъ�"j	t�D��/Y�fy~Iu5LTꒉV]C��Y唖 �hB{&�L�5m	'��R[�oF� ��F�Z�z��@�Z(�^t�y�']v���iY�4)������\8U�L��9vrvr'6�t�z9K�wI(�I��WL6*�Urn�X45u�:8�]��jK���[��zh�W.RSE:&v�qno�Qvs�/z�6�r������1���d왔:ȉهE�5C���U��)�2i��I��ʺ��Y�3,�ĩ�_cg���\v�XP�Rgkr^+��8^��i�.��\R� ���5+�&R�%a�<ы��-�'�4ڵj8c���5U����.�d<���A�$��hu	��Z��G9h�R�_�J�VQH+׳Թ�@{�f�]@�%�(����!�,�9���ҳ@�4�.�V�a��W湤�6PUSf�$���4���s����Y� �Ĩ�<�q3�WϞ�J�G��tթ���1qu�W��m��pŽt��݇c��M!M���ϧ���)#��.%!3��.P<7>�X<�~�7Y.�����У�me>/(.+UOj��Tt}�L�or���Y�,q�-�Z;���iG5��$���2)��qG�3i}��0M����l��xbh�X���0�^8J1�j��5�S

���$�\9�f��4�J~D�;f�ge�Sm�ʑ�m�3�aU���:��"5�����Gfj=lk�g
q����F,�n��S�j̰ �wuaM	���b�l�y睧wW�}�|L�}
-+�-�H���S���a�4�j��O�(QiD��|�%"e�		M�����kБ<N������D���-��|mR���m���1���x�����HiTES�WD+M$���.�K��0&�a��@�����J�F��S���~��Zݎd�93bF������
7���ch��$gɏ��+w���ʲ�Z7��)����|���.�)��~qn��a5O���5��U�p�?��0L�A�#;3"U?�GE���YO��t$/����������1�\�s�a(5��Jh��1���I�=Y�J�X.�	k/�1Oj�m]t��ڽ�C�#24bW��RO�Qk���lU�5�����Uŋ�jj�̮��p=�[X{�C�����Ω�:'�3��K�s�9���������o�~���Q?<�o���l3���.͑��O�2�E����y���z�z��ܞ���{�Ipd��O8?�S��J�O�o�O�t6�g2��&�/}���*?��M?���D���Ы��ү'�#?��M}BӇ�0>�U����4���f����w�c�5��oM_��I��6��;�Ϙ~w�;p#�7p=�U߲���ҟ4}-�1}��g"�����o����6�O�>���x�W��`� �?Q�e\�U�n�m
���(�/��	�/�O�u^廒���+��$��*��oz�_ �E��b�ԥol�:��L�KHW^�W�%��M���~�߄�O5}[��;^��}Kӯ}j��'�m��o�Ц/c����U>i��!�J��}3�w%}5��*}M�h�Y�?E~D�����U���c�����2����:�����j�I����q~#K?��!M����N��LH������ox�W�J��*���J߃���ϳ��*���SL_��~��$��*�f���o4��s�W���l��/f�ڦ�n��om)w^姛�Z�#���^�#����M�����W�㤏K�Z����K��Y^��e���J�����*?�N?������g��.雔���7�ǫ� ���^�o��kwy��t���?W�;��U�z��Q>.鯓�^^�*?��O��;���%�_�{7���T���N�������e�7�������N����� ��J߽�mO_��e��Q����	��/ۿ`�_�7Z��e�~��^���E飔~<�3���雝>���8��ӿ}���-��F��w�瑾G���]~�O_��sN_��QN����L��mE��3��W���o��U�S�ߚ���ߘ~��tC������XMx��Z�,�_ܷ��o~+M������W}�F��^�;�~��ӛ���/?��?�U��鳛��鳞>c�Q>��?���s�ok��:���ݫ~o �Q>��ڐ>��s�>��c�^�g��h�;D�R��}~s��p�˘��Jp=�U>���~�ۼ�79���'H�� ���2�Or~H��^���@��]����Y�\��y��?j���x���Oh���o� }���^�ϟ���ߝ>@��/}��w�+�>��]&���jZ�i��M�h�T�zM4m�t��aM�5ݡi���4ݭi��]�vk�t���SA���hMs4��XM�i���$M�j:]�BMgk:Gӹ��j�״B�jM�.Ѵ^�M�kڢ�JMWiz������t��k5]��FM7iִ]���дC�]��ִK�nM�jڧ�>MhzPS���&k��i��y�N�t���j:[�9��մTS����j�Zӵ��i�NӍ�n�4�i���5ݡ)�5J4M�4U�tM34��t��Y�fk:J�њ�h:Fӱ���t��$�PXb��������P�.Ŧ�GJ�5�沋4I�Q�p�bc�@��25�i��ٚ��t��9���t���wCs0?�@sQ16�6���<�)��L�&��b�C
e1��c~h�T�zM4m�t��-���t���Y����,����vR,�y���L�p7�g6�\���u5)Ց����ca�{�`m�t�u�6i�t�����4��Pl7�b�� �2VO��p˻	�IӃ�z�S4Y�MS5M�4C�LMW��P��|(�H�8Nb8�jblLRl��ؼJ�l��P(���a1��F
)�R(c���R�o;����50~+�)6܃�FM����a�,%�ⱋ|�&�[�NM�4��4��^M�4ݧ�;˅2�����#�Һ��R���L�2���^O!)����c��U�ޫi���5]��ZM�4]��FM�Y.��,��(�J|�%������p(�~��^O'�#q51�R�o{=�I� �%�AT�t��z��<(&�C�)$�25��wC��c:(�sH���e<���l�� á�`z���
�F���9��F�Zb(�ݔc#��P)��q��y="�h/�ø���`8-e8��v�C�S7��.��w&�Qׅz�AN#������>�h7)�σ�Tz��dR�)�P0SI� f��`�$�1:��\)�lRS�Ha,�&���C
�)�䱤0�Ǒ�X�#��'�^�T)�)�R���P�f�� *%�a�'�qTA
����`=)���z�C�PZ���x\I
#m�w�O�Bo%����RkI��:NJ�ؤ0B6�By�D:�U;)��'z=;�~��C��yM
ex7)��.RU��cR��Ha� ��z���b��/R�)�0jSIa����hɐp�)����?žD
4�F�(�	X�Ha|��@C
cg,�q�SR�y�0������Nz)Ƈ���0�Y���~J�0oIa\T��k �q�$�`ޒh!�ºD
㨕��j�5XWH���%���@
�u)����0`6�^�q!���Nzƅt�a�?b�!����F�̯a0�w���)��.ҵ�w�wa~��x��8�#������g�c�Hi@c��a�L
5���~5IaLf���F
�{$)��,�V��h��7��?��c���c�"�	ƍ4�yF��<#��<�����lR^���4�F�RR����a�H�����h_.�?RS��>=���j�b�+R��I��8�� � ]�q ��I�ǾGz�Oz,�%ҩ�/�w{={Ia���NúI��R�Ii�a}�1�Fx
)��T� �O
C/�4	|%�'�J
#r)�������w����d���Տ���d����T>�L��S?��	橅��zZ�����������?=��y���CO�`����
�E�����	��flO�`F�i����wU�\�,�L�g�z������`f�󸡧�1O�����,��$�̓=��_0������	��U�/�U��H�����&�̪�����˅���_0���.���]��_0���-��S��_0��H��W
�}��l������6�u	^'�O�!x��?qX�&�6��2�ĭ������!�O\/�CƟ�Z�.⹂w���o���	��'��-�O�%8"�O�.x��?�Gp��?q�A�}2���d������K��U�U���'��_0Y�_#�L��ۤ���:�F�`������<��o������`>���&k�]��<%�G����j��_0O�������~>}���S*
q�`�?�8,�'��L�6�q�`���G��P�s����,q�`�?�x�`�*���P�����?�8G0��?�8K0���'N�D5�G0��V,��1������9��&�`���[���W��K��+�/��N�_�/x����_�&�ఌ��_p����_p����_�.���2����2���]2����2���Oe���a���'��'�O�OƟ�M��V�e��[S��9������W.%�#�+�U��N%. �̦�g�� �O�d	f��t�ؓ.x$q5�G0��_B�w@�q��_0��o��M�"�̮�WI��!n��f��k�����I���������������_�t��`�¿[�/���K�/���G�����I��U���O������%���w� N'g�	&+�Yĭ���"n�@�C\/����%�L�z�<⹂W��^#�O�'x��?q��6�,��d���o��'��$�Oܷ_柌��_�����]2����e������K����&����������d���_p*q��_0�¿[�/8��K�/�C�H��$���P�H��-�OL�=]�9t�����ӉÂ9��L�6�c���[sh���[�#�!�̡��%�\H�G<W����9���<���-�l�`*�E�wf͌���M[���z�{����{ꮰ��4?���Wp��ze�����j�����{C��e�)T���j޵��ɗ�p��� E*��yn_�� ����/��-�fd�T�}�>ò躿��@vsp	R�&e'��d�n��-�7K[�Ҭ�Ɲ����HU߱������g\~�kd������{ǆ�������1�Uo����;`ձ|*�kk�k���Nk�|kJ2[���QqN�W$ �	HE@��zꮫ�a��n���&���C㲑6��e��Z�t���{��+�YhͲ���WlQ|FՖǪ��8����[��<���E�����6�3�y`@}��uh�3��(�\�{(/Ҁ,ے�!m�׍6XE�lF�/*�Na�j��a�"֌�PA���fJ�<��`x*+��)���g1�
u5�C7SoKk�6��ӭ�T�MGW�3���c3�ܱ�:���myC����P����h��D1(�C��-5;r��5�&5f����lϣ8�_ݾ���'��B5�j�r��SQw��2Z����^�鄑�����W���M�y{`99�c�eБ��2?>B�.́8����@�d�C���9p�G��K�4�֠֬d�/�:c&Dn`~_����2`J�0Q�2:�O�&��Ҽ(V^6'���������K�G���s>r�˷>���R��"/��E奷oyy��?����b�E�O��%8��rӖ�?�b\ҝ��lZztMt���Ǐ#�c1��j3d��p�z!�q�T�@�o��W�Q��[F�[�C5l3�l$f�Fk�>t�\�1#W�ר����x�B1����1x�����0:>?���I���o����a��x�o���;e�~�|���ɏl˗f�ϙ�B�4��	C�|��dHa�}��S��)��'a�1a%�>�ބ�`{6��{\����H#R#{eQ��UV~�ŝ/�܂��y~K�I\FPj��R�>���Zdu/�rý�j�i~J�g{�y��3r�T}�^�[�ɩ\kr���y�ɽ/���42�����k����lB_��{m�	��lS�G2��io�6:F�y�X�S#YQ'Snf�E�H�9��P��Kl�^��(����4U-�)z�"�������%�L�M�uERNNQY�#׸;�RP�y{U�ӂ��A_Wr�O�ys������=�~���'6����e�;�y�1�D^w��������g{�`���u�߇{���-ޛ`�����V��������ۢ�g=}H��������sG�<��N��0.t�漯�J�����1k����s���*N���X�G�~<?�9����q��?z��x��~��|�':����ߌ犞���Z�ǰ�ɏ��791Fړ/�28��`��҂�E�$��易����_�Qw\��=^1�\�閬�V�k	�e�����Y#�=�Y����еt�%c�G��)���Ub�L`K�iP*�]�m�y��	������W<����M{i&R@E�s�Gʥ�O"^�t+t]r�-.�H��m�+�9.�wu�nk#�G�I�h�E��l�=�%�P����"uhk��1e�S����f[�9��\���P!ʽ/"%��|ir�M[�~Z���i��S@(��<�k��f��϶>�+�-���d?���̩!\w�������V�XOQw� ڴI�5����z�_��)�b����B#O�+@�#%R퍬6?3Tw�m*���C9�ޣ�ﳆZ��٘���L&L,N�|��:Ad~�u��=-cP��j���N�����Cx[d��&�����&��[E)T���N?��[��_nX����J���IW��oK��������� _i�`4����x�@��݇?���]��5T#�s#]�g˛��J�\#�?@�+�ome���4�"w�+���?9������ c(*�?�˄x�9���ث�n4K�\�:'g�ʳ��oHT�+J:�"Qs]Q҉��ͷH'>�w%���@���̺w���qH��.���-q��1�l���5�ރ9YDro����b�@[�����'�.�6�	�J��ފb��W��?��܄��v�n�u1E������:=���f�iP�M�Df�C�PnU��v����F>�C�q��Xu�3HU����lӎ���[i�Q7��cU�=�l�Uԙ�~�(+��;����Ҥ���ͪ�rm_�Mͫ�ۻV�߼�Tu�.���2�hW�m�Q�jΗ6�WE�|W�D�Zm�O�C��{�j�ң��@�E������PQtޞ��*9��]:#8fL�29�z
�UM�%r*�����P l;Gmx����;�@Fԋ��p��|�;�6Op���No��6)PിS�G�/��X�A+y��\�s�߻������D�#�^|#�����^�s�L��J���"��~'!!��;�e�i?��ts9${�ȝ%]3����a4P5��`i��y�jÞ9hC#�{��+�Z�Wǿ��c���6`����W6_r4>�ɰt�fF�����WIlc?������g���N������E=UN���Ŭ;��{�B���z�2��!�7Ħ?ڈ�g����kBJ�N���M�����@Ѣo�%:���ԙ�^�]@���%j�:�}X�S��b��8�}�R����\�:|ш��S�n~SL�[8{V�G�/7�;!eJ�#��������>W]��>���;�gZ�q�{D�.�T:�}���9��U��JB�|��z�J��{~B�Y�1h��F]/w9��j�ً��m9]�u�vP;�I�˹��䧇�����\�$��U9F����H]r�j�|��W�y���lZ#?�P�EZ��^>�fL��R�e4�8Un���P�N�_���W����f$���ETe7��yF��To�ҳ�]�#o��ϞLU�r_ԝn�H3���١�����/���i����y_��.ڎ7~�=.N�ϼ9p-�˻�s���7)�e�_��`��2�R����	��w��_rb������>p���)=���Tٻ�*UĶ�#m����p�κ�x�'b�l�$��7��wWح?C�d�T䗧��ס/�6ސ���}�)iC��ᑘ����ߏ�事u; �|ԕ�Z6���EF��)b�".,%�<e�{>Y%{ސ�)���T%w��a䲚��)����Zg�reX��N=V�������^U_ZÏ� �����nH2;Wѩ:�����������ZTz�1�_��Ƕ�������|�?:OT=�ԓ��X����zz2����RoU�������='sҽछτW1�����[ߩ��4��|&�!Ny�V�3X�w�zf�u�IwK�Lo&z#3�����8�U:��sJZ��'ݻ�������do=��V���-�=�/L~ݍ�5��L���F�<�R�%O��KqƩY��5����r�A��S��hk>�:c�����됓��������l|=�5.oFk:�ȷqOL�U��ͷH�.v���?��o�"[v�-��N�J��Jg�Y����Q'����=��ʹ��g�f�_5u{��ꓑ�uF��&�7^_ghVj�"Iu"E!���{�&"ۜD��'�S���'*�IT?ѧ�����'��9�F�OTf�âܝ�'���r���+��(��?�A����n����Ӎ���dw�L�AM%����d+ȯfyy:��z�XM�*��
_�f�T'�s,��@�"<�y�L���K�,8����i��|�3���M���<۾�8r��(FlWVM2d�qg����?�9ؕ��7��+��Ц3۳��6�FƚR�^���ǉ�����Q;ʷ�o)�3�c� W��l�;q߳�(���6�δ�R<�)s��T�;��-�d��T��&�\3�۝v��ȶ��7E=�?h�ݑ�W�Pð:�e1�Tt�������<�j����~�m Lg5�T5���&�e�+]r�}�n*���Ր8:��C�JZ����+ĞR�xh'%&Ś�f���=5�/M���j�Ok�=JNrSmv��"9��^��PD�����ˇuyɡ�������(�޳�l� ��F��z��"j����e)�#�I�����5q��k�[�k��w��3$sPV�z�N�������r39nV�&�5�_�<�P���,]I�y�,���̞��wAooxgH��W^v����i2��t�x����e�p�W�ݬ8���j�_%��e���3ͶC�~��r�-�� 7�]٘,;�ee�~�h8nH4�W_�6����N��K���\u�+�!x�4��V�]�nI��Ƨ�N<VǶ��ڥ�r��;D?�����v������%��J�C)�Ck���zE��Ԙ6>���/���&�T�d���Y�y�g�I�{6E�]�=/��ݨN�	�O2k�m�X��'o�<����U=��ܰ�R���H'7��RW|m��z�rO����\N�i������['[��]J��:�x;ߞ�$_L��e����e��>�/��3��M\~Z#]�X��A�4��h�W�$���*m���i�,z�t�Kd��P�c�#�7�M��R���g,�n��E)���73�Z�J��53e{��cU����Z��U��2O�y1:}�PϮ�V��C6U�i�6�se���1�Ψ�>s�Bջg�Y�i`S�l��sq�=�2�'T�wK_T�R�PC���۷���O����U/Q@�>�9��A$��v���7��\/�;��P�cS)�]���ƚ��}"��c1�7~�O=/*�O�dDܯ"~'�FD����6u� m��^�uV-:j0��)h��A��Q0u���g���o�yd �ݓS#��tӖ�^O�c�=�G�\O}#>�7�ڞ�wl0�8/�O��I�?{����ֵ�Ԑ�ٹ�!o32�aV�_�[��ui�}�^׽���n?R)_���|9ö���+_��r�=D����W���?�`�i�?�ۄ���m��7_{Z���<����G����&߆�k���¹�i��7���kO[_�msW�濧�aO���$s�G���l�{��n9z�����ȶ�����}@l�����0�~�O�h7�7|��8�nQ��B��yZ�5)r��F��d޳�^���2���Σ��i��b�)ONn�yrr�h�a�/E�H䯳K��/U�q��o<��Z����n�7|a���c�׌�H���I����ͳM�I�k��|��! ;��'���i�Q /4�
�b��aQ����+��}x�� ����7�v���u�}���K�K�˒����y�w;tc]-%��)��h�Ml^O�6���	D�M�ؽM��6M`c?h���~�4a����e
y���ÇZSa������\�)�cDu|�u��(�k7: 9��ħ@���v���/\��vYw��ދ�z�}d���Z��7�arrWZ#�n��Ø /֍��g�ϧ�i���<����o��ͩ��N9�#�"��^�uW�m����s�K����m-Z3��[���7��K��vIR�/UI��N{>�>[��T*�-�;�ZB엀�ޢ���W��=J~_S��:��.rQ�<4=tŁ�E?#C�����A%��;�Yj�e�X9�y-a>��*ʔ�іf��OV۟�"Z��4TDt���JD'qJ�R]�,��%r(���<#+���y&���\��'��T� ��<��˖C�s\ߝv[u]G,�ψ��9��w��dW�3\��d9���'��v�V��F/�A[D�懼��Üi�j=�8����ϕ�
����O0�����|�n#^��[޿l'�:5����uHů��VI�����$�8X7�]��3��`;e0O�u�G̷�-�ۚ�ב�7���?jy�'��a7y�v�W���C��6g� �G·��6ߺ�|3
Yo�Omu�/��ɿ����_nچ��!p�)q¶���l�}�)q_�o�QV���/ٕ�忑�U����m	��v����g\�j�l����G,olv3�h�(o�#o����/n>��͌#o���W�&m�o�v�f�M��$|89[v��g�S99s�K��9�B��}a
�a�l
�ob��4����v�����C�͗�1���j�;M}�m}�e�;ꛯ���m������@�}���D������ݮ��ϟ$s�k�~AT���3/�rz�qO�Ҥ�Ui�^��-�[�&l�V�.�>-�����o���	�k�N�n����7������sL}�Џ�'揌\{+�'���Me=����蒑��$z�n�wohF��P���V�G[]h��z����p�蠓�:Y頓�:y�K�Q��f��󄩇~牘���΋m��F�?��F?��S�}r��h*���]\}T��[���'4�c��.c��e��	���eoQ��^{c���~�����T�N��})}�,�$)��M�aNT�G����h�%�c6k��+c�������>�O}��=}���>�.���ї�t飭��,��c��O?��G�����ц�b�Q�_�ɯ��k_Z��A�,�oJ�ox��Nb�}���'��+�ϣ�_�����E���*����+����_�ݿ�'���>4��(Ji��>B�35��G�����烞�|ޣ��/���n&?�zT-�zHh���ʴ�Iܙj0����Ǎ	�M�����f���l�S���(sgb�Pcg��<�#��@(_��د�G;�%���c^�e�|oe��M"���x�ϯmr�g�s<��a�x��x�Q�y�F�x�7�ôg��t�=��7Č�|�V�i�'7�o�z0�u礭?&m��!���I��B�%I�a���_D���������;�������R�}��q�_����!I����<���z��5���/ڇ0 !��'r�z� ��q`�����#��ܰ����?{��V:�����s�<�^���[7"m}z��<�<��+=l ��<"O�s×;���7o�o�����G]�M���	��������֣G�����k�����ߎe�F�#_���=<����q����:s��e��j�Z^kF��o��=\|^���?>��r����J���E�,�]�b���ꚍ�u�#����~��t�{��.|�����3������/��EK���a�_l��/��k��̈�/����kd����/`�\s�˒��E襁;��|�E�/���W�/���;�Ofϧۯ�������|��b��G���C1��C�eL�����wO�D��C��|
<$�i�9��_�_Gn��!�_�o�P�+�i����m��(~������p�C^1[����͇N�݀A�ӭ���Ѳ���C�Aer����0��]��ײ�3R�P|)V�e�&9�S�TUJ�)�~�(��8(���R�[m�sy��n��Yh ����:L��@��	i�R�mf�2�D�l���D������t�/���w����_�����w��s�_�/�վ�#o߻�Y�e�m_����k)�����w�k|�x|'K���l��/ɿ����/��+���9.��@�}���R찘���۾����$�w���q�7�վ�Gܾ�R�����۾�8���������o"m}~���ZEo�Wpv��l���A�[$彺�lϤ��Y�=ߓ�?_m��=S�g�a��n@�?�=��gm�������J)^��Ǘj��Y�?mC�����C؜V��ច��Z���g�~�#[�XK���v�}���,%?�'�}�q��9H�<RJɟ��w`�f�m_����Z����͉۾��}������U�R"I���������+����I7[c��F�����l�e@~�����M���w4[S/o��w�s%��h;ychsZ#��:�9(�f���/��_����������/���j�N鿓H���W�U�jlm�-�{Z���ie�$���CP��n�I�=��W�T�u[�$�M�RyeȎ�s��@����X�E���~����!#�\�o>��9�绉�8C��=^�c/Q9}�	����Z[>�޽ͷ[����d��s�����p]Gݟ�ک�l�N=�1���ww���A�h�}>y�dKc�P):V�^C�	�qv>�yE5�ZRh�uA����֊0�Ob��IU�d�Z9H**0͏�f��C�:CI�����PF�q�R���g-Uw�8*���f�1f�!g�|��V��X��)�j^�⧎�@��^/�����U�����vݩN�o^w����ů;���ԝ�٠ug������M=���F&���m�;��ap�v�-�vZ0v�dl���[�p����}��u�r��ݼ�&N��֊V���F�o��c��1xr����-X--x�h����`�ӂ-��`����k�=F�9H&9-�l��l����`�����;-8���-��ໟڂ�[0=~�K�-�;H
�\=x
��>~ڤw-�k��qZ��[0;�o�<�Z�8�F7������	V�@����e��!=�@z�ʒ�<�Rz���
s򻛭a��.�XK�ҋ�y�����<�����g�ˉ%�ü��M�98�S����*?RP�핅JC�^��b�:-K:*�r���e	��S�S��/��
�벂M��+����g��o�Jr�������V�A-(�/�&�Z(�춂˥�ݬ��O6[��zw=��t �٘Լb�A�BdYq��C곕�.![�?l$~�N<"�XZ�b���T�RQ��~���U�U1�;��]���k�o^�7�$�3���U�W��I_8]��"AW�d����*�l^1j`..�Xh��F�����^�.&^�����#6j�=�0S�K8;r<�R�*G���fDu'�t5T�2yrTV�|��a�]�K$}���+)�ae�;T};k�t��c]4�O>o�V�4�LT��h��Gq��l�_i�L�]�|���<����?|1@�T�p4G)kZ���ej�fʔL��"�2m�f�!��?12}�(ӎh&�Dn�H���ҌP��]�:��r9HXuM�JPӮh��5�+F�-T��α;��!1�>/Q���������D�������aB]6xú�96��]!�NTG$�cI��c��u���vl7$��/��]��������+oL+�q ��Ю㷃�q0����:�%��?��r<�т�>x�:G`�����B��{�k��*�?�_Mؔd�P�H��"Mܮ"�_fy���z�U��=E���4�v��\!����|��5��3�M��y`�|6���|"��Kp�|��"�Ӎ�w��|�n���k$��c'x�GI�J#���oɧ;Fp��+$8��a����_N���J�J#x�7
��o1�\�3����	���	��/��`�ap���/1x��2�c�??7������?���?^��������~0�'���<S���g���Tx�VCC��!���3�2��鑷�Y�ğ��BQ&R���zAc8���;d;4DqC��ʥ�VA�uۛW���r+y"O��/ް\��UG�3���4i��7��mեZި�5>ZxX4���KaB�b:��c��,�һ���{��y���z�?���?����.&:����_���]v�N�����P�h��ȖF�G�"e݀��=��Z�֧�;bO�y�众"�{�
������u�Mq�׫�<���y���-R�{+m~����D���gFfI�*}sp�!}�w����|~�ɉ�5�t�J=1R�%g�7�ķ�����c��_P\�?�SN�2R�T����?���a�ߔ-��D��V������om��{�����ƒϲ};�$u�S{SB[E욃�(�j7q�!_����Q#�����Z������Tf*X�����<�xu[�n�>��^�����C�p���h�Y�QCs�~q�7����g���}�����%���5�oȷ��Ƽ:O͇�g�mW�ĥ����+l�ͷ&������E��]9�WV�K�%�v~�ާ����$ɞ�m+W*�4�����C���^�����J��7��Pm�������>ǘi2��`s"I?����$Ku�W�5���$�"E됖#��E��_�AU#eȹ�v�R�!=u�c�w�Z�x�i�]���w���]^+�y�;nXs�~���y�n~����"7\��ⴕ��1I�x��m$K����uLZ�
���_k�g;�~Z�>��D$#;��®�Ɔ��oy��wJ^y)��Lپ4��w�T�DWp<_�qh�ۯ��& ��I�?���Y�#'_��׷x=�;���c�����n���wg��8���ìs�}�<��;g���t�?/�W�x�0w'�\��7�o��h�ћ�zV�p�~!���g��k�?�)�������7>h�w,G�gc��	Y��K�����O�}�-f�wd�_i/����0�[�n_��iFz���N���_����s������n{ƌ:�3s��3�i���oW��Go��2�ĥxJ4�:�=�!Ino�b"U)"��Ʌ��O�F�;F oQW�o��^Bd�,y�ݬ�M~1���C��Op/�|�5��|�|�Z�I��)%_r߽\�*��Ԫ��f��$+8	�ѫ�R.*u��n�5�dݩw�tYF3D���
X~�A/��E����u�֍�C>(��b��韪��B�;{����\�>��h�g��?�M~���D����fF>(d�����r
�;��;��d���7�8�;���q?�]|D�]~���.uv#�.�k'�rCq�~����H����sq�*�N�1G��,�<�i��j�;�����d���W�u�����,6v=ɢJt���ʲm��L����@\>�����m~g��U�+�&�>*��f�䓬������|������Ca����ߐX�x�a�xHAx�2�|��A�I�G���J4�.�Z6R��da���TѐVR�p��]�.\r�0���֌�����;����[Ի�;����I��5��uy��R���W����Q#y-��1�K����J��!q����`���7�����7.r�~jCp���q���Q���ȟ��}�e�|�GZ6�W�-kI߲q�b�S����3eJ��l�H����gh���yX�7�Ok������UR(���]�U��g+�/Zrف��3���2���J��~ßQ�S����
�m�_���?�������k���M�&��h���{Uk΁��L��ظJ+�|�n���<�t�����D��B�G��@���R1"4%%����6����������$[���2�91:Z���;��|�_�*V�du\+Z��Vg��OEv5sQ���������z�h�)ly'�ZRjdr.��D��.���;>���;��N�d�nV[��Д�~��d�nl&(c�}^���W�t��!J���nkZF(�Qk(�mۭ�s޲�����W���m�|��Ik8HPS2���p�d��%=/#�)��)=O�����qO;���
MIUe�b._\�w��E�))=Q���d~�_$��6�?}
��7���~�����:�������^c~�\�݋�����z ̗�Gq+�̗�z�`���{��)�=��+�]�|���j�%���,?h�c����䳿5��m7��D0~����(ڪ��o���Wk���Wr���Wv����	��|���/߂0��_�5�+?���W֏������A�v(U6/�.�(G?��_�D^���[�P��l�F�&�z�%�Z׋��jN���:�0kFvԉ�l:��i���ۨ�T�8��iI]P�+�>�2΀�s`�z�%�������G[���}qM�nԱ]qc7�+ve��T��u�q�ܡcwč�ұ�qc�u�vWl}��uB�o[�����} ��wǍ����㖼]��T�6u�|uL���(p�+�*.b��E������6��A���O�b�������V��)����U+X��|i�dM�Wn��;4!��l�fn�I'�`���4a�֦	��1�J����6����Ҍ�ce���ڴ	2J�}�y�Q����&egY�u@�4��_ ���,�Ց��^��	��DCs���=(?���A3�< 
g^�y>>J[�Q���L�t:#h���ת�4���y���ͺ�?�lŜ'����ў������J�ugk���h�<+�[��g�Ęs�/b}��5�������mZ	�6޳�c���/`\�r�]�i+(ݡ��V�}:٠�L0>S?�r�jy��1��i�n4�&a�|��0�*jM����R�סFO��ѠT�:����巵���}ݣ��K�}�V����q�n�,Yۆ�ܳZf��NE�_ݬ�����X�:6�:e�бq�)�C��]/,YM�\�T�v��=�z�[-31녵Rg�g��,��nc����I,D���IDA�Qd|�z���R:��t+�*�}_���,
��#������׏���+�9�3�<ζ��#�����;b[���\QQo�F�S���
,�u��[Cu�-˼�]~���7v��:�oK.B�7�Ũ)�ǥ����o���7���j����̶�����3���)��ro���-q��mS�dY�ַj}ۮ'���I��t�h�������̒|̒�c��_�v��!j���Զ;#�<&GP�I���!u<�0�.ql�ܘ 6(��ۭ`{�b�VpG�Xk�g!L�\��vXAN0�Z��-:�&+(s,~�+�w`�2�o�=n�Ǿg�%�}�
H�>�vYA����vZ���E��|��׃�9Wl���+�=�)�Ey|N�ʰ���]����{������i�gIQ+�4�H,D����w������τQ�	5*� AA!$0�a�L&B��<0����!�qDS���mJiK[ۦ^E�T�C�\�b��H��BmT�h���������d&/�������f�?����k���>k�^�Tr�1srܮ��c�r��m͘���[�nY�0穸�˪�	���_�UۮV�0�'Bp儂�9?�4���r3m��e7o�l��0�M�瘊�里؎��c�}	q���[�˥Z*��������@ ���XC�둎R5TGf2�F�Y�B�>ჩj]��#��H�����M�<[�!�\kȳ�	-G֧�,w�x�^@�C��,��K�6ܽ^J�N�K�n#�r�ޠ�R._���)yx�Բ��$1�῭/��s�"y8��,wR���(!�����$��	ヱG�t{d��G�E�;��Gct��#�=�G��H��G�J{��0��g�E�G楃��FԹ�#�m����#jI�f:�T	o�覊����r<�1"c�T�������p�1���n�$��HK�%�&���p�A3����&}Q��'�"�n��_r�a�ۍY����J%ɲ(�d�ͺ����y����s��w�����#���<���#�t��D���)�/����j�" ��Lu՜]R&��K�.�H,����W֙łq?�Gs���G=7��\��U����cC&6�C��W�8�,_��Ug���*��V���p?�3$`>oP;���uW�G>���w���O����@������y=M
q����Z��u��:����ܭ@=Q������?wG���k1������X}���[���_o��V�9�wG}���*]��G��h���].�����}am��~�2����s��3.S�T_L���#���5��<���=f�G��G������3/�z�J�s�]Z��R���TE������T������]���@�����i���X��Yڏ\�] ��MtWsK	�]'�r(:��PIw�oYf �t��{F,|�ɓ���*��)�t�T���׎q�4=���S?�/���"=|��q��&z����s���҃N ���ɻ�M��j���ⳳ�����U�p�8�8�_�(���3"�uq/�|��/jt'z�Ӿ�c}�~�2���]���J����Ӳ�=��/���H1q�T%,DШ�r�XO���M��?ڡ�瑻���j��R�׀�K��.�_�R��9Q��b���������#P���D*׸';�6���?�bG�_�N��qA�ׅ���D���#B%���[_W������O~�JW��$N`=�Z��q�gʅ0�{ϡ����߮�k�����9S�?��>��hB�{�	5�C�J�h
a�J����u&��X�����|���T�V+Xc���	���<�r��!�m�/�ׄ�o�by�ik�81;����/�8P��&���νO��M,���=�둎ދ�i����8���s�*�8��R:�v��X�xYʱ�ކ���	ʏ���+?�͛��hiƯZ��:M�����]������{�@,�|�J6dek�����-�k���W���S�����q��|;�ݘ��Oӑ�t ��84p��k��OLǷ���=-�OH1�<��K��V�1#ޛo�N�W&�n�n�J���ۥ��h�4�/��M?��'��&�)O]I�M?�F�0�Nn���<4��@b��Ȼ����5ɻd:`�u>�GI[�%V�%g��}W@nI�)+��G���	�d�������f��2����j����AW���:+��Ƅ���ס�&(3c��G��c��HZ�ן}���WW�A����M'z��2,=S=�@^b}�'w?��1B��'\�J�Q�ݞ�1�m����aG(ݖJ|V�F�G���}u'�t�A�����Z�H�c�W>
:���1�ID�gD r}�Z�mT��~��������Xצ(�)�l>h!��r{�v]J�㤗��Q�_K��h����#Z���c�@��/��'��tк�gt]��^r������o5���Iy/��OB��A��0�6޾MD��g�? ϫ��U���A������؏T����������T��Ua�{����!��m\ˏ��-�Ƒw[mS�I�M���;��ߔ�ަ����NL���~T_2.0*Pp@'٦���}+b����D�^��vY@ɸ]���3�UC4Z��B�=-Z��w�i�{nB�n+�����G���2"�E�FB{�O�7饉�]�J�0r_Ue���aH�%����9ݖ�^oY`䦒nQ�~lP�%�m����ˌ������y�� �Fy��K�!��xI>I� �~ZZJN9��A�/�Sg�ƚ_�'���`�_O�3�l���s(��0�~x��$��Vq9�}�@��s(���~W���l���âU��C�q���s��}��w�Mt��s���W?$$r������S��C�d"�V�<?@�]ʫ�B��sq--a�x^&����)!Ҟ�T�E:b7�Jek_�0�_�#n�b��aq��w��j�ס4�v��@����%;� _��H}(�LEw*@*#U<,S�E����9 v@hJ:�0��� q�����/�9 ����#/$e��Mb`觸�H��a��Ir��ϊ?֕�+�v���9
�O�yI�yA^�q�=���+�}�zb�'K�`՛��H�b��>�&�"Y`O<ײ�TYt�怿�)Է���J���=�������y�_�.��NRb;�W�����������:�)P�a�[���G1���}�:�<3��-��h|J,n�ȸ]q��@c�q	��`@�Yq+�
4�N���$_�����O�ν�a��I>l�c�o���[�QJ�c�{�~�a��Lv�8���n���:����=��.r��(��*.��7n�{�"�7�Cϲg|�o2��7[��n�ܢ�p�x^h�M��7�e�'���$�4Q�(B%[�<��y��ʋsӷ=_������7��Y����u����P���p�����H�����oE�.4�I�-f}{�����?��o�:��{�9���}���Mt;�����շ��s�Y����a��=+"��V���ʁ�c�p�11��	-t���[7�A���19q�.�۵��|(J_}U�s��3Z����Z��_���_˯��G��o��/�r���-7���mв<�������W�m�_�}_^n��@���~��֖��U�߃���{��x�iҊK�㣴�J`4\$ߩR�/�>t�f��ko�WVD�J�[��~�Ը_��{��Ko!zP]�XB;��9�P���yC��,�4Q�e�J02�|���k���_�|��|�	�����W���}��œc�;���a���
��ϲ���e��l%g�v�����q�ϖ�eɊ��r�za���+��}����s���^�_N������mz�qd�牯-7��-�E!뿢�~���V��FtU�so������D��߆"�ȸ�{�ԱO���;���3���%�qo]��y�@��c(�9�P>K��������s����9W=������~��趲�������g�A��B3��(�~WA?�������_���f�oK��ǒAΟC�?����E&>(\���h�@���P�O��i���罢�ϟ/
�ϟ�.#zV.>����g��-5�-���튂�ΟD�D������Ú?o�G�oO^"���i���O�7޿v�6{0���%ܾ}�fn�n������־]�پ�ZѾ�0���כa�X[�(���ٷGu���`�[�>9 ���ٷw/���m�os��}[��۷7.2۷]��ڷ'�>�~rx�=:�}�#쿼�۷o��Z����`�Yh�%k�پݰ0�}��hq�e���ۏn6ٷB�/��}w�����۾ݱ�l�>/�?-�~�3�</�~~w�i��s9=��H?��~�g(�m�f��{�������#��y0���>��gy&�5�p�ݓ3\�<� �/��kK?���?�o����ߛÓTA�}�H�����y}(�8�������6�n�@����̟b�9V���g���ϟ+l��ϤX��l�8R�̟�\�Ҳ8��dw��$��e�?����23�}}!ȑ5��4��Eb�}	�2���<M� �Ӽ����ep{���v��ٌ���f{w^ND{w��D�f�k�;�ٻ/��4�Vz}]��#E��'i�������g�+���q��%��1x��1c�Gj����s�&0�8T���"�]絷�s���؈��$7|�С�>�PAǰ����Ke_C�����U͊گ�<͙�O?��~�g�c����i����P��ʰ������!���Ǉ�V����}�?2�a�c^����b�c�9ꇴ�����y!�����Ǽ>�����y�#Z���y���?;O�r��i������+������s;Osќ��i�K7���rӀ�iha��r�f�d���4OƵZ��i���Ѵ�!����0�o�)�������6���������d߆@#�US�2Ḃ��۳�Aa�fD��0N�3��v���N�������Q��9��;G�6�s4��.z�����֨���k�X�9M�9�'#���|.��65����n��W	l3�����NY�����&�~I"�W�#��z�fW�?�M�����������_��������4��M�E���c�{Y�)���3�u����wh��ߪ�ovHb��ᒘ��E��f�ᖜDn�*��6�~~)�`J���O~Ao�v~��D��?=���	:'^j��I�����#d�x��C�1/�a����qt��"�?fY��O}�N]���
�(jFs�͗�QPK����ͤ��ug�r~:��Ϗ����~�J�|`���͇�2�6ݸ��-eʚ����-�&�8�{�<�RxFӋĻ^k�	�HY��█��vΓ�N���(��D�V��o�<�B�Z%j�'�e{e+��Kq�T�w�}������O����vj���|H^��hi\�>N��}�������9��B���?��yϛ��nj>�u���}�±�DE�s"�
I�lɖ3�2�O�C	�c��M�r(�Q���3�������W;_�w��>�D2��)�:���eH�b����^y�G����<X��>:�Pwzw�%�Sa�Y)��kgɛ������ޯz�����G���Ī��i<�F�����M�-����=��E%G��V>�EX�1��h�H�Ľ�G	Wp�5�e
��7��H��n�������G���NP��G^�{�����_0~̑H��u����٘#�_��������Y��#&�L����������\��>7�G�Rb+�[����GwDǿu���<@{������.�2�(�Hx��}�K��yħ�1@|� ��� �p����W�����x�-6E�	�	��Ɉ�n���ޛ���������@&�wt˱M�ǷM�n�ɞ��aA���QyA9'���?�O|L��;��P�j����6����'4�����m����C̗���o��R���:�O���T��W�c�|���%�
IW��r�ّގCY��&��h>;�;��l��;��I�>�@�D:�8m�=&|F�0����p���wzY���e��M%���l���󔳂�}�&ư5�9#�"�\~�(��˟4��7��v'���O��1�`�!��������(����|f9e$�����͈M9=�LU����~۳Q����3��,���=��=gc�<K���rf�����-�ａ�olsG�,%V_i2��p�����>�������o�ȵ4R}WG�O��GG�����|�]!����(�;R�GʿP�_)���w_,r^v}�~����oQj�Kz6�S�3A�RS��):���+�{�ؤ�;E򣘱ĉgB9�����B���P�ZQ@� \,���o�3��^r������	� �O�õ_H�ψ2~7Y�0A7��D��È�;C�a1u�y��6�.��R�����Ni������F��A�����Of�Q��_7��4}���%��i0�'i���X��}� ʿ8��D��S�5C-_��XQ�U���/N���>#V4�b���E�wN�O,}�?��Ţ<j�~%�"�r�]3co��P�Y�m���x���nWZ�剺�B� o���#Q�wD���������V~�ԡ��.�?_��?��/r�o�����ľ埙"�?���a���?��-��3��������jQ�u�}a�AW�!��b}z(C�B��6��tkgA|�޸�w�����Ɏޒ��x��TK�|0���h�ȿ���	&w`yt����b����I��M,���c��֫M�;o[�P��,�զ�������H�O��Tk4�d<����4/~�Mk���T|i��l�����7)n�ec�}t��G,I����x�k���+�{{O],�'������!�s�J��#��z�hۊ��xҞ��"����b\����>�l�k���}+΃\j%��)?�r~Y,7�I���{B0�l��/G��N���?^K;�)��G
�t`�8��Qp�k^b�bp0v��M-���O��&�&\k`9]�#���;�E�87 .��������ύoj���[
QT\�!jNḖcq����t�k���#6Q*�fܣৗ��S)���g/�.�F�[���V���w�����@.��l�;��H?�>/�95��J�4KR_��$��YO�.�8<Ȝ'#�ˣS�}vw�?7��w �8@䣇��</^�ύ��^��U]���9��W�D:tA���B�w���GU�����M*��������a�Ю�EB���� WZع�lE�@.=���z���jRo?yPGb?wD +����ͧcS:�c��61&P�8V�s�r�76���W��| V��D����G�x� �)MK��osW�z��?��nt 6��H�ss�x�DY�z*�_�)��;C��5W�W����r����3��M��x�sz�.,�?!�S�0���F�E�o>-z�^QLJ`]t��D�{�z����1j��HZ�FT�ha�~�����ϊ�\īi=�%+��E�͟[�����c��Z���C׏}�ל�O��:��[cc6B|l��eݯ&��>��v��v@(�������D�C�����[V���Bһ�I?G��ӕ<�7�I�H�Ӑ�q�����ӵ!��9��E�!�]����㲐��~�/�߿��ib��R<��ʰ�ʃ|�ȍwq���
�H�CV&�:Ο9�i��{Y�9��P�x��)�ج��]E��/*��q���ך��!në}ɭl�
<�SzS>�/��+��ɧx��j�"e���vly|�Z�����z<��%����5}Q᭾q����[��%��S�="����=�w'PK[aϜjFz� ½ͽ��?��謁���E��)_�}�S��}O�/�xa�80�>H�z{�=������oY���'�L���_x�Zv��ǳ��CʍېI͔e �N��*{���������O�+j�J���AY�h^��rO:�n����릍�{D���C�t��	��*��b|�=$����WϞ
WkEK7�,��w��Z�h>��[?�hiaoa���-�J�Q��tSIW�N���{��
o¼J��y��Q��٢��E��߈��VT�{О� v�3�e����m����s��?t����x��&�'�"p�(����5DO���^�(�[|J�$Qe+������e!���kB��<o�$�~z�����&k��{�����:_}��	;�l��8ǅ�b����}t�m` ���������#�M�OR��Qdw}���z����w!BB������N�vZ�
6"��u\%?)����;>���*�?��d�B��m�.G|�x�ٍP骭u�����.p8��E�kJ	���߅�:��݉?	u!�#�!GЮ��w�
�m�nC����g!>߼�NCZV",L��7�a�T4J������3����6 M��נ��M�~ۍС�ކ�S�/Ri�T���.��U��	��M�ގС⧩�J��{QBB!�\�P�ЄЪ~oChW�W�P�B�{2t��o�q+#���'����_����6�;���0��uFH������4�a��W�9]��2ha��!��O���x��a��W�9]�{]����uY�1���V��j�[k�o���a�����:��^�R&U��-�j��5��
*���z��:���Ua�w�8��������q{}��VoiY�̜i��p������Z��2��Ya][�F�*��t�lIe��J�U�:��kuUZ����Zb�k$�d:������%������R�'خ��ڮG�'�^Ԅ��:�i��ƹ�U^�AM�媇f
��8M��Ȧ�7�bxZ�c�����}�^��Q�vx�_��e���u�5��>���t	�A�ӂĸՁ��T��)��W_�r{Q�:T(��9QVM�*QP-�3jZ���b��MVU����W[�}n7�â� ��QZ!
���rWM/C�����kK�V����Fk�ז:���h0�N!k[���o+�P�qn��q�VX'P�e5U�R���@/C@D�sV��И�( g8>Qy=���\��K�"f���)#z;�z%��^�w��*�?n�T�M�����]Z�YN�U�TB��n���?d�U��kK��
�NC�_M�<g��a�y�i�/���8�C��jf����2��/�������ZWĪ��7����[���<�\g�g	���	"������)����-v8*<��_&��2Ե֓_���ݮH,ڟ,Sb��r��`���T�!^�$�o�'O�ykj�/Z�W�O�pC$Cߠ̹����@��7ʆ�pU8�;�4`숚ʚ��$�Y��DS�Sv4�.eG�Rn��$�kK���u�g��r���ͱ�4�;�:\[�pZ�A릲�V)`�Jm�n��4#�A�2��6�&�'ҫD�<�̉V�+j]�h��O6��UZA-���ɋ���X$}\�.uV�6*]����� ������7��<��祺��)]J�ƁZX�A�R櫒�뗭��L��>��ҞS]�v��^S޺-'�n��\�����֜�\f΀�HF�n�-*e�-v��Oi��:�xI��)��AE>�l�#8���>f���J�f�P���I*א�M��B���^+-/GQ�Ѳb���m��Z=���U�.-����$��a$l�>�C�G�{�f�>�]w��y���G1�^��y+F}\R	��H"�\��T,6%��D�|kJ$~��ڕ�T9�hF��N�VL��VIx�`ɡ?�$˪��(v��o��e!�"x��u^"v�V�/*G�A	B2�\��R'�ܪ���*ۭ!�d�i���R�=�i�@*��g��Ys1�g�Z%}S�ry>����v�$sek�ʕ�s�D|��aX��q��>�3�%Tp�������Hs����L��:M6	s�擆�5#.��k}?��V��#&��qFV<W��d4c�����U��z4�cm�Z����6�X
�g��Z��QY��u�b�׺��X�Ӄ���"��� �-d�B�ժ��-B^��;�ja4d�rEc�XPhl}�����*��g-�����my���Lֵf��5n�j}�Y���Z{Sc�&-B�x�n�i���Ǡ�L&���ф�v^�t��u?^[�Y�x�u�bkvfъ��f�C3i�PJ-�Q:M!���}NC���L�9�r��:��TLќ.'�a���;X�cw�VB]�������֛��ac냱��գ���?���y�g��t��A����F؇p�J�1>�`��A��0!��B^{a3�v���!C8��1B��h�|��0!�gjp��A����F؇p���QkP��YEen�6#l_#�zZ}���1��>?F�Z��& �@�B(B(Cp#<��a;����!�@�!��d��9���W�!�!�D�����v��4�>�c'X���=j�A��0!����� �f��O#�[�������q�_��	��c��{@;�	3����"lF؎�4�>�c'>F���& �@�B(B(Cp�+�z���+�4>��۷M��o'��1B�}(a��,�����e��Fxa�}}����4�>�c'>F�jDf d!!�!�D،��i�}�aڭ~;�Ϗ��q�܎��2�,ZG�E|�٢5!d t,�o���g2B��ֶ��'�_*�K��j	>�����8���U>�*��oB~+����r�|�/2�_�?����N����-!�a�	7������/��GbN�:y��=m�q��<�#�gC���	Cm�7t|��Oұ8��%ަ�Q�3;��+mǝ:>_|�:t,�:�7�t|����ѱ8��ů��E�iQ�b�Ĳ��8^|�)��h�ym��ǈ���eG;�Q
�SZ�:_"�ė�ό �L��ⰍVė��UA|���}:�R���4�7B�ʄ�6�kLت�n��YP^9p���������D]�5��-��"V��X�j�12�tS�͠��Y��c}�k}-�o�f��z�ɤ�Z󈢏E��ܕeG+�3|����r�B�'�������f���8��~˔��ǖ���:���F�g�����
����,�s����W��FYB1՗���,gx�)��&L�!��x]-�/�7�O�y�T�/L�;�p��n�k�H[�����'0L��0���qWw0LG�v�	5�=��n �`������+Y����?��	��o5��~�]�B�ۀ��?��2�s��,����?C�}���S��H�3L�>L�3�*���ǈ���?�f�{3�q~ ~�����d���)������u�w��i����b��;��,ƛa�z�i�w2L������g����]I�f��T��H�m?���{!⏳�x`��|	�S?0���|�F��W1<x2�I�	?2�L�n�����������J'��~���2������It3|���[��������:J����&~�1ɫh����b�����p=�Of�*?�Ng����up�'7Kn�`�	`/�ߣ�3��A�w?���0� �k�_ >�0���:��?`�n���ǀ{&On1.�|��(,��g1L7�1�)їa��T�pL�5�U8-_L�l1L/ >���?e���x��k��0]4�
�3��e�����ᛀ?g���7�"�q�M�S^�����s&�O�W�2�v0����{�b�	�I���Ï ���f�?1�������Z"�m���d�����.��c��Nc���m�[��,����_���?�0L>/�~�;�;�;�����{�
���04{� ���?�ϲ�K�-n��cx�$�'Oe8	xé����az��\�5l~ө�:_��a:P���;��p�O^��a:�|��5��0�|�����p �Û��d�;��{�F������X����0�,�\�� /`x?�b�_���׀�>M{�~����{�[�;p��O�7�6�4�[��a8�p���[���ᫀ�1��Um����\�p:�����U^ ���Ŕ�a�8���픿��e�O1\\ϰ8�a/�YF�{��0�����!�?
|��s+�i��<�.��v��V�o�ϰ��T�/o`� pB��_�++�u�l�?�����x���p���πkYy_oa�<�N?� ٫�M�^��e��_�����O�gx:pó��`x.p�?�	�������^���-�^�����>���3|7��a�1����{�L�g�O�g�1`+�[�������������/������������H-�G��+&�W����/������7����~�������S�U�?*4����J;s�����p�\��Tềio\�[�i_v�¿����
�L��z�������J���iK3Ϣ�*<%F�OTx0�/T�A�o�hs����Sx3p�;c�>���Eʟo�d�O�b8�|M���8���u��|����{���L�t|���S�e���q��:�yA�x�?S��'և��2�5a���3��h��`�'��T�Äi]��	`�O�A�?p��p!�/P��
��=x}���~�t��0���o5��p�m����w2L[�i�<�aگ��0�W�1,T������,��5�KN�^<���1'_����z��/0�_���x�nS��jꩃ�����e�Y�G���f��]?<�������᷁G1�7jß�������������������N���&���>1M� g�Kk��i�F�;��sF�.!qp�V��?���4���c�b��Y4z=�����|��������K�E�]/�gJ��&��j�}4F6 |r�l<�l}_ӮR��n߃9����4�\}�h�w�5Ӣݬ���O�E<9!��b�>ćN��M{@�?�u�%���'�kn}Ǡ������Y{�	\��8����m7Y�I��k	���+<8��xnA�vzd��Sv�ڌ��<�շ��W��Q\h�����*�E��ڢ}S���^��*�Jd���?�	����L�UG�&W�f���.�z�৻)~��?m��3���a=JR����Ѵ{ϓ�]�N�E�P����?^�R���kopg�E<���3��/�#��[�>8�l����ēO�N��a��g�=2�x~F�}���(m��Wh;G�ҿ��_����-Z���3��xrHx��|�Q�
��[M�S�o�nSP���~�is�W�C�͇j��VM{A�x#��f����c<o��j�Q�#yp��oӴ�T���a�����/)=��Q0���x�@��)����\�vM�^շ�����lDT������ ����&��ǋ������_��a4d*|�Uk?�8^ysTŧ �`����h�~%p�/�W���t�	��A1�E|3p˿��3�3S�������[Y����6�=�����c��6�t?��*<�)��t�V~��o'(��������� �Zi���;����?��ִo)�����x�Mx/�G{�T����l>���M���9
ik�4��xM�O�a�6�gx���yU�}����H��6���4����_��M/�}��� �ϱ��:���e����s�!�3����^	���t�'/2�����������y����g��O���y2M��s�E�ʻ�[�U���x'k��	����s�!?VgtiZ��_I�Y������Ǘz(��T�'��z���M�_R���V-���Y�>nc�y���3Y�)���yJ����g������>��one�IG<�ĺ���C��5��}�߬i[?�n�΢ݦ�O_N�W��X�1�k1�� ��o胋1��-���+�{ L�TxML��
�q�Q��^�L^o��z��.O�>�B&��GY~�׀����sO��8~��~&r2꟪ʛ���O>����vgt��6*´\�6������s���~x+�ǟ�3{p$-F�l�}�l�h�W	�d֞�6���*����6��n�ǰnc��	�d؛��=�z]Ď��x�ΰ�����W�h�/����S� p�#�8W#���i��~����/ѰO?N��&���fG�h�/�:��q�W����;����y���ˁ�}��mԿ���#��z#�5��l|ߧ�������w�5���w�7����������Cf��Y�VV^!p�s��_�>°_��K,Z��;�	-����1*~p�|�_NR�l|0h]��9�}
����m��VC4 g��i!&��(�7��PF�
�n�݈�0���ߦ�`O���p�#����j�?);b<�w�E�P|���g�����0_}o^���nc�*�Тݮ�8��1_ܹ��ߌ�7�{�P�>���'�SY}#&h�Q?����d�v�7TyӁ��7�m�P/ v3~.�����	ti�E�D�cpr�%8 .d�{�����E����#^{E�w_�C�ޡ� T�c~,~�����iM���7��}�]�XV�/����xh�<�)��W��M{L�?����}_�Q�����8�0�O���<�:��R�>��	�2��^�X{n{�X/~������W0�1&���S��^�&A�1<��y�~�	�c5�Bஇ}�nz�H�	8��^���q�E{Y��n����o����������/��.������V�o�,ڥ��i�_����p�O4��n[j̷��ٌ�?�f�����/��m����߈��Ga�:MKd�]�v���r5p'��x���a��w���R�U\~7���Ne��o��~�)p�� �e�;�<�s��^�.�_��:��/�wNPz�נ}N��7�����K��՟	���/n�g����;��( \��a�<���\j̯?���D��+��x��oִ�*���|����[F�h=�i���~���&�6����iY��Z`�7��8���$p�Lc��0�ˍ��P�^c>łq����j������7�U�<�&����Ni��
� '_f�&(��;�]���tz�Þ}Cᷩ��u��&��)c���Nc���_�ݨ��o�Z`+����o�����W^�+���������T��A�ذ��@�C~/R�����_q��o2��p2+/�6���z?�:��r�&f��H02�kk���g=�����V��O�F�)�����N�e��BL�=���
�|����3���XI�_��p'��ng��m�|@��W�A��T�� ~�+��IB�)?M�����<)�v����`�y��p�#l~�������3��.���,��ͪ�{5:-�V���n�f(��-֐w� �2zm�x���4!�O!����շĘ_�'c=��On2���O��L��W�P����i���������[��}���s3��3�s/p'�����}y
����h�<V�E�Xo�R�]le�=�m���PFx�|~Nxp=��)�p�a��OP<�?�a�|D���*%���P�l?�e��oa\T�ZmM�xk:�����ޚ$������4�\�v�*J��I�Rx��Jz��n�/)���-+�ہ�CP�B{nQfA�=+gA�b��"��p٫j]e���
�����rW]}���H��:Q������L��]Z�W����i.��?~�1S3�AÒ�m��O�f���y�3��I�fj��s�&�WB@��b�����^�v{Rjʬ�(x&U@5�!!!�����jM
�M��)�z%�A�fR���n&��I�fR���*r&%�I�S)q*%�A��#u��7�檫s9	f����J�BE�P3����}#�	�( U#5�FjÍ�WT��T��T@�H�i�#�r�Q�4ʑ6[[�8O�e�Qfe�����#�"��$(c�����l��6�p�h�M4�&�n���yg��3D��A� �MP�&�lt�	B��m3%�����6Ar���M�&�nd�	��RE�T�7U�ț*򦊼�"�,�W��m�dK�w��;K��d�%��yg���E��"�l�w��;[�-��yg���E��"�W�X�Y�Z�[�\ۍr�D^1�61�61�61�61�61��4�>M�L)�E�tQr�H�.Ҥ�2�Ո�!O���,�;Y�q��d�R�����'#HH�ß"G>Ez��9�i�����d�/R$��H�I��jUm�I*�T\�,+H��%�ʓ%$��\�q���ei3ë���3U�,Tr_�d��s)�S$7�HLIU�F���2��$7�HvL���"X1U�z���d��>b�f����.�Ob�SE{R��BHT�*%�hJ�hI�hA�h@��?Ut)U0|�`�T���/����Sç
�O��)���d)*]+���J�'��FT�p��O~���w4|V�s�{i}C��*��\}���N��|�7������R��E�����x{��7`�:Oh�4�T="�+����D}&�M�ƨF�!"����S-/��>�o�p��g����Wr��O�V��9�f��Ho^�����Yfn�*s��t0'
�rs�p�4!3�^V�q��]Ʈ���rˉE�p�o�-��*���Z���0��@�^�~����H$�
~ee6�J% 2H�̐bFH�$K�1�m��>�]vO�=�L�J�.|*I`+^i�R:�^:�sK@Y��=�Y�^N.�|�����&�4d�6Y}u;��Jp8u�L�lLH�bI�ݓ}���"�.��V������"��	��ZW�}m�a��,���4�uD���ݰ��K��ub!!��K�`z��.ɦٗg۵,W�twWQ�I-X����	ƣ���YA?�l�l��KW��B���)5����vT�KH�,���]�^.��QW^�N�������Gl�tҖ�\���Wa��%�`�	WNުXk4e��3��s�`H`��;Y p��VU\�ٱN��?4S���Ų�ˉ�"�wb�e��֡����[�b��S�p>��!��[a�Q�r+uʳX���WY���(f�t����[.�0�7|ҷZ.�5;��繊�\�FR<����t�K���:�ѥG�s�x��g��hl8�g�$�����u�Z_��BfI���hO)����ٯ���V�
�0B*�^��L*z�����o�o���P��aZ�v@Nzʅc(�B��h�� e܄v�
1'�³�خ�
:LN8e����#=WK>��"t�& q�l}pbɑV�
֯���p����:�Y�!}��\m/�Th�e_y��u��P���`��b�o	�����J��c�٠H/�l��*S��3Tꃋ��c@{a�[NvIQ�=?o�͙r�řY�9�Hbصơ����IU��mT�c��Le.��(6 ��Pj����+�+F"9���u��@���~ۗ�ʴ*��22�	N%g���L��VI���,�B[�(�k���E�ʰ���ksA��~0��Ҕˬ���@���	�����L��<5U�r@C���3z���<��۱h�rG-��ciP�K�"I,{����[���/��̷/��]�S�3X��L7J�ߩ�!ܞV�ϡ��:�b�I]ʬ(�G�ew���u�I .3׮�]!<�R��c�:M�l���]#�(��P�\�$�D2��Ay\a��E��\�*�s��[��ӯ��OC�I���j%=֟
�	2��T�S�J#N'�0
ĸ	��9p�*u۫� 6�쌴�Y�oA�a#�;1�#*02q�3i�J+*"�RyHF��Z�ǡ!�����A�TE�k������	X�&`x1L�d�"r�V*���&'�1/핐a� �]e.w�+��Ϣ@��Z��`�l�sP��t作x6!���Ro5Ԕ�J�ס"��Ɣ��Gw�O�S���^:����1e�F���>}Y�����G')����9�N�*�bu��w��C�U5�ِ��qb��#�U^��܎�b��>@CtZI���J��P,\�cm�B��q��-�~t�#����n�c�b�f^~���ЉH�>�[{F�r�ю �#�y����ᶕ֗��xÒGJtT'aP&2��Y���RS[7uM�b�W`���A����X%�v����-����i��J��]QSI�%l�^w-8��Y�|��H��5�"5��vp�[�p�v��/�djO��z]���X��B������]C�F��6?��u���}F�ʼf���Ќ}Hb�:��H�*�7L	�� ��a�]�V�A�)
�{����r���j�0�Ⳛ*ˍ�����A�Β w�a�r����c�J�d$�j��!����)q=$���Z	G��� �."?ی����k��d���PXz��$��[g�٨�<Q(����$�ٯ��Cc���6���O��b/��ġ�Ү��e�u>'����R7��7I�������u����5r��[G��FTx=#���^p7-����j� 6<�ڝݓ�9!z87x������&��@�xл�rI��Hd\�1��2�a�8Nn��!T7+H*�w,Ț�{kb�V����e/q�MI,˔%f%�D2j��5t�P���y>�D�6IcL���&b���#����.���0�%}�Ψ��U���"��
Z@ʸV�H�5��m���\RB�?[?�	�"5_R�$Mޒ��*E���v�k��¨?ˬ�����KH}���]ª��?�m�>��дS��o`����C/���"�슕�4o���9E���@����Ą@�b�Dd;]�h�}��,	`��潮Ѓ�m/=/�;*�}?U]�b����ժ��b����84mØ&B�D�=!&�`w�ٓV[�Ѥ��d����fY�l��� �^	�
L6�k�^8�[�(�/W���k>�#�5�Cf�|VF�T��bKS_�S�U1�3P��Vd!�>B�CWё��h��Їᦰ��F����O��V�n�%��<=]iW��iL��-$�ΑH���'I\�U��+iQ�6�^�[[����6��el	z�T��R�[�Gxj�%l�,��t�TKJag��@����L['p��f�OA�>�HE�DK����4�V���0���w��E �j�, �[O���h�ԓ�t���!�bw��N�D��3C}�%"?���%w���c���c�>d���o�l��Ji��["�h��'\�w���s������S>���Ϋg=��i0F�(~��<�3;���ʞ��/Cɉ�$�~�_�!��B~�_�%�.�C��j]ؚ����n
j�*�F=���Ɋj�e�\\���� ���k�=�(S�����3��C�?��m�u��%S��I��fh�s��\�^���}y7=����8<�i�'����8��T���9�YI))�R�f̜��iI뜥uX�&9����pkIե�j-iY���Z$�v'�O�[��}3%@���Y- �\�t��6��?��Ib�&�J�{*�3	դ$�� ,�x�y��k����l �cu�[FP�Ʒ$q���T�IBS��eU">�a�q�$O��i�~�cE�=�B�E�tw������@��tt���.�ۏ^�:O����(4]���d:
�N��^��{�(��m�7S��w��5�Uyt_��+d:KG�ӻ���;�cD���?�����J�K�Q�j���'��ث�ѽG�����?R��>$
�#z���F8_�{�(�OP^�٫�ei��$
�Γ�bY�6v��Bg��JI�F���ۡ��;F:�M3Ow�%��9���#�>��s��4�_�1
^�d�>O�t34y_�զ~P�OX:��£̧�E�g�'��L�k)0W;��~��x��j�o�jS�(f�ȿc�:�ƒ�c��ޥy�g�����u�'�H�KG�*-���=���MF��K'�3E�6v'�U}����W�g�h��;�"�P��2�n��H������jD��T9�`1���c�������1ԋ��"�뷕�=a��t&��+��E�f	MG�PK
    +Q�Hk'
��  �� #  org/bridj/lib/sunos_x86/libbridj.so  ��     �      �}@UU�|�RQ\���)����i`�����~�)�����B ��QZ4�ۍ"�g�i�r&���ʌ�
�'*2���Ȩ.aF嘕ʻ��׹g��m������q�g����{���9���:�4�������O|�0FݲKŌ2�hc�q�q�a���Z�&_G129^�EqH��XcC$����_�8Dp�ǹ�{)l����-��?O��~m�M&�8>*�7�c�>:�0�=�0�Ez��FvE�a�@�dPT6��]�k�8�h-e���xt�a��-y�a�E�������_�gM4�G��0������<�Ǩ��zIP��{*�OT�iD/�>0B����<mХ����i�+'�1��h��L��i�т!g��q<]$ZK��v�Œ���`p��f��]g8�$��c�΢+��s�A�O�:_�$M����(�"M��r?F(��+-M*]����M�k]�_!t*]��Jp���L��Z�����ʘMׯ%<ˀ2��ͥ+��<Gx>]�/z]��*��UB��WJW]�ҵ��[��K躍�
���7t�誢�NIs]~�t�C׽Z����ҵ����;����r���?�� ]�ʪ��!��7G���N�?�z�����']��tO���a�AOӵ��g�j��Y����7��]���-t5�����BW]�j�^s��J�tm�k���%�m������ߣk']�����u�PK�)��A��	�k7]�ky��#�K��j�����������:H�!�z���|2�k]G[�9��芣k���@�D��:���$|8��u��D�g�u]It�#����ܟG�|�~NW
]��k]��K���t1]�hac��2�������j��7��[�&���O��+�J�k]�tM��3�~&]���Q�u<[�Bi�3r蚣�˓�|�7�UH�|	âUB��t����D��-D��u]��U!�!ZIW]wJ�_�=Dk�W�}Dk5����p���R���ZEן�s���j��F��%n-��Sn����	?Q�IB�iq�
.�t-�LG9g�u��B�yrO��3��������B��]Bץr����F߿����W
M���麚��t���g�u]�"�}���5'B�y���B#����Bha��E�K��!�W�[�q��_�_!��BW
�C$f��/��j��*��h�
]�OOP������t=O�t�(��^�k��7ӵ���^w�7�����v��OY���H�?��Ю��8�Wt}��}������e�4D�<-����=���\q�ܻ����`��5L�N�0ǜ�������Gh�?���t�LK��/�����.�'|���':A�':�^!x�~��_-t�-�G�;p�l-l.��jx�{�*�����"GY�.����b��
]��{�`�#�.��v7�� k�2�[���������?�ч�����#D����D�!����m|�{��;p�co��S8�V:��Ns��r�B.w��8�
~ҁ7;�6���_8�A>��':0l�
R������4�.!��2�Щz�_{�-�4hR���j��G���U�?	�i2�_@8��'��8Zp1��?\E���H��P���D�W��Q�q�?'\��hSߪ�K'��8�p���7j��]W۸�p������)8@�n�ˬ����E�ԁ�!\AF�K�_I�v�-�Մ��z­�H��p���Q>�g	~�p2�~�Q�>����z�/�<�;���x��w>�g7+[�J�K�%��ౄ]�C�N߬l<�e�߭�P�� \O�!�K�W�i3r�ĿC8���_��F�O>}0��K��\h(YţO�E�E�n©�՞�o"ܺI�] ?�C$��L��s���mE~Z����	���j�����lЇÆP{�V��M��:տ�߫�w-��N[>	���s�~�p��_=�D-~#���j����	�f���N8�&�?
>*��S��N \��/��F����{H�N���1��� ޫ�񈟇�is�+�?�]�Ugt�[��ӆx2���W���~ང;^��A����O�M��x�Bث��k�u2�!�v�Z~��w�!cm�į&\qk���l<M8���	�3�NC������O��K��k�ԙ3�0D�Mބk��.$�Y�N@Q�%�)>[�>&\���Qӯ�	ב9O�#\ҥ�?��C������pc�:��p�_٪����M�%G���b�k�%���a<'�Jx�&�K��
����[ҾX#�p��|p+��?�s=�������i���K4����{��u��I��iuFlƆ�3���^u���s	'�����Y�G����1�p�gFh|�K���G^O�A+�U��|�"�����w^�a����7�}�J�f���a�+�RgG�I8Q���;��;��N������������g?+:(��D��Y�o#����S�U�x!\;��]���� =�O�$������$�%���A���S�G��V�O'�U���Y��[�y?���?���E�6�D�zu���Ex�����k$�ۄ�h��M�N��>k�Jyg�Q��L~��gU���g��(>Y[O�%\�/[�s�^�q1�i�=5J�^�����o�ϟ^��UԱB�ѳ|	�j�i�ԗ���ZWx�d�?=��|W��F��~UN_�Π��������	�u�g�M�'k�~�Qާ�g�&�}�Γ��O��w�P��.���s	�ީΩ�>�p�+�<� �H�y���HO�O��U�gi���p�֟/����s#��P\�ǔ�o�_]_W�b�w�!��⣩��F8q�:�G��W�Ԗ�$������Cẑ&��:A=+��K��?m��^��{��������6vQ���}����h��HWa�6_��pm��O�nM1��\ˏ��x�:{F��'�g��@8�3u�	��QZ����l�Іv��O�C��m�b,�t���
���N��8�p��p5��h��C�+��ោ��y,���SG��u�p�ֿ'�D�n1B���w�K=����ŷ������l{h��޼���B[^�O����@8]�m�+���}��5������G.�_=dyi���/��WJ8�'�}��鏫�W�Ǵ��a����Qߵ6�;wh���=]�z�K�^���aT�0�����5}�N8��v�-��h�[��Ŷ�"���׏�h��y�p�9���No�{_��ZO�Q�V޷x(�z|2Md�1���L����(�W'��?���g���������	�l;~�$M>����Sh<�m�g����|g��]G����,�F­����-��j���P�vy+w�o�W�b?SJ��Z��_.�?q��Y�O�ַ���F��x����p�����M7��O ���=^����cם^�Z�'�%��+��Vn��Zހ�5�{�pk�z���P�f/|D��1�����vM�cI��{l���u����"�<��n3������E�&�S1�����i��˾{�p�A�L�u�����5�Z��QG��y7�7б����@x��~&�V�^,���Q������Q�
��	��R����N>Ş��!�}�=~6��m�|�/�������v������$bd�&�фW���$�=�zv3��3������~K�Z��	�k�y���m��v�c�k�B05�z�p:��f;�E�[i~ɗ�c�i~���_���\B�R��¹^��+Գ$�/���x��[���C�ߢ��({�5/�g���;���;���	Wk�F³t��&�ƣM~���S����-��Nx���7�㻉p��~�I�VK��m������D���ޡ�?	7>o�_�	'���c��
׍���&��K%ʿ�:o8�ξB�G�}N7���x{�p���Cx�V�g�wk��k��#Τ�y͞�F.�c�'s0�2l{�±��I����x+��j���2�{��3�.m�XK��[�����p���S©�G��^�k��'���'�!�p�6-}*�����̈́+N���{�o���ӄ�H�=r~D<��$�W����� �����	�H�p��������P��%by��\=C���p�v^WG8�[�MH����	�}I�})?����30�����9�p��ޟ	����)�������S|	������Z�gvi�]L��>�^��p�.�Np�p�6��b�/���#ܪ�_��u�~�C�7��س)^��'����ĳ��s.�o������_�x¶7
�K	7j�} �]b��������p���z�-�k�-&m̲��w�X�h��/	�j�������!\�K���"��p�>����(�"[��"����c�9��9�Ƙs�O��s!�F����Y�k5��K8�[�w����ʣ��*᷉p����F���~�޿�ƽq�=ߝE�^�ו��|�s�W�����&���������� W��wkP��Ʉ~�������"��s{����N�S���H8U�oJ8F��Ho�獄K4y�F8[ӿ�Wh�n��z��R�袼V����w	7�i�?K��Y&�s|�Z�/|!�:�|�W�]����'˻�CI�ל.��_;�+"�P�nq�̙SZ�{��e���Ro��eƂ��򼲟��9.�ʼ���t���[�5��xNNaV����,+�|��_�3?/+�|��������99so��S�[�WJyƗ���]ZJ�p�hn^����`by�\���&��̽"gA��D��n�ϟ_\DWL�B���x�K�������r��&�.�)͵
��Oi^N���9��2��(2wqf�h�,@y�s�>�4�,ϛ�h�E�²]�����2��S:oJ�3>k^Q�a��/O�^\P��+uTO������XX��䖂���7F��Y��-�4/B�z��923<ť��ɉ��q�Ņ���vM�G�倉BL����'@J�ug���;E(҄���99ey��Y�7�f	@��k�e�-�6�J�1���)/�f\����Q��|-<�½��2N���nH�*�Ɲ+��)/�1]�s�.r�rsC�M�E43�+^�Q0?/��3Y��e`��*.��ųhMFYs
�r�Q<ޚz�"��G�F�\�6%����47�4/7RB���sJsJG���7n�b#�p*�v�t����iD�e�Ă���)�Y
J��9�S�r�Q��[���ܼ���J,�Y��x�����%�����`��T�#�+3�e�]�������Ҽ"�6�O����3��-6R8�bUQ�'Cml�<�aq@�Ρ�L�0]j|�yIty^�{՜i�B�V$)�lA�?�t�&c�x7�oZ��SL�Ќ���|+d�x���2c"ZM5g��/��--�Kss�D���x?�?��4g��0o>I�̘RT�u4w����̪��X�-��� 0A�����K��Ӧ iH\X���RƳOJ�9�
P�c�B�g북��0���h�H�h�J{莗Fg%�	�U@��Ai^a�q���r��e8OU�
����w!婋f��b�F"S���ꋲ�Y2�Q�n��PU�3P7P3I}H%Hʦ��$ h��>4�TO��B�[\g���) *[L�p�wt�'kNY�ی̼��b~���	Tđ��3Ӡx��ey�<��]m:�QD��	��E��R\=ü����ku.����J�~�x����S�]9v�;+c츩�����yTBL��8�7n�7/lPM+�\$��:��&-V��	��y�K�2�D��ʬ��(�������m5�vg�(�CS����U�5uZyaa^��yE�ujf���ȒK�ɛwM^�M�x����q&�����B3��,�-��8Ɩ��~R���Z�e��О��'������e�rT?� �I&� �<c��@��S���Y+ɛ[�_0�y�V�����h�ɬ�D�Z-��O��Ț4��qc�f]5q�w��`�Es,���]r�\�Zqn�pm�,�Ф��9%�n�M%�y���Ͳ�.O܇`��7!�c�M�+�[Z�[:��m�z�"�%J�y��'!�0˃n����^���|j0o��u|zay.m+(�n�V�cMB�u�����R*#��/!���Vi�^}'�ӤV�5ehTXЍ�q�� ����x������Ȥ�u '7�.�@r�����Z��v�g6p,dr��d��Q)�5 �i0�4L�a���+��i�x5��q��O3D���Ľ+V�̼�2��)����ZK椘j��G�t^��9j ۄdm��x=�Lϳ���)�5#	XS���b��e�攰�D�۝��-�o��髪Y�0,��&�Q3���(�0���X�k���Ц�*�WP�M�:�* #�w�ej����Ҽ��b5��KV��Ť$�>G"�Hi���/�aӥmk�Z~,ã?tlD�]ݴ���x���5M	����+�>����6(�N�_;��������J����-�F��y���Cs�|n�4�x�k�'C�2u�6��HY�w��g��0�d�wI�W��:l;��尓J��4� �K�������E�BG�ֈ̺bA�tB<������o�~�"��.(/�G�5�ߔ�X�Bc���mٵ��~��ƈ6>,�L�ˣY�,�4���ӳ�{���`��g�A���pU�*+�o�$���M�dW�3��������pn�^&^�7�m>=�lb?G+2D�4�(	i'1���H�򴜒ڢ�o��"t�,��6E��τ�)R��p��A�����(dبS�N�����0#kµ�ƦM��p��E7f#��s@�I7�c'{��tr��T�gii�iR��������E���,ꖺ����g��R��f��e��E�P��>[;���Ψ}s�/t�6�h���y���i���d���:�	[�ِ�C��D4��)���ȢG"�
r�E��3u�۰H���.��%`�H�ybkJ���y-?�C�ڧL��tbNAă�2gԨĜ�B��k��P��:��@f����'�р��^Z����|�a����P� ��~jK�$���2�G9ċ2���r���B��3չ~_{@6e`sI&��l�0;$Ҏ��ϪB�4��L3�)EԭEs��ye���<kOy2�2���O=#
�:��c�hU��?�c�|��9/7t�O��U6���'����"����̸��R���pL�d`kwU~>v�*����J�W�4��S2�>XX˾�E��Ÿ���y[����rՓ�<�Bm6�G�r��k̳�8�Şk��`�F0Mx=��
��	G�#���BS�� &O�}�h����2�f���#�[i�b�zѵ ��aJҷ+G���k>0���E�Y���L�H���#�aUi�����RX��48|m?2S+�a�q�)D����	�rk=�2Jh�y���7e�������-)�܋/��U-�8�yEN�y�4�J��yJ��}ؼ�v%6u���K�O,�Qi،�|��2mI�F����#y���f�Gx��b[v�l�XN���d;C������%�H���5?Y>}�ܐ��[w�w ��?�͝;/.�͆6�{D�D� j�լ~��s�q�n�'?���H&��#�W��JK�����?{3��Y�=�Q���������b��)�P��x�<�.H�J�eVJ��a5N߼��9㕟pE>��0��Gvf�~X��T��YO��t$/�DX������1���s}�aT(5�e&�^��x��I�<,y�x,ikM�aOj�e�ḿ�{C��G���BF=TG��"5ǶUm�ѽv����d-�+-�mv!ǃ��e��t��C��1��e��32�]��|��������?x���i��ߏ���������w�4GR�����Q��pc�ˊT��94���FX��[`�sd��o$9��R��J�o�o༇Oa8�;W~�>i�1�e���Z����V���T�q�����XC}����!?�/���9����B���d*��~>��5�k�҆H�{Ʒ�����߁t��	S}�
?x����?��5���6��P�(�?|m��|(���VS��`�M�?Q|"��T�n�m
���(�/×4�/�O�u��]	���
_��������� ���W����_���	~	���j}�T����o��8�T÷5��}l����[~��S�?�m||Ç6|�gt��|��;C����=�f���WM�o���]4�,"�	��E�N�b*��1�o��k�J�k���_|5$|���8|��&|H��1|�Ï�#��|��; |;��T�R;L�_~A�{~���yS�&��b����3�'���|��;�ф��lS���l��/f�چ�n���om�w�����ZG�IS�ȅ#���~��|'o0�?N����|	?��ɜh*��o��w+����v����:�<��*|���2|]�7)���oh��� �������;L�;~�����o�޳���:���-S�Ʉ�I�_o1��K����n�����p}w� �
�o��\������(�3]�J��^���/v�2M4��e�w,����X��������ÿ(|�'|f�w|��g���p�7�O;����Ӡ�~g �M��|5[�+�o��K~��>���>��/����~f�2��[�6�{��
���e���c�� ���k���ݦ�3������g9���:��7�������c�o��W��T����>���<��ß�+��-��������C�����L�����{u����T�7�h(�pm��9~�1������M|�_��o.�.|�?X]�2��r���_�zS�&��NS�& |������9��o*�_,~W�S}#���1�G����	�w������P���f*��������}��s _p��'~�n�r�����	�Z �D��5�\���lE=B���
]$t��
��B���#�V�
�+��Z't��5B�
��Nh�ЍB�n�,�Eh��Bۄ���)4(t���{��z@(}�h�1Bc����M:\h��$�#���,t���B�M:A�d�S���:K�l��Bs�z�
-��H��B+�V�Gh��BW
]%�N�j�k��Z/t����6
�"�Yh��V�;��	m�!�ShP�n�=B�
�/�PQ��Bc��
u	�� t��D�IBG)4Y�(�����*t���B�
M�!t���B���
�-Z"�+t��%B+�V
�z��Z�+���Jh���B�]+�^�:�B7
m��չ���#t���B5+-4Fh��T��N�.4C�,���f��Z(�N�j�k��]'�A�F��B�m�"t��6��B;�v

�-�G�^������Gh�P��x�	B�M�$t�БBG	-t��T��N:Uh�����f�Z(�D�W�"�K�V�Z-���B�m�*t��6��B;�v

�m��V��БB���:Z���B'�,t��
��B���#�V�
�+��Z't��5B�
��Nh�ЍB�Ȟ���|���ǐM�xԱT���qd��u�s��{��(o@z2�w/ JFy(�t!�����T(ړAɰ^A�4ɸ^)t��:�����Vh��uB�����L����h{9ՓBv*�M&����$���})�w�+��7(��HO��X�G�dP�|�E�Si\	= ԸU�h�1Bc����M:���)��$>���m%�4���E�I�Y��4���-%#u�G��xē���&mX'/Vt�И[�m:�VE��K� J�VP��V���r���.Z!�Rh��{��
]!t��L2��h��0�6+�?�����w�_Q��^Dh�TE�z��B�:g���*t�г�R��BzP�tE�$�s��]�h�����?]��{9�o���?��Q��&)�63�H_G{��g(:S�߄�:d�����`�{������ͺ�>Fz�8�3�?�}�s�,��&�R��
������(�e�?��J��\����E[N�hW+�(�6�ע�7i<MW��L
����vQ���~���4�C�hS4K�l��Bs�z�
-��Hh�I�
�}E�=��q���C�~�;P� .��0�����3�����2�$��6�УM#�z�i$.4Qh��BG
M:J�h�[P.m�9ӆ<��O�X:�4j�/?2��w�i4A~�	�C�٦��y�4����Lc50m�sAn����c��Z�M#�i�P>m�WӦ<t�iL@���L�E��ɦ�,4a���Bc2��?�4zP>��٠4�F�\C+�*ˋp�{��3����F�X�tŦQ��4.C��Z��B����Ɵ1��J��~ڼ�4��+zh����뻨�Pn�iT��Mc�ݦQ���|�4����A�X��:��A=1��g(Z����\���i�@5��ю��q6���H~T��AP��4����^�C4�@'�:B�y��{�n��hm�y�砗S{@ǒހ���L�蹤������L��}d��>I�(�-t(�Wo��\Z�@ϧ�
�q��t��w����8�"9����)�u��^O�	h���i= ��� ����Z�AsI�AB�>�Ǵn���u�Z�A��qz&���e��t�_�+��=���D�h��M���E�(��6�[��-7� h-͇�&��AZ�A[��@q`Jz2�V�/Љ���2�X�<��A�Ҽ���o���~���G�.�A4o������7��7@/�~=��4���si}��������WAi^�ͫ��[�Z�/�Q�Q	z'��C�蕴^�Ӽ	�w�Х4π�1�5�I4���X��4��CVѼ ZB�:���f��c�_@к�(���z	���ِ�����9�O��@i�u�>@�t��(��@�~�1�3Ы��@q M�|��4�Aϣq�N�~�A/����7�G��@�S���:�:���}�7P��M���y�l�1�Ag�g�gQ������3�Y�+�8�w���m�=����|Yz��N�?��i|q8�(�V�@��=z7�+�,W�OF�S����0��O�=���西�q��AtW+c�$�jd��su�3�D]u�qz�A`W-cx����
�8�����1n=��ٌ�k�̐]��$ǃ�ԮTƈ����+�1�rO6p"c$��A].�x���c�.�1�zp���sO;<�~�(�S��g�'L�Zn?c�Y��g�'1�:n?cT�Y��g��p�zn?cT�i��3�/�z���������O=��~�`����g���n?c��	r���r==�~�`ճ������w:���ne�����x#�?p=�-���u�����k�p�W0n��.a���8�q�?p:c~��{]��;����w����8���b����`����s x/�?���~�n?����~��g%��1~M�S��g�y�p�Ct�zn?c�����g�'��Fn?c<a�4s���Vn?c<���q�C��n?c<�����!jO��1�y�s����=x���1��xb�[�+<.�F�x��I �g���$�1�Sh��Z��*O2pc8��.a���g3��-�d�t��JO:p*c<)��Nf���d'2F�z<�.�x��)6�k�����7<�~��jO5��1�*yj���Wr�s������3^����g�����g�����ϸ�����x�?��q+�?����n?�6�n?�v�n?��n?�N�n��<^�����ws��2���nd������~��:����kC�<�����G�0�N�f��=������2+�Y�Ɍ��t]�����z�\��� ���gp�~o��~�`�S��g<����M���3\��g��y�p�����3FS=�~������tO3���T�Vn?c�����g����g�x��~Ƴ�{���!*�~n�7,`����`�yb�[��{���C��D�:�K�G �2�N�`�zF�0��WO*p6�������p��2^���̸��8��:�`��`��F���}<������[�����[�����wp�s��q�s�	Ð��<sFO�����/M÷�U��o��7|�tS�ԁ�������O��t(ʷǼ��,���_���d�+|H��\�S�I���ªj�_�k�z��I�K�֭>o�����������\�0�>>�o�Vm�&��(�BR��0;)�iB��(��z{���j����o������'�����_����͵�����_z �4������zM����r���A�����U�q�x�)0)ܨ�U�P��v�
���B�����F�c�lL F`�H�7)�?&�Һ�x"���HL��r�� q����������A�ޟ:���"�X9�b��
���~~��y��P̰>��c��5ϵ���hHi����޽��M�����$��`���g$Š�`�	�����������r����d_�dT�RPw��1�" ������qU�.Q@�+�K)�S��i�\�T�c-2����F�;��0��I��c����S��@� =��Xl�I�;�^�1�5�ǭ�ے
u$y���(����fK��
�Ku��#����
��27YgP֮9$�|�o�Y�X�I��C���m0�����k�I�ϭ�%��U����jk��ҿc)RK�igFс���H�=_�ݝ��+ۉ�I�v@�tt�H�بHz��WN�Y�/���ʉ�+}����������˃_9��O_�@}i��ї�_�����Зi_���r�W����X��8A��w��}�&����c�k�Мh+�I%J��G%��1A�c<�cwO�����(��nt��X���$�o{T�Q��g�a=7R$���蹏z�z��:G�� ~�ɊP�8��/���o����P�l���g��j��?D9��������^ƫ��7GA?�<���̣��$��^H�pυ��x���0WXX6�ņ�rK���K��mI�&tW���f"6��'��H)�bX���\ѵt�2���,��i�J�P�|.W�W����گ&D�RTJc���Լ(�ٚ�Xy���U�������Թ��.{�+ك�/��^Ds1D:��W�k|�{��e{�s�H�%6��� )�Kq�;y��<q4��)Yf;R�����xS\%Dx*�O�؏>�:�����ƪ�1Fz/x<��W�ڟӋ�	��4�pʉ1*kt�CgP
������)���������q^��E�]��"}_Lx|1���k^&b^@����y�m������Ϗ`�&}��g}������3~O�<4~���3~�܍�[+�0�>���>q̧��"�)��N�܍n�^a'��Vk��͒��ʰ9�����ֿ���"����o>>|tAft;�sF��ϸ������P�����?u��ǋY�vB���oF�D_p����LK��t/�k;�ޏ�6/=�~i|�q���x�D�=j�px��0��=wut��8�"�����r����$b����#�����:�������l���e4Mĩ����`���h#�w�Ǝ
����/X�E���ipsh�.���:���Q��5�'� ���t��
�`e�V��k�GV5�?GSf�6zkWW��ݏh�)k?5�m[��?�$��\�)HR�q�q�)_�����Ϗ+���V���c���MmKd<[��T���[�x=E������b�'W��G�{2;k�Mm܄�j���!Goz�����>�H����~��`W��j����S�^Z���ʿ708@8#���4=�����r��8�u~�uO���QTv��)g������ǭ'`�rǇ&�z
�_���@f��>��t�R/�KiT+:��C���CًĐTkʛ����}�ob�^�g�Po4��c�AdƷ���(Σ������Ԉ����tNՂ�M��98[����P�Z$�F���l˪����]��O�l�B�A��f[;�<�zŚ-�i�|���������9*��X�Qَ(n�������2�p#ln�1I�����گ��7Go�Ǩgt����)`��Y%[>0���$[l��)�ߴ�: �x\�{���ӹ��?�_����'���ٙ���@����?ir����I��ǺD��:�
�R�N6[�c�W�'E�3�}ǻ:�J2��ݽ�����*�*�|Bר��$ԕ��~�@Z��;a����k�U�����E�f�o�Z�C��w��B@��f��W����<Y�uۉ�Z-�����S%�m�� D��mzl`�˟�A6oקd*=���f&��H����ï?�,���y}����d X���jbz�����Ƹ{��K
�<�1C�Q�K�V�T೻��#S��u/���@�oIס^���탆�t2�3;��k�^�s����L�k2�xa�hv_�O!��;�⥮��<���!�(H'�!��kD܊FbP��zhj���ˏ��wf����%�ʾ~%~g(~����@]ĸkt���E���^h�f~��S(�6��������'������.��Ŀ���j�I�W�nݡ0>�&q�`���Z��!}ex��Z���g]���������8�v�E�l�!$����6�Z�ԙ�lTp���ҔFf�:�}��o�U��B�����:8l���oi���j|�kz���[�k1z*�o	�_J�c�IZ�t=�s8v���T�p��.��p��ˊ�3-^�+V��+��vi�Һ��|i�*�T�!v�qQ2�u�]\s�uЛ���+o�����Ia��:���則����RN�Is�MU��C�r��ã�-�݇�I�����a���M�xtVm��§p*4S��n��:�Z6ꐚ/C�KU�����z���=���Co����7��P4S�j�?�t�j�)]k���!�����G�gv�4Vm��i	c?��ݕuК�l�󈯮��q�#��Z�b{aG߹`�a���:w��;���E����������u2�j|��U�i���z�����h�P�sަ�gb,�]��)b��T���������O�ﲵ��o>Ќҿ��3�O���-�{\���-����E/�l�;!&�rP��[{o/�G�_%|P�Q������LM2�v������}�2��<K^��L�&�*���M.��>�1�uz+W4�6Ӯ�tU���MߝAʫꋫ��&���kQ`\�mQz��w���U��L�+x���*ݾ���jG�X~���w��u��74NT=�����9V�綝ROWB�ڣ��������� *x-tNf���N���s��d����y_�=�Py)������W�E�w��f�y�N�o'o$ڙW�M�����o��S�*7#���f�[���ȏ�xm=ޒVG;�F��+xP��`�gM4Y�qU����F�6�b�$O�	z�Q����d��J�\Ê�����,n�6��q��
e�s��������+9�eZ(ߩZ���V��wr(����(ۻa�gY�3!��$�c|/E�gưL����͎gav��	J��m�]�鹌�߿��_5t�na$�'>��n.x�!,��v��X�4Nu"T!���ȉ 6;��ȉ6��4$r�ܰD�ލ�����D�GN����(���)�O�]�b�=�97rU�z�!㢷H�II�sq�R�>�t?�N���Sc!e�_��� �!Ϡ��t=�wMI*5�
�3[8����J��)���x)��w��U��nO|��~{�g@�Y��1d/����\J�I�����(�M��(߇�?m���*[g���J�J�:��2��*j��,��r��[
��x�m{��F����{��qU'��Vf�aD��	����x[�sM��-��S)[�o.ݗ��Aw��mT�Xݷ�7V*�7}���i��r1�x;�MD�Z����j֩j��*�$P�lɡ�q�n�V��G�U�aS1w㈻�x?��q&��m��j�K���51��;�z㪺���XKܷ��9��&�woR7�;�@Z��i���~��N2�6�?J�G�1���+ϣ
h��O?�}��I����jKӦ�S�&�0gMݿ{M����%-Ԅ���N�w
�s�BU~��U� �]!����2N�����6s5y����x��
U9�߶^�olAU���P���[	���7+�G��n��U�/w8ԯ���tȶϕ\�!��V�`8�0²�|����_1.*��zf��ֵ:����Ma�jES��������P�־%&�706�W��jsli넷�ZN[���ސO�u+Q����~I��RnP�j�p� vE?��>��f���7T�4q=�ۭ�th���=ig�Ɛ�"����U�A07��GY��@]���{�%�g���]��bB��p#�m�R��#�z�rO�ʽ����������s��a?���]&��Z���|a��������]4��[��鳻&�p���ˏ��k���~�$�xW�bc�v�-�U��C⫫��y҇�1����d����T�,Q�{Q�om9fƬ��~��Ő�����&{��Ǫ�Ma�!�I��8��54�$��!;,3�l�� ���^�c�pLEU ���l�P�N	�7@����c,N��b+����=��V%,���n	���-]��ϥ'bXA���9i� �c+ùop�;C�<�lߏ�/�<9�����V��0J��^�	�#�Jު7~a�?�M֍� �V�8YE<��Z�������2 /��^���F�����k	7�L���T�9�Xr��﹇�G|�=16�wwl޽�4"Ly5tl�x�����vl��j�c�|�<-&�ǕS偱���a!uz�R���]�ҷ�L��\�����w.��Mc��"��F�:��g؁����V>*W�C虏U!�0��r�����x�Fj�>��A~w#���W��ď���ƈ[O�S�~�|q�zwcJo���Mq�˷ĭ�l�ԑ��C����R��o6}�p�W��c8t��́��G�l��qm��u�~N��b6}�������62 w��v�R����P��8-ǜ4_��� OO���W�<:�7Pf����*���
,�''��=9��H�a�;��H���U�ݤJ�L'o<���*�jk��֚���n�qz�����x������&�l���QD^�;�HK��h"�V�=��k�cy�z쐐 ,}F������ݗ��4v�vf�����,���6���E��B�	�-��<�v�N!j�3�1�A����^W�80�Y�8���q`vw�80�y�80��z���z���edu-�jM�]	��µ�r�T��\w�")�d@rWp|w����W!|i�����a��Ri���>���ϵ���%Ӏ$w�U��5 Z��z�hR�j�i�ڦ]	G�>e�.ߜ�iW�ѭ~��;X��u�o��d�,�;�ri;���h�I���������$.�XU���϶��g��	�$���U�n�^�|Kmm��������]����ZE.����7�N��o���v�a�fn�<��)�k	���@f3�B�e$��'��ZDE�;���NT*:Q���Av���o���`=�W����������/,�8!w�#=|i��a���%�`~���w�Vne=��s*��{!��FL�<w���y�вH�:��/�f�~�zw�!�F5Q?�~�P�3���>*��������J?���7�,�6~��eȫ]�U
įC*y]lq�,�$��Q��Itw�,�k=?�t0U���#��T*�{M��k����@�g����O�I��������ד֑���#�=��o�����V�zm}�iv�/y�.�_l	�_J�3��H��q,��-N�j�5��-���~����3 q�<������Jm}s�چ}��WJ�C^�f]^Q��X߆mv
���R��_:����s�a�mF};���mH�Dn߾�[�&]n��t8=nr��[�[=[����)/�7gC�.�C^�o�µ��ZhQhe{�����l֖ۦ���lo�A����5{s�no�۲7߄�����|�ao6������^ߖ�bӱ]����ȷY�ӛ!�f�|��f�μ�ٙK�Ҹ�,U��V�2�Vx�E=��ùN�k�1��:�ek�n�g�&Ү�͝��|_����9[��5�kb����Љ�=���N�i��熦���j�+�H񰼛���m� ��T�:-�u�f���Ԗ�-�l�NT6�De�NT6��!�F��/9�кt;���޶*�8�}�F7��Fo�l�S������%T^���Q����D���h�6@>����~�ъ���ٚ{��SOl
�GĘ�y�8�z>�8�A��ﭒ��[���9!��K���{4�P��/�z��إ�3���l��F�G_��@{��ۣI/�`{tl��um�E~�Ɓ��_ltڣ���=�wC�=j��^����!y퍫
�t2s��@�v�!�;�/�E���۷��h_�e� ����}9T�N#��{��*M� ���g��G�C���̘_��X����9M�������IE���k>������x9>x�o ����}/�/=P^�>
+S)u�C7���D�MEa��� �7�Z���%����	���)����_�����,�z�?�XѤG��{�M�󽕥�w��?u$��NX����?����sγ}����;�?�?�_��靁�������g����w�t�+ �/�4�������~ܠM&�|���sz[�n�wP^}���~8�A�����E��s��?��oF���?�(�/���ntȿ�]���q�?s/@��oy�f����N����)�Iϰ�S�d?\�+���"[��Xޒo���O��f��[�[�j�o����������t<��z{~����m��{������X���7�#߿�w���G&�O����;j}D��.�4���0�^�t_�Z��m\����?�ɗP�o�\��[�yʳ9'<���ԧ��\(�/3�i,��N2J�B��M��g��G ��ly�l��{��޲�N�ޕ�w��|O}L��b�>�z\������zq3M0W��7[��ͼ^ܬ��q��(�N�fZ/�o�]1�Nhƫ,�~q��§x�@���l��=�5����Z/���
[��q��O���O�Om8M�����N���O����IO���D�E�-�Ʀ�j�8'�z�FWhш$�o��;�F�������\C�Z��-��kצCg�߁ �R���G�Yc ��o��*�{������w�.F�p%�SCL��F��c�T�K�)��{�}��m\΋�����4W�El���_b3�A��	��.w�?t�� ���_���?"�/�!��#�ߝ\nӣ:���.�rn4"��*���O��s��K��ߖ��A.烿G�����<�������w���?P~q/� .@A��=� ��H���x��q����������{����zpMD�F;�[}���b'��7&"u���_����o"n}Zl�����9�+8��5}9��?py��g���������/|$��36?�#��0�|�e��gjD~�F�Ƿ{���K��o��;6���}q�d�[���i9��3�K�bߙ���Ȗ;�Ԓa}���2�zG�M�����_FD�����R���{��7+"�G����X����7;"A')�}����U�c�Ӹ������X~�f���f�kO�D���BlM���Z���T��ž�&Єx~�,�]���s��rXɫz����}��k|�ivZ��D�;=A}]߄����/k|A�X��.C���� �jR�����xOkG�=��� 1{j��O�{Z;���Tm«���I\¯Y���
�ߔ�+��ZU�{b��=d�I�N��%����wH��!�0{���	$������6����n�a��C�	9��yZUcy<G���Z��l�J=��ѻ��7
�����?��9���K0���{�	��Œ��g�N��k�A�X�a�uz����ہ卨?
����OUe�:q�T0`j6���������bk6�K��記�)�)u����Q/j�.Fv�rd�>ȇ���r�pH�@LfG��i��>,��^�`��*�����Vݱvݿ�u�E�;��n���u��\7젚����R��q����Q�d�8H�9xf`�r�Zd*���#�w\�Gݝ5˿�Pwg`y����n�Q����Q6��� �/g�����(���p0��`���������a<�p0��`�����62k���k�`����s0�/�D栙9xO���8Ȱ9�l`��r���z��u�� �@�̶9H<0 �Bs�E���7��q��qq�ό��u}�e-o��疨�x$�������,��Κ������ �I)S9��������?��j}:	��03�"T�{�[�����HA��f�
��;&�n������
�}O��[�{%R^���#�����_v���V�(g����ub�&�T^��rpȵ�|�p-m����[��;g=R�r8�1F�,?� �WeY~��C곕�%�G�BK<�J<,���Z���_�t)��J?�o�*�ʰ��V���ү���,�)��DJ_��K$�Z��_{W�e��{+�?��f�#}sa*��6J:�����{�RL��kC��05�n4R�S8r<x١*'��6B������׉"O��7E�X�.[����7_Qq�+�Y���?$Yc���B9��y[����7�P?u4�r8
s��X�iO1����dJ�p�����Q���.�8�G�T��P�\Դ��CvoO�/ӖP�Δ�e��_��P��hdZ�eZ�_��P&x��	,�L5���2�u:�򥠓h����_M;B9��T�.��š�Vg��P�?
vCu��r�4�E�J�:B��a�h@��Xg(�&�C3�g���X%u���ݡ?��`u�r|bJG�X��P�?�au���O�C92�:����ǆ�qAu�}���!�2~�:�%�wi`Ú�DI��0�,7�g9|ذ6��:*0L��')�Tc�
&�i�r_���ʾ���ve~������ ���Q�BnF���?����{����pp�^;؇�|�\��A��g"�9��'A��7sp��v�����`�?�Owfi�߮��v<\ޅ�+8��+;���J^����l-�O.���Z��w~i#�|��[��Bpj�c<����������]����[�����%�bS���%�8�u?S���m��h���1C���!Ý�3��2�5����,�{�2vY��D��_�.�j��9�Y���v�X�RPL�������`¸e�<����ް��U{G�3���f�����U۽��cf��-<��E~�RQ����c߯Q�/���+W��������P~���.����P�|T�
��Gk���x�Z�Ѡ�����L��?�~Me1?.ՎX1��4�%�4'H�{)ܾ�n��?���׵�UG8^/�2"�����;����,y���y)p�������S�k|e�r��G��g���$�L�4�>�M�I��&���G��{�-��˳ʿ��qʉ#R������������(�(�hIp3%�o������t����$��'�c�g��@�:q������VV�_�>��7q	~w=��QI��S�>�+ݖw��ej�E���)H�8�e�kཱུ�m�-r.+^��Ϫ}~wcܽs����j|�tږ��#��yCM� ��mM�<�2��i����]�̫��4����3qn {f�5*�筛{�_�����}��Ӭ�+�A�+�%򉜹_���&RQ�(��d+W*�d�G�������WG��6�i�f�l���R����>m�N�!P�='%�$h{(�i�j����b�C$s�E������2T�p�rLB�6y!E�ö�z��v�Ŏ�6Z�h���"���a�v\��r�R�.[�b���Z�/��<{?�Hi��$+nEcͨ�����p7@$���_�f��TH[kp�J;������R����ЕpNa�}{emȷ<�(��/EA�-KB�ݫ�J�*-]�����}2�(�I��~���
M�n�����������]=���)�>��?4��,~��0���:�<o��'�a~O�>����|<�^�㡌�������v<܁�����m,�c䅔ޫgm�߯�P�P��Z�BP�
������e������l�����[>mv������~���$����J'��i��G�Z�/���̓�P?a6o�[^�iD�6r�X#�%���	X�Go�^�2�٥xL(�:�`=ͤINod�U)����_�7j�:�7������\0��W���/������C�Op/�|�W��x�F�~���d�R�%��{ٮ�7�b��7��%Y�A�^��`R)w���Y����rY�\<�Ƴ-����������نI��xթ�Zw�2��(���O~�"��*H�����&��F�>�]e��d��?w�������i��M��@��߅��18�L�DZyQ;A�?�ʩY�+���v?N���л��7���W]Ү�$�۲R�Y�E"//cc�R�.NP�-�s�μ���Х�F����0�r'K�����?�/�,g���I"L��}W�i�� �{�e�1�|ls��[��L�U�+[��04��@���
����^�'�a��(k9dQrki��A#�����
｟����Tj�����98���*O,��u4�oIR,[H+`T8����/��	��& u�o=߹_�4��l�w�zp;;�W2�����ί<��Km�4�����b��~�����%-^ٜ�/���q�95�%߄��w���۰�ސ��S+}u��׀_Q��&\���$k����O�6�W�c�e��m���p����4�L�p5�<���y�}�����Υ�{aվ�ʻ`^**ދ0���i�5���!#hj�r�/��cX��k��Rf5�{�����?���Ux��Ꮹ����@���}!��|7<��sm#��W�����#����{a�=��
��x˶n��<�t����D2���'�Y�DS�0����*�F�i�������VO�������`���P�k�θ*Ƚb��4�G��2�E�ju���Tp�}��G�'%�#?=�?��z	��)�_-�wHT5<8���@�����3>���wt�$�|-K�v���ۮ��di-&T�H� �{Mf��/��5�A���~60޶-�g_�����K���+^h|S4��q�� jR��:Xgi袘B�u�I	�&�O�t=o��~��_ƚvr -�?)V�1e8|q�.Ï]&�t��"����b��[��1�g��Vc+��ĺ&����4�����M��ѽP<a��������!Y�!\����R]��6�KY�����uk���E�u�dc��u�����TXkom����z{[����*r{�:�kڪ�����ů���ů���ů�����z{�։�^����ꪷ���n/�����������C����py=z,��^"o�'��g��>�60̷5ڲ��Bhy7�(��
.�<CW'���̂��q	V�`�W�8�yE<s�y�W�}���KH���ʖ�mQ�{G��k� �c7F*vE�T?5n�2[#��"�-c;$�=bl��6;b+B�H'T��"ƶJ�VGlm� Jn��#�6F,�YJ~1ϙ�~w�f��C�<�
\�Ȃy �oG�?�E�����$��,ٯ��»����X2:"�[MK_��?��'_���)8��ӷ\
ie����i�l�7����q�1�J<��J�6m��'3a����k	d��d��}#qڑ����&$%��Ѣ	ld���x!��ܠ�����0�<Y�{ l4����>��b��}�~ �dp�&���#dw�	��d��������.���:ˎ18�ZYz[���[a�^.��[����\|�n/�7�I=�
.�K�Գ�R�c�����.�QUW���!h4AQ�E!X�	Il�I�$�\�y��&H&q.\�@tH�tDS�J_m�Zjik����Zjå\,�)�-�����X�����Y�=k�}�93�������;3����k���>��M���j�Ox���ީ�X�o��}:���8'-�?�ݡ�sbߧ�J.�d%�'V�sA�B>�c�h�]7�6�r0r�{��(?(HT��+<!G�[���"��hWcu��g�M~[{,�bs��i��9���?�L�[!���ͳZ̮�.Y��TlDi8�b#ʩ�1QN�UlDy�d\����GTރ��I)fB�E`�ʲ7��4UݞH�)@;�`��͂�E�O�-�a�)q�	OdM�mE�"|����� 1�~	�~���v]~��sv_A�Ncv�������ޢ\q�{��G����-L��R�r��+`0ߡi��ڦ���֤�o���?��pc�׽�r���(���OS1r
^�!�L���)���<�S՛(��|N<����[a*��?���p���7t���혔oG�d��z�O7#	Q�(ߪ!�K_�YR�Y�5-�pG�#M��,IS[����09|b�$ru�y�P��vE������(|����8!�YE"
�ܪ�v|4� �L�;T����c�c�|gë��͹?
�����5�;=�ŀ�|�Xߑ�hu"�����Z��%��������ed9����Dȃ­m�/Ҕ�P�JI��%n�zb����(|�z>�|��wҔ��e�H{�Y����)	��/��5�̩m�?����Kr�Kh���*��D��!Y�;ժf�$���P�:�'��t�T�ц�h]�o��f[����	>�T��FSq'�ڏ��%%lj�PnA^&�jq�L�P:ߴ~��LZDg`] �G:F�PY)T�g�
���7��uA����$Y�^6�7�lC�x��eȳ;�I�G7d�,o�x�^H�Cr�,��K�6��QJ�n�K�d#�r�ޠ�R._���)yx��Բ�.���������<�s$���,wP�J7
�A�Ca$�`&�/4�o|(�H�n�l��^!��l����#�=�K�#{{�[�#Ǥ=r"�=R�!�=2/���1n�D�)�h��%U���PS%�1��*fsc(���(ƈ�}MŚ>��g�� ^����')&-)����G"�͠�M$�b؛O�E�=::��o�u
�ُ6g���/;�$ˢt�Yw�6Ngg�A�>��<wɃ���y���S��"a�	�S������>E"@��Lu՜=R&��K�.�H,�R?��o���o���N�܌6siJ��>qC�!����M��P��ŕ?3��y�y��#��_4)�v縟�90��v�X��+�r���w����
������Y��kI!�����[��c8��Ǻ��/�v���˷������]����1�7������ߋ����e��E���(��n����:zׯ���������[ro��~j}X��5���5���{M�MW�})]�?Z��Gך��~�c�����%�������Н�6��]Z���k�~*��3���S���|�7a��&��赿��_x��{25Vw��#�Fl�0(�n����[J����/���JB�A�eY�ܳ�r�9��Q'O�$CU�Uzu�\��c�{�L�i(�̳��[����k��c��D��NN�E�!�cM�+�fz�q����s��������L��q��$p��\Qbs��D�O&���>��o��ѻ�+����#�p���M��5��c�,��lx�x��d��RL�&U	4ʤ��!&�"�Q��r��p��a��O���,�5��҄��5��<���
*� &*�����q���g�rMx�+��S��g^�
�k�o!���9!�5}N�����4�Cl�=���2����}V/��!H���ܨx��3�©;�=�ޓC��Z��m~�j�'�,a�8�>��hB�{�	5	�C�J��s��
�Lm6���U�>Xe�O�����9�bk<�
N����	���?Ŀ����ت�m�-���ʒs9ə������b;�,y��ԻA��b���n݀t�^|C��=� �!�Ծk>Py&��ȗڕ����e�W�o�_w;�>I�q~�w$_�^�y�|��~�|?��i�,~6�<060>9w��X�w�J6dmGơ���-Hh���W���S���o��	�Ӽ;����}g��P:�	{r8�
��X�$���۞�Ȟ��[�ON6�h]L�j?�Y�~�s��9ɉ����-Ө��	���\͛��E��GQ���d=�OP3��L�b���j"5��L=�y����_M�.�q�_@�Q���b��|�9���El��[R~�J����q�-��'��+���l�ևؿ���B�8��<誚@?�S�c��ݸ�sq�:t�ef$�z��!�9�j$il�@�E�?M��:�3hp����D�ݕ�&�y��[����$ߝ�"^?�:M����6u��n�k9�>���I��ת�h��H�����ĐN3H�^����jA"юa�_{QЙoE܏)�Nz��D���Ck��Jt�/�P��"3 ���Vo)�8�J^Q@A�!��ߝן��*r'��.�-�C��)z7=G�����'ˁ8�/��'��vѺ�t]��~r������o��]��g~��
�胒���x�<���P2z�_P�{�J�����6����������4��e7�W��D����5Aok�?Ȼ���������_��]X�o�}cK�_��nL��c~T_>!0&PxP'ٖ�W�}+b����D�^�Gv[@Ʉ�����3�SC4N�	��^� ��D;�t�M��mE�k��{I�T�*���P�^�G�륉��D�|/#��z��8?C/%�J����{������r�c�b/�n��']f���8+�΃�7�s���1'��K�aHZ� I����RJ�q��|a�p�:^8��:O�81���|�S�>o�5D��=�PI?d՚�\b�s�W������w�Ҭ���~x�2�~(�*��CJ�~�0��d���*F�R��¬|�釧+�ꇴ)D �Jy~���N)���W?Hh�d����2qe�G���ܖ��{ Wj;���h����Eu?BQ��;J5�t�	(���L"�udl�v:�Wx�b����NHe�J��e�#��cHu��P��܃2a�f��	�H�!p!w���!Ȼ�܃�p����2ARVao�C?%<J"���n$��?+�x���c��i?���c�b��#�Z�.���|��S{u=�W��=�UPp�)��7/�������/>�&�*Y`o<�о�TYt�怿�9Է�����S[��������C�|��/�)��Rb��W����m~�&a[p�(�4
ڭ�i�Q�80�����0��(�x�ZwA�%���;!��h�i\�qPqV�����'��������z������V����6A1V����y����d������Q��d���]���<к)���/�!g���2Z��b름G/|�8�,{�����
⛭��w� n��?�K</4�����_����|�^�({-��]&C��V�ˋӷ}�����M4��ٓ��הQ���]I������\���3+ӷG��o�d�J����>r}�hed}����7�]����o�x��n�+8�V����b�ȱ¬o��gD�vڊ����U��[:�z,i=&F�5���ٰrK�D��������,��1��֟�F���ӊm���B���&m|Q,��k5����?/�믿,3���o�޲�믟/3���+������ח�=i�u�����kCݖ�7 �x��o=B�4i�%��1Zo%1	.��T�՗b�Q�[����++"z�?֥�VϷ�м.�^��羕Dσ���/��T�|�P�A���ã����Dٟ%T~��q���^��A��~|�wd�=.D��ۊ����?oK$��w��-��ê���������2�s��s	��q�f�8��r�,9�B]��\/����2��Ű�9'���`�r������o����GGz�����g�X����rS?S�j+�u3�*��Zf�矖����J�s"�~��'>A�M��s�p�sf$����4�Z)�GL�`��k8�9�P>�%f���e#���*���s�%z~����5L?���D�#K8�^^2R�l5H��%f^s/�~~xI�|a���=#��پ-O���8g��D�?o����k1����?�3r�ر�<���|��Zy�\t5�3/��Or���a��n��8�>W4���l����<f��h�E�oO_)���о���Do���m�P���%ܾU��ۋ
/̾��0�}�V�پ}zIT�v�x��O�`�Zۏ*���ٷ�t���P�[�>� ���ٷ�/����������0���wp��w�����׾=�����#��Q�[������}�_d��j�7�.ľ�Xd�%-�`��\~���q���m��me�ɾM�y��?�}�$�����۷����������!������"��%�q�.����p0��w8�y��|������D�ώ��Y��'���k�0ѭ7���oy#���%��k��1"��\�ľ}����L�Q!���Rq���C�?'�3�"͟q���/s8��l����)3��H�y������\N��39��Y{�Ο������v�8ݾe��I3H�u�y��.��i�E�oc/!���y��"1��$r���?OS6��4Yy�޽"�ۻWf_�y����ݏ����syQ�ݭc�޿�K�n��d��D��i�����}�8�(�4?I�z}��������	������њ]b�
+<(��3�9�HM`�q�f9E�����ݏ�ݻI��$t)��Pa׈��|G/M��(��.F���4+?��4�>>�pnd�a|������1D�pr8�ay���l����!���NG?,g�����.`���(����G������,��������#��l�c~��G���?�G����sFx����e�i��<�?��Ӭ����4ͽ��4�s#��Y:�|�&6s��4�����9O�M�@�y�'ڋ-��4��H�hv�!����0�w;�)�=����N����M~o[��wS��-`%�Cb�����0V3"�i�S��+кSn쨓3�s4	t<Fr�ep�f����t�����ޱ'��a�&��uY2r���6�͓Q��4�'~٦�rn�6�/�	n3�e]��NY�莌
��D�3$�z�?�?�=G�;��_�|�����k�Я����	�B�W����"���1����Ԯf����U�h�}#U�oU�7{�!͈щ�r�py\�D��Ԡ?���ȝ��&"����v�����v�͟=���{|�ĉ����k����z�
aAm�>�+�f���L��K?'r���O�37�,��/��ќ�n������~�i݉�I��f�r>����o�=����E�e*���(%;}G�2�3�y��B�&���y~D��(N�y�z)<��L�]�5��HY��▋���n��N���g(��D���v�p�O�5��n~����q���g����j��.�)��v��h���ʇ��m/��&���d
޷��wM��>C:���(D�l͝/��^477�c���0��ڴ�}����DE�s�
Ir@�s�3�O�ÙI�c��m�r(�EQ�����x����������Mk��-�)�2���)W�}���p�+/����(x*
l�����ٯPw���%?��<�S��������t�������}��'� �7<�+���W�N����M�!'G��Ķ��^E��B��m����a���E��ўI��#\���d�z���G�G�5tK��=�\��>
�>s�:�; p���X�����^#>FD��q�ώ >᥂��Bގd'��r���������T~� �O$�:H|� �S��6H|� �i���$>}���A�s�_8H|� �Ńė�|���"�Hhd����ۋ{f4A��>���z~�DM�E;@�rH�>`�H�q������%lz?l��w>&a���l,j�Z7o��81j;|�&�?JB�`���1f>m�y��4j��i=�;?�s�pv����Gy>�;��M��h�����=Tzl�aKy��K]D�V06�Fyݐӑ�ˌ��o}���o��3����/eJ W��Q�jZ.з���2B�F�?�?�>I��$�+^_©������ߤ�};���G��B��a�'bN�(��m!G�!�����X�s�F֠�%K�����=�Jx�0s�_�K�Њ�V�i�|l���t	w�@�u�R^�O�������>���8�������bK���C�/�>�=����ɛ�������?�<n�A;Δ���t�zX��ۗ�{Z q�1�_���_7ʑh��
`��}�b}o��D�}H�&X@�܁���Cq�7���Q�������@q\�%>�.,�J���;#VC�'��Y�+mL�D�~⢪�@i어Ĺ��&���RvE�g���}�-�I	�-�c���0J0=7���y�k�ŖQ��e�Ί�g�,���	?���c��-�=Ұ��X�:���}±ʿli�g����;�L�~9�R��Q0��0�'���H�␴d�m���
�Nnn>>H;�t������CpZ�x�)n����ފ(ɖض.��o/Hh�/jN���	��ׅV�L�_~��2j��7ԿD��I����?���3:0���[�%�Y|��P����Y�?���֧�l�\�~���@�<�\�-��>Aw[,2�?������~[��ov<x�(�?)6���e�b���AG>l�h�4�{$4����m	�s�q����ؤ�e����Լ;N������}�~Ҩ@v<�V��q�]��?!Y8��$Ǣ׉@r�x0N闟\���ܰ�����`Īv����;wQ����c�]�㹋��{1�#g^0���;~Kn�ة��Z,���c�M�w�K���S��ɻ�"0�o_�Q��_��ZN1����C��$��'�BǾ���/�=�������0Ɨ�j:g�mk�(��/ˆx� ��8�>�Qb�z3�}��Ę�8��� �A#��1�yb��ˏ�w%<ѕ����/��h�WE��ޟ��?W��_G迥�z�@��!}�Y�r��5��6���YRDe��;�{��cv�X�>���$<z�K�7'l��F_�j;�?S�R���{q�&�ׅ�S=徿e�}����	���'?�Xa��RwH?Vz��m�x*6�}P���QLB;=����2����I�]�qgGy�<�Ϗ,߅|�h����}�|��`g�
y�|֎�+r��Rh��*E�)��U}��OT�I�>p'�����)O�Ve�)����Tz��J��3}�a�ZaAZ�
An��Qz����N��3��G�r,W]wΈ?w�@�~�ja�Q�OM�tū��%[
�������J[��O�N���L(YR�_��?�bE���QUIK�����yk<�ϫ�$ͫ�����3� R7�@ &P{�՘�9`�G�q�?3�pf\E|��8�@p~N����eb���1���DR��ţ*���1D��Ԯ��'��}ii�tM���ʢ|}�����\��{�U��b��a������&$�1p��W̎� �{���{�E�w=`����$�(R��O��s�G���R�g"Bߤ���U؉ЁЂ�q��g�����oB�d|�g'�6|�,;	��ɏ��Z�!�A8����D��t�͍��km���N���zQ�J�U�իI�M���BʧPBB�y���/T�aBB/���3e��l��3P�,�a&����8aT���$>�3��)H��6 �|�x?�����}�o'zT�߻���U*M�
}?����&����gB'�N�.�{7>{6��B�T�A|�� ��>�::v�߻��6?_�:`�|aǝ2�D<n[�4)�,�����b�;L������⢤�Ӎ$�������ߜ�^����UDI�>@���x����ߜ�̵��Yg�4[�1���V��j�[�nO���a�s���cu�kqT{(Ke�T��L��U64:j��:���wX����kKs���pYk]�M��5.����ꩬj������o��7y�k��Z��u�X�6x�Q����\#[R��B�JW�����X�k���-kc3bo�Hl�t*_�ߋ�
DEՍ�nw�]7Fj���zPb(s��T������JOj�Q[�zh���Q��D��lڍ�v@���X�h��=.o���r��n�W��T�^�޺������8�͂xbPŸ� qnu�{��J����4�<�s=*��(��F�(���5-��P��6�MVU��TV�[��.�â�� ��QY#
�R�쪛Q��f��k��V����Bkf4V:�f�h0�N]DuOY��(�t�a�j�5։�����Y����b�����0��5Ճ��'*�{}SUscQeSԬ��:aDo�]�d���+�?_��������T�*��K����]�J�����9���M��f��JW��F��p�W�7�Y�X7¼e4��ֺ���o�ˆ[�[w0@~L`[vcsԪ��������7z��]g����e�p���A���7��ǫ��7��ɢ�m^�.�t{r]��h,:�,Sb���\�u�C��I�ϱ���zg,*�/ǧ�d�!��oP��;�OJ�OO��!*�kK.7P
;�����0(�� �r��.є�����F�Ѩ�9��{qc�S����l� ]nI��۬��-B��w8���uS� ]�0�Y���~r���kF~���dP�m�^�T�H�Mv�2'Y�v�ilnAk4x�a�͕5Բ�n�m"y�c֠���˝����F��1��<��Z������6��T׷`JW���q�V���Ty�d����M�[no�m����׸n��ao�oݙ�o�d���m�?ߚ[�'���`�s��y���.�6�L�j�;�v��mw4�N��X������z�5%blK0��4Fuh�f�C+"�G7����26��1�nwe��:�lq�⩚��%^̔&G���4
ڙ�(�1+Rh\�5�B1<.7��D+��0n(���0����j��-+#y@=ЦL]��`~y0�ի�\���[A��s50����vh�h�ܮ�gmhם�|C�6��(Cً4���j���ka�q�L��˲���e�D�7��V�bM��osY��A�:�����iي)���*	�,9�'���l�bK57}S���1��y��{���Z���<%�����t"�J�J~W�V�d�Q<��VR�G�ܦU��6�1��g�����i��M����D�'��+�+G�_U��K&�C(��"WM��ۤ�Y��P-�Y�~Z�~j@��uJ�3���?��4�$��RS�7��qY55X:���I͵�f=bJ~>g�`�s5iF3�L����^5��[s:��"��c�k�5���E!�����YQg.�ycs��1�=H�)$a�' h�ja~�"�D�c�A1���4��ьu�Ɩ%���Т7X��pZ�A�3_3�4�Q���t�[�Z��q�X3s5f�j�՘]��v�j�iav�f�̴��&l�'���Anݮ�Q[�URt��hq�5'�dY~������E+��R��b�N�G����J��rL������.-�ߩ����s��]�0a&B6B	B��>��!|>�����#�Bx!�~��0a&B6B	B��!���7�������������� �|@�6�3�J�\!<�����#�Bx!�e LD��*��V�%��R�]�|�1�g^@؏p��;1P�D���%U.��Cxf�,�|��`��8��Bx!f#�B��Q��o&~�F(A�Bp�t��c� ����8�)�wb�P6�D���%m�����U����8���@;���Axa?�q�S� �<�!LD����P�P��Bx�1�g^@؏p��;1ɺ.��D��
g���6U��\�|�1�g^@؏p������P>�D���Rh��Y$XlѺ�,Z'Bw�Ek�g>+�}wX�G�ߩ��;K,��%(�bIh��KT��3�`*�姠V|���n|O)2�o[<����N��d�m�QBB7B�	k+�q�
�3a*G���*V{[����({΢��%Fǣd;t,��kW��"?]ǣ��;u<F|�8w�=w��Ǌ�y�m-٫�K���:g���/���X�L��l�� N��t<N|No����ˣc��nO���e����J�>����~_->�q�,/���=A|�����>a�L�:�^[շ��,(���*����o��s�Vo��KYy�/�Mت�����X�-��B���T3�g�=,������aE����9��7񹓥�{�������+�����)=�O�6�)��M:�\��.g����)5>��'Y���w���c	�T�V����7��Ʉ���0^�z$�����Ԟ˜���ڿ����O�5\�-^�E�Ng�Xe
Â���l3�*�.���N��tJ��u��g2��:V�g�w��?|�)������@�g�O�0�	\������w���M���������g�μ�3L�m63|��g�౬��D_V�o�O���"����>�w0�&~�`��i���O3�w|-��Q?��6�E�_10����x3L���0���i��~8��������Ͱ������{&~����ğg���_5��Ƕ�Z��o��'�1<x!�Ӂ�wxp������������>�P� '��� '����֯�N���� ���w}X�W�h���-3ɟf���|}�įO2܂���aoL����Ɠ�o�u��	�',��&t3��g�� �.�O���3��f� ��w��gx�t�_�1L��K>D��0ݶx�ǁ70Lށ>�����09�����0ݚ�K��I�e����0��=��z��_�0�ߺ��k�ob�|��3|�<����|�gW0L�k<���a���Ë��b�n��6�K���Ề_d�܉���z������ �1|��{�|ß��ᇁ�3��R���1�e������o�3�����n�6�������0���`��2�?�{�G��pp���o '1|x�� �`�<�\�?^�pl,=S6������H^��ncx�#O����o3<x�i�����ӫX�3���7�gY|	�y���r�������*�9� �1�8��V�o^�p xÏ����73�I���7��b�������_dx/�!� ������2�K�S�~��?�<����`���^���w�2���[��Nd8����	���
�.��Nf8����7�`x&p#��S�>[g���1\D�.���]����U���^ǰx��b`�>����m��d��,���G�O0z>|�ᧁSV�k�5����<��,~�1��0Ç���~��g� .`����S�F�	�$�}��`�}`+�#�&o���${���q�m_���u�;������ ���l����u��Y��/ �a����R�
�WP{�SvP�^M�g�^��k��c����3���ϰ������?A�g�)j?�_��3�j?�ߡ�3�=j?�?��៌ւ�Ⱦ~ل�b´�;�����]A~�B�_���c����G���	��L{���F�5s�;^
L����x'�_����
����T�L{�z�_�;X|?p7��e
-Z��3���%
�.�h�
;�i��f�7Ӟ�4���f�y*���0����Y�6�Ǐ��޻�3�iO^���r�^Ǜ��g:�L�t��
����pm��x�š�U<�\�K�����&�5�M&���r�;Q��`�����m�.��n� �>�U�cT�
�6I�_���O���bM�ӿ��c0���8��O\��o�O�$4�LS�ہ�.���ݦ��/�Ԯ��.S}�?�����e��=o.�����1p>�G�m�8���Y{�~o��y�76��������!>t��fª>�����Z�+�h�2��ۥ�z��/R�����]9J�o��V�'(��&����;/�h���K/B�ؚh�z�M�]�	�
������k�5�9e���������S��{��9T��Ry�ܭ0=��i5ʋ�̳hw��I�}-�I���� .���=����\)��� ?������}~�4��ρ?d�8���`+����&�)�7.�-�������oOx��*�����x/+�܇�|��$!��_ ��w�M*�E�����;���'K�G#�֟k�;s,�3*~p��5m�·��b�OS�1��.�O��p ����I�+�B����_��"�����ho��7�~̏D��*�}|�e���.��}Jp����H�x�߯�g w��bT�
��g��xV��q��#��`+�+T���B���*�_��Ңթ�O����'c�?�����K0�]�_	*�T�L��]��<���*�.f�/�xk<��	x
�W+�_dԷ�r�y�8-^{��Đ?����}V��%�4�/��>��
�����l���ac�����7w~_�>��]J�E����?*}p2�7�=���T��(�Jc~|��oZp~uw�CӲ>���� ��ysL�O �a�7og�\�KM�c�L��= �6� n�nW�s[�ڀ{Xy[M�w �����������o<�7j�6�J�'�E���8�n���w,0�+8���B�!�F���+C�gp�J����p#pO��=��V*�3
xg�&��~��/0��x6�P�nM����p:k�hL�.������~Ӂ;�8�x�D�뀻�-��=�<���t�;����ST��}�'�b��)�k�3�.V��$��y��X�s��ي5�N_�n6�6 g�7��SW���3�})�w*�AO��2p1��-*����W`���,0�:!�rU�X����W&��781��6�
��	�g��N���D|�ր/`�7T���3f��a`+��f��Q�CF�J|x9k�k�]l<c�A}h���ӑ���tJp�ඟ�np=�ϣ�^l}\�)����l��O�~O(~�p�4�v����54���U���Z��)�C��k�E�� |&N"��5�'[��7)����"�Rz&���;0޺<}�;բ��~���x�%�#M<���W�S>e��7p1꟦ʻ�e�9�w1�x
�wW�ݰ/|�ŐG�
(�@�g�{ �oU�e���>>�������3�?
O��$s�1^���2�.(�޶�`�ߩp-n�3��;�6�o>h؛�N�m��<;�B��o�b6>�@P��3ڗ
��������k�[>��s%�^,���+������jا�W�P���'�\Z���F{��a��F�7}����p��F�>���g�0���`�{����?\���?�ێ����&��߿6�?�݀��5-�On�d���~�i7��ˁ����܆�����7���_��(�������ی�E�6وONf��<��<��Ɇ<���Ƨ�z�Q���- F���w�e��wBߦ�Q*�Q�o�{>o諿X��u� e�.�zu��_m���B|&�o�݈��G(	����8�����Ģ���.~Ř�� �����7���5�ؓ�*� �6V���1�p#�����]1�}�I�w-�����]���T���?Q�[����o��U��pq�%8]�}�=�)���.�c�<�x�/��}�&p
���
����ژ��X����h�D}�A����� ?��o�f����yEi�]����ӴGu�w�Ҵ/+�k��k��/����E5�q|r���#|��_���0z�ܵU���}L�}��&?.��$��X���p?���a�]?�n2쵹������+�;��wC�Ԫ�>O_R����|	x����5���C���pf�1��H��[��TyI0,�b���B24>e������f�=���瀗s���S�Z�S*�K�O���O�3�Yz�H�1��w3�y%pK�
����������I�	����~l�_N����owf�?�d(��������^�X$�w�}l�d̷��S���	�X�Ӏ�2�	ܕe��U�=?7������d;ͷ2�^�oZ_lC�N�1L��8ߠҟ >��π��xx�4�Te,�T�L�Ӂ;vjZ��o��X���*��,�C�}������ۮ7��{�?ḑ��;���j��S0��sT�4�&�>�Շ1S��x�E����MdX��h�uzw��}U�T>ۯ;l�e�s,&R�?��|�nU�m�)�߭*���C�g�g�����v�d�c������B~�T�������������y԰׻�31y)�
����_�J��ўS��l�> ��e��'A�f��W\������c�z�jZh(�Q�>pk���=��ƷM�ww1��*�6�=�>���/�º�ZC_��`�-6���Z����=���� p�:��/�ͱh�U�/���W��.���OI��/�w�����o�$sj�s}�w��	 Oc���;|�����������z�i�ޱ3п�A'��������
gw�3�x'����B��$�Y��.f�}a��W���ۍ���Q�_�	��Cy�J��$�����N�����3��m�c�m����|��ѫ����o�������1|��c�5F�wy*�g�}p׍��C!p�r�6[�Ww�����k�;��փ��l���T�>��?Q�bj(��B��~�N�� lDU���P%^���n֪]���n�b����ӫ�WsM��r���n���<M���%����2�('�.��d�ڳs����X|M��������^�iv���uZusSK��㨙>;%5U�{C�:B��ZWe��^�mjZ�5�7����Y��6���BR5[KK��3��l��Ffi�cr!tRA@��a�����^�v����ٷ��YT�DxB:BB*5��jM*�M�ĩ�z&%�I�fQ�Y�n��E�fQ�Y�*r%�E��(q%�Ii�#m��7������$�-j�"R)e*�JE̤"f�"(��s����C͜Cm�#zE̡�P�#�r�S�tʑN9�)G��ڢ�|9
��F�m�ٖ!�J�X��+�IP�&Hc�	
�D�m��6�r�h�M��&o�)��yg�\3E	�:6Ad���M��&�l��	J�fIy�m��6As� �MP�&�n$����i"o��3�7M�My�D��"��lɖ"�l�w��+x�6[�-��yoyoyoyoyoyoyoyoyoyoyŸ������������������y���� �����������E�t�2]��i2D�"M�H�!��P#.�<E�v��9�)r�SdJ��/K(�P� y U��T9�r�S�P��zf)N�H�H���*�'u��U�A&Q<��Sqm�� EV�"+O�4�,.re��e�fH����R��&��Rq�P�}���R%ϥJL�ܘ*Y05M�YJ�� �ܘ*�1Urb�`�4��Yb��R�_!|���7+C
!������I$���0MJ є4ђ4т4р4Q��R�`�4��i���n���rç	�O�&>M0|����
���r�tR�'�]�Qe�)S�d���Y��I^�-@��ee���S�?ӟ5TpM��n'w��:0|���k��f�k+�]��w���uN�i�ܡI��S����d�ni�&�=�cT#؏�Q�V�rD���?`�#7B�	
��|��J�~���vF�!�r�D�F�Jo��
%��ts��-7'�DPJ2S�U�nYC0�м`��j�.9��[��M�-��U'������7@.�C*��k����<Ģ]�/����Z��A�����\mw7�� �B��w�3G[�r��҉o-��Kj����&�a�jr9�m�x�����͊�)���Q�P�édR�dc�@���.����47��<��4����~T�=��nll���]gX�E9�4�v���j׿F{�a��<N�D}L�n�K�i�Ҳ��2��ݼN�3��΢,[nv�;�^�ଡ�˚m�wGJWћJ��5�fW��娉��DUAC��ҵ>Rt����e�V�X �8�����+�-uy�B2���qI�9S���E*��hJ��#��3�PH`ӗ6� p��VW��ñ^���0Ӗ9�Ų�K����wb�RT��P�
�Me�-@�U��\8�c��"��1� kv)d�sT���U��x'f�t���R[*���7k�wV�5�9�Z�g���<�FR<
����r�*��6:ȑ�[�w6x�Ug��hl$�V�$c�k�UM-Z�O�HM!�#U�۳�VRsc��VM\h+k��@���tx)z�����o�/���P��Z�r@N��E_(�B���j��%d\�q�
1'�½�̮�:LNeQ����'M�Hn3�t�& q�l}pbɑV�
֯���p����:�^�&���Ro�r�h�e_h��Mn��P���`��Bb�O9����J��c���H/�l��)S��3��郋���7{q�b[nNyI�� �莬�����\{41ܼơU�k�I]��MR�c��,eG�(6 ��Pj�ՠt)+��E#9���q��@���~�K�UZ�ti�����UGM�ta�$�AUS��-sT�^ �r��6�$�8���\P"����4ֲZZ.��uB��z���.��5wC]��2A0�^��B%O�t�+�����D�H�R�H�^+mA��k����
���Js�t+wV�F	���9�[˚j�R�ZgY�3�KY5�-HW����lm���1s����C�!5�<6A��4�q��]�On��L��N�K$=�'�5� �[$��u�"�1'��XQ1�j8v4��t��V�c	��� C{q�=u�4�tr	�@��P|ѝ�F�R���`��fg���
��UމyU���3�I=PYS���.�U76���Z�nQ��IU��J�(�\��ulF��+�,"Gc�2��lr���^	Q��UV�RG��=,
�����i��1����`LGީ���a��.���CM5���:T� �Ҙ�P]����~*sU�HG��56c4�L#]5��'�U�P�<�$e�ؚ�ΈӸ��XT�c�,�Pq]���%��F��pKy��&����Yy��!:��?���P()�ӱ6T���K�8f�T?���MQ}UW�X[$Ԍ��ou�:Q��ްE�g�A)WZQ�R?B�g{kk.[eKeu�'"y��AGue"sj�mH�l5�uS״�}� f	]D�p7�*Y����Ql��WM�*TZ<���Z�.�����Άu�G����/Zc/QSH�aW�ա
'���~�$S{R|��}�c�������v��_0G���[��9r;�F�μf����Ќa$�?�j�e��9��*js7�U}Pf���^t��Mc���/�������l��)"EЀ�$ȝhXa�:9�+[Z�D%[2��W5D��RNZ	����	SQM���WF\Z��mFQA���ܵ�v�Z�JY(,=��	{Ί���|��/
�]݁�$84��ahl;¦�2����^��8bR���yl���뤹9�b�[�f?�&�4[���HR�ɭњܹFNy�D5߈��g�9����;�Y�Ć��W���{Rr#'D��iP�4U6D4Hy�Y.i�����]�2,���_6��s���yǂ�)��&�kŹ/Y{~�b]�3ȲL�PbV�L$�V\NB��D��Od�h��0�$8h"���o���n�A,�]v7B�4�\5Q�U�RƵ��0����JsI	��l�;$Ҋ�|�C��4����g�8ܞf�C_�DFYfa�/c�3"!���0��U����La�VдS�l`����C/���!����4o�E�C���@����Ą@�c�De;]�h�}��,	`��潮Ѓ�m=/�;j�}?U]va���������b�ځ�84m#�&B�D�=!&�PwDؓV[�Ѥ�d�4�q�,t�T�gA�G&��y=�^8�[�)�/W���	7���C��!�H>+�u�NS���/�)㠏����C�A+��E�á��h׳�f��HSX^#VB�ꏧ®��i����P�U�o�rE�B	�s$�z�I��au�v%-�\�ً��+�}bٺ�&["��-!C�xSjP~��O���-��Z�N�jI)����ϴuGzn���	�Gj�&�X
�:=X��ض����~���3j�-�@T@f�݊z" lc�aRO~L�m(gb�����r9��%����
{�d���&*���vf����6�I���r�E�Q����7O}�̣�*�pEޙ�`���C�3�O��CT$;����
�����ك�H��4F4�+{.|f@��_IB�0ƀ�C�'�u��¶HKX]\�<�1Ժ�52�i���B#T"�zb)��L�V����5:�A�U����]Q���A_�{�E�0�6�m�)�ʧZӦϞ>Sk���Z�\�9�їW��I�O��m���ւ�jknM��:{zj�-��gΚ��i�k�;+��8��Ws��ƥM��t�k�Kˋ�����=�z\*V(� 2���j���\M'���4�G�<c�����%���9դNO��AX��Љ�f��z�N �ȏU�hnXd:䩬Ҩ(�Y��Mw׫�����סw�轲]*dZ4Mw_I���UZJG��P`.邾��5��T:���_��qd:
�.����fJB��P ��To�JC��kw����~
}��t���*л��Z=ݻC�[�=�s�<��T�t�Z}�{��*��C�Q���8z�m�����1ڠ���z��*��C�7!�<��G�#��t���2]<K�����P16t<�.�,�C���t�2>�������7����F��cN��f��F�ác�>O�t35y��U����gY:����#̇�E��Oz���R`�s�w
T:��E�v^Z/�#,�k|n����4�q���{���BV�U}����G��-��QޟX:�'�H�to�~ ]����wF�|C��ޠ��l1��4"���	���%}un�|u^���k�[�_�w�,�}OQp���N.OGa�%���F�+,�����PK
    +Q�H삖=��   8   org/bridj/lib/win32/bridj.dll   8     ��      �`�� �w��� hT��h��1�Q9�����b<�/�;�J$��Ͳ��
�|Dk����[��"�$�H5ԨQ�N�TSM!J�ｙ�_��?����ݽ�y��7o޼73��e�� I��@@��J�/K�����/�vx}�^�����s��@ꊕ�ݱ��{Ro���{�s����ԕ�{S�75�湩�ܷ���II��w�\�������(_�3���/]�|�}�����3[	��L\�xa�?��m��k�y���5���\�/�f�]�f���j�\-�Yҏ� I��$i3O���,p��I��%)Q�ѮR���7dB�1KG�,���K�;:��(IZ��NO��ݺB]���X%iŋ:)�m�:'��'�&�o_��ݿ�$��H�T�}��巺o���n����"g���Lr�b
� .�u��M\�����7�
<#�t��;����} ��e@̧t�ˎ'������
Զ�j7��<�z�N�����I�g���b��ry삁f�� ����mp��:$�.���&5wR��l�Ht�Լ�|Q��J�
�{��T��&�a�c�a��'O��Ks�Aի��P�
ThB����H��?�$��M�2�@l�k�F�!�g]Yo�,��Nɲ�
���6�-,����-W�;3^uz��˷c�r;S�V��̆f���Eu4C-�^{��Db�ұ��hT��l�2�Xko����.� ����5�g(��#�Ѽ'�oS�������M�7���<��x���߿�^O���5*�SЀ��ܔ<�0A.$K
Av��{�\�$��@�ܢQ�������gC��x�5:�/��a&�ۗ+IXゥK�E��'��*�;�U�=���2����<B*c�g�-�q�:U{��72�O6�)�.QP���.�B]Z�RW���'�&���t@k���@1��<vC2ig���i�+b������/�����������<��/=��ϣ.g���;���dثY��m��؀6 �ꞻ��5J��)uk��x��R"y����jj����i��4( l֦|6*��ck�Dj4��M�vn�g�J�Ӏ��������	�Լ�|�^bD�؛�,���%���ٍN/�,s<W0�o]���>g�R��]�Z������|���JM���bG�\�%y�]����b�\c �3|��@��p�u�R�)�vJ�!��Q�v��:���On����%Q��Z�.���a��$�X���<� Vd'�T��	܊�a�Y��%�+�!�v�0U�V@7S�vʭ:"�K>`P
��Ӄ�'���k��j�:��|�019�PLA��}Z��˥�g�+���V=���Zth�f�m�N���St��CChh3��0U�2ly$J#���X�A������s�/Mh��4���pa��4CG��_Ќ4�Ag��_����_����I�_����B�_�z�/����B�D��	�@3i�f�H����t��2��=��V��P��D;XCC�g���o�wn���o��>�G��/�1V׭=�N�K{�o�>�	�O�޼���[���V��	�KM����"HF��:���Bn��-p�B�=F1M�P��ͮ���5\<U���I+�����d�6 �`j�	�C���K�%]�{� Nʀ�Ľ�h��mV�w���= ~���'?hѯ�j�Ws��G�R����ٔ�6��Z{;o���e�,�
2�9��Ac�ŇP�TQC(�H6��Y��֒�����m6�$�2f�
&K�X�����0,�q�DrI0J�!��N�N��*���P��`;����M ����N���=�u��6!�n�y���7����_U?EO]��s��� pT]#�<�+͡0��NU��'6�i�ܹ�@���#��6m����މ�O[ ��zj�`��?���j�'c�<�3|��S!�R�~Z�<�܃����_)<�|VL�����NȔ�wj���X�S�tUt*<K�T�̍!�6H���+�O�g�@}@�ӟ"��H��iN��n4�q�N�uX~ߐ��Q�v��!���v���q�a}��5qSW�!�ʂO�	��.2vm6z,���k�5(h) ��r#���a���P3e��|�En����~78�)nD��O�p�k�I���Qq4��UG����f�^�F����:����!���ސ�,��d��u
�lޓ7>�F�ȼ7��p�����6�j���X�mv�T���!l�.�*���"31�����OG}�#�a1{G$` ׁ.�i��h�J-hS
a��@7ʥ��O���j�y�Hj�5Nr؜�/�kWҘBf��+B���uX�_�9���=7K�����[o�����B�qs��"���}S0A-`����	" Zp�a9X����B-��& ��8��G��#��V�o��N����w�����mՑiw�r���R�s��h0ef������`fCM'S�H�e���+tB�&��� A�_I����\j��B��)��so�?e����PР@4�UW�2i҂'���+�U�@ݯ��\Z�s���}��\�r�SK�y���\-������s��|�@T8�5:����J�>��i�pW��Ar*y ԛ������!�qC�Ц�%�
}-���-
om�B��S��.�`���ޏj���a'��|�r U���8~��� ���8��x���q��Pfi*�"|D���߭��z�@ǥ�ɊRq�+��e��{|`h�_�k=�@��8Z�Җ!�>O=�%����b���$��I������唋�E�)y��	�#�f+��%�Y��ZV��5'<�`�ɑ������3����YJ�Sh0�7�ח��	@סLBׁ�X#�,�FQ᭠70��������k�b�Z��b����Fԡ�4�>��&m��f�&Q�B�<�U���G׉t��Q�6b���$�z)�R�[���$3�-C��s^Xz+,����!+A3�T�gV.���q��D��s��&����@�	�)F�A�Gs���˥6��Ա?ٳN�=�u���������mz��Z?�s��������$�&k��LH�m_���`F�@o3��0��g�z����\��&�{,��+������<��T��9����baz0��-���b�F���m�B�X#!�����#�daf6��"ɒ���4�Rt�dy��!�B�_�j8^��Z8^��q8��������B�&�8)�6�\�Q�Mq�����@��\-H�d�pC�u�æ8�D�v�m O���D(�Π�<���۰	a�9��h�:"N=�|�l¤��/ܢ�N��N)���L;�EO&�>A��aw�ozs[�,�S��W���T�M ���*�B��xm����'�����d��-�KAd��u�i(-�%�60G �6�G�\*d���`�Sp����ʧ?~L�i��U�� �v��b<|$$* ��(��CN��?4,-��ٺ�$ܤ7�A��&��ץ�teC(�,Ok�8��
��[��#x��V�Ҁ�p�5�k�%Qc���3�P�F�,2��{�k����h}t�C�S羈ܣ/rDmp��
|}�F:.;5(�Rp0$G�V��7�4cmU|����5�
B�Oc䗼��/�tI`�V�>�`o׷��vݫ:�j���#����T8�ς�Tn�����c'7��i��.�`�j�f�sA�.�Ο��.�]C��9vC�.���p�>�hZ��i����џ*��9��{���s��UC8�j����ڬ:6s�*��R�M�o'5�v9����FBƜ {� �I�������sI�d�*����c#��M8�`�\u��;���',��m�|n�5^<sF�qa(k��lY����*jL�}6��G8��]����/䑢z�R����`6g|�Q�.��Ԃ(P- R4�,�A�R���'�������t��g�����<�����1ʱUV�G��x���ӭ�ܻ7i��D��F [�_��Y����.D�����)'+�Nn3b4Ʃ��M���x&�r��/��։��`$�!��e[M�e�h�eXMOC���C����2��}�&R�{��]��ko/й�Ą�2ҞeB��l�`>�\-����{�J0|,�'M��� ����v2UK��fɍ\�/�b䐣�
�ҹ����=��0������%�g�$Z���[/�_
�r��?����k���2e�is5_ BGK��Zw&B�_�(��PD^CRǕ�[�H'=�;���'I=]cߋ��"�����B^�I̋����� u ����1摷�����2h��L#4i|e� ��&8�� '	�S���/5�\۞��aPh�{�k�� 1��
�[l*Yz�P�\�?W32"���*fCzm�S�oV�7NB�Ջ�L/�����mq��ox �1S*rH9�hr�$���u�	D����-9��c�6�e��$m�����,@V����9Q.g_���i��vU\_S���"#⡧��ҰlvGf�GP��|�'|�sķZ�����,���w��u÷E�H��3�v��e�,���(�[�/d�G��~/�-��p%� pqy��q���6�����#��9�oJ���^y�8�ǚg�*�)�,�7%.�i�L�fLDO����ZWe�R;>$�Ѝ[
�{-z��ٍ��E������0���Z}�j���s�@[	�u	���©�?N�,/_*Yޟ Yp�O�,k�����%�r~�~?�|8j�r�dy��r�����$Ϳ��3){�ҽC�?ݓ�Fp/�z�fH���u��r4��춏h�Pf��<Kk5�����P��B#
m�,�x��O�X��P�Eδ�YY�ݙZ���K�(qqd����J�2���%��U����5�%*y[��yD)od��4�3�w+��ax�BC��^*va�N?��M���N�'��A���&���g�Qנ�o�uk$�v�>�_�<����.���k�� ��Hdm��Dm�/�V�&�²[pN����b�����"�d���dg&$����pƝȥa�~���ķ<��t��A�ۨ4e���3��8פ�4��C?UCOq�V�>��DW�M��F��DrP�;���B���ם��*�FT\���F�/�[
��Oh���q���)E����w�eE��er�MD{I�!�O�"hn�!���N|?�yҠt�ԇ3�v_�|#��X�.��ʱ�#�Ǖ��1V�v�;��}�}��Og����a���Ҭ�>k��fMw����lpO���������fhf�X���+♡�m�:m�X���z%�Ǣx>~/L<�K( #�������#J$��5O�L�6Md����.���eLJ΄�e�d�:U���&Yހ��z�$K=wL��S�{
\�8e�a���_�>dS�b*��rM��s��T����?�[���>�v�޹Z����U���m���J����z�^�~>ͤ�ȥV�=׌s�p����yG�����+�o�R��������*r�)l2��A�K����Z�8:Ԃ�̂�F����G���P�6;E����Ԯm[���Ө�mDY�>W՚�z؈"�3`���8�)|�Q��7���/i�+	y<���ƾ�7m�wVm滠6E�"��v�����9����]��\�{��N�ώx�q	���F�������ݽ2������������?�����G����b��;~�F�7Ā����8=M��Ƹ�����wv��nb�2uT�x-=W��qz������;����	���;��g��;~���r�[�ŎC�]kw��TWf�f� �r�o��rmB�T�=\G	�m16I�y��â78�����T�-Vi�����U���L��:$�3L|�`D^��V��E���:�n4m?�m���5H:i�cĖ1\�����%uQ�$�i��Al;��v�Wu�F�L�mJ�2����o6��ƚ�?A�i}N���d��0Tj�F�T�t��m�MO�ko;J��7 �$a���oG���0W��k�T��4���B���}p��A����h�]+�։#����c������&��Au��]'b�]q��q��Cl��M���!�U�P����N{\�q�ı�eH��NU�b׉ÆˊP��X��u�x䚜�NM\9�-�\D�8���!�����ΝԞq��M��ʱ�ݱ��G�P;��ݱ��K��N�'b;�u�b�YG�P-T�/v�8����։�.i86*���Ʈ����҇c�Gc�YO�9<^�8��r�l��1v�8���#���l�]'���q���͵�m�:[b׉ÛkB�:[b׉c�k_�:۩�[���N�\��Iu�Ǯ��jD�:��DZF�3�l��x']��Vj���[�Q�vw�Jq��lv=�Mj��:�|{#�U"�F8U�S��6#�ND���!�6�C�N��U'�ߎ���`C�g���fj��j�����`.K��]'n�w�A�MX�%�u �6��Mu�����Kdb� �y4�l;[=�1��hl>���,#{��봍�����̢��F�`�p�������m7!����th�l��`��->v�r!�ڑ1d���VH�g���(*g������M���Qy�(ϴ�nQ>�<Ԕ�z.���/�s��'��eX����˨�2Q~�V��5^�(�o��r*�\�o����Ǐ��yT��]T�%����/ʗc�'{)7��[�ߡ��,�3,��K�*�"�K)�Gx���?���T>U�����-�o��O�R>�ʧ��;��nQ�˷�R~<���?Z�_��>���=�O����|�|�a^~���K�IT~�(����廰�4����dQ�6F�_��?�i/�R����K+?Y�����t*?]�ߥ������z)�C�sD�N��nQ~�X�c{.�K�s��;V�_�_���z)�E峴����,��c��^�Ϧ�5�����7mnj��T�)�OO����b��^�ϧ��5�k�ݼ|��JuriX�5�XV�z�|(*~d����w6�kU�)�L8A��O ���3�v|:9��������x�ӫ���܌����	*3ĵ9Up3���l�|=Q�T�n�8�;�i�5��5�$>�E��4�P�����S�_2��&{^g�t��^Tk�I�y���{��+�38\(�M� b�cf�G�?���jr�G�ӕ��W˗r튚^�|W4����Qh�<���EN���Q؟q���[���Ӧ��y�C���j�u�q؅ꔂ��}'=�Cu��0��ෲ}�������3Ț`ߡ؟U�ҲwK>{Ѣmv��u�>�p�����q�k�8t��ҶX���!���}X�iϬ���*��A�7�'qE��V�Ԃ�̂f��eZ��M�-y�o�cՂ���z�s�g��8HE����Z��Z�����m|(���j�j�gbY���k�<]e��1թ�����I}Y��%��Z�F��8�|2�86���J��R�$�.��uu@��<��>Zo����z"���t�q|�?Y'��ߡ��p%�`���#�p��$H�ƻ�/L�מ����NW�����D��s>�p��
�UE�[�~W�N�Wl��ʾ��Spӕ/����3����ʩ�9��؊�,{��]�������q���Z* ��6A��1�+֊݆k��v���D�-�{�	]D�m#��]��;�<{7e�f�ݱ�}��//J
<�?�ޕv>�����a]�0�J��z�7�'�{;�_���&�5���Y͞dײ��&\�n�B�j�#�@6�[���%|~�H��)��
aQx��8����^� ��=T{�C^��c?���?6���J��s$!Trd��o�G�I �T'�D<���2=g��@�>~Z"�������� ��] �d�;М�(�����¿-��G�^�N�t���]�g�-r��9ѣ۱��G~9��M0���;��;ŒqG�a���Q�`\���/��&K$W�7P0ٲK�	��2u�.��}p�XnK�~W�]����7'8نA�[B^L����5��
��'�E��J>kь/S�(w����Z"��t�����9�{x:B�DrX�@�-��󒳮�n�����)1����z�������/h�d;ف��sa����jϮ��|��)���z�I%��Ժ�	�WE=���ܟ��+����7Ơ�HA}N=d?���m�kt�
h� e�Qۚ�j:���z	��b�	m������@O��tt����z�Ot����I.m���k� Pm�����:�[�)��p��� a���ר���*��/���q�C�wp�J���$��$O�_�q1��}��/w *����?�F��6�H�ag$�D��x�chu �*�?2����	"^��4 ��*���vIkM|�{����ѥ���R���F��FqH���^.EjSX��E:d�*(H�U����Ю���w=�`W���]��w��Ǯ�� })w����\�����v&u�� �N�{��E&�I�.��.t�%��z�凹��H�ӽ"��ɴ 68�p�0�k�2���t+?��w�pX�~���'��vo�a��Z��x��54Ps;�{�l��X��s c����1������	"�2ha��-4X�Oى�SG����Sx�$��E�x�3��-��-\'�~u��!��{"���T����Ү4{�����iJ���RpR%�4� ��}>y�xY���B�88���
Ƌ�r2�N��d�LSp瑑�b���1t��2� ����\O]4=��� �6�\����^�|���y��zGA=k���ɴ�����K�N�na���6���$��$�N�����T�M8��(VzSL�p�!����G5��Z�#Dgފ�a̘c�X�)���+_3�P�}$+߿ݙ���]�9i	�L�tMHOӬNW~��p�C:12��������P�7��W4~��v�d�v�7�>I9����JIl
S�c+��(>�����o`��_PA`�����`�7W0lq�>�ןV/��J���c7)T����(^�`8�.]?��f����?�Qp��C�*��|䩒�B�4�[��5}N��T�"�����t+���4z�������q�I{��Iz�ښǚ�p<X<��I��+E`��\��7��1�]rG4g'�c�i��$�W�l�d7�I�z�ޭ&-���Ydӣ�I�{A�WMr��ݦ&���ݨ&M�%�EM�#���+�gԤ��d�&����$��R�����OM���j�ݽP��_[�,&|����Ћ������8V2��k.B�T
�};/��M�5����Xs;C[��;��1�q�Qq_ ��}�d�����M�'�V�N�	�^ɶ��E��5	���8S�;n7�?�̞��P����N���L'G�)Ӧ>X^�cm�a�𡦽N>����{:���g�#���6�o�!?oRx3m�C��>���hS�Nv��n�U��1�������ՊZwj���._����j�h�v�>�%s���54�En�5{Ki��$`����*���A;�K#�v"fvS������y�l��1��=�1VW��1��ZL�GC��mZWk졫5W9��@�x��Dռ^r?Q��68NT��oW�1ﱟ��y���AzW�c߆�]�y��nd��\�������\������<��Nt�}�IE��vF��aǱo��x<� zT��;ŉW|$ᨐ�<6���EH�?����ڣ;^�|�0��\��1b�"w�"�tDf��K)q'������[�ְ���U�������>���Z�|~����b��v"A�����v������>�Z������q9f��`w���+�cf��c��jRZ�lm��'���>V�|6�acf�S1=F�6t�68��������K��jRV/�5Ac�u�%�^J��&��%�è�n���SӢ�yv�TfNs�w|���`.�ȥ�=>yA��)�`�2���Ê�he
^kV�I��<����Ǔ��� �oz�州q`�9�pH�������y�x��N�w�kl�������bDXU��،Un��m�b���_���	���]�M�����m(� ն|6���f��Fb:�x2����q�����|�7�r��.gHh;��vn�"���Ug�m�bد��Wٯ��^�tz���qNj�%=j��m��%�u/��{9?����4V�F�� 	��{���p�f�΍a��8�p��L��4�aSF��Kvs������1�C�I��=����vM����d����K������]4gM�,Ή�9�IyOaF� 5�l����`�o���5���A��߇+�yS��f��4�r`vPx�����o:0;��௤p��4��QL�p�v	=*����D�p`�ED�e�901��-=���ԧ��;������Oq�]��'м�o�s���Nk�G���߃��+�Y�hF|(��e��KO��,R����E�Yײn�+����f����/MQK,�SN<� 5+�m	������;�����*J#�B#���WQx۰�푫(�jAK�e��'�\ޟ���Fj�Ьz�_��QWVz7v8'8�Q��3|JA3m
	2�D��ݿM�I�ÿ��}Ǣ�7�W���Y~ ~���bU_�؏��b�����s��}uNL7T�e���>�rD��t㿽7�[�5v�M�}�xhA��Y4�&��͜�::��x�k�77|�C���j12����A��}�G>�D+x�w>��������������K��_���v��[ۿ�y��ε�V�>���k�?ӗ.�"E�WY7�z��F���p��*��� k��7nm���K�Zfo<-8��1����#9��^�ԭ�,�.��bI���:�Z��]S��_S��=����̂�����8?>�n[5 ���_H⥻�hs*O\Omc�����*HW�6rtm0V:>����A�|@�﫯���v��m릭���=����\B��������?ɬ�W���.�Ӝq���x������@*�.A��K��������u=3�/Z�7����P�ܪ�u�K��A:2�mk�A5��L[y9��P�ɵϼ�h�_�I�pV|��������߷����d몛-���o}u�Q��0���"uE���?�M?�ε��-����m}Ћ��B3#V2�i�6�'���Y�����]��W=N{���=v)�J^���.e�ҹ�;\��=v[u�ͼ�1��}ˠj��?0: )�UӞ!HM��1v<�cSh���'�r$���]"v��v���ĩ���;�i;_���^t����GE��=Wݬ��+_7~�ɟý	��i���	��(�_�Uĩ��m�/�����5�%�����H�K�C{��M�]=�L��t	~
���&�_�f�&]��AGT|�4��<��1-?a�06^�0�n�^E���y<�ch��¼���rb���m�T����C�g�ɳW�1R?�m{���Z���@l���Nߧp��0�0|DR��1�uHn*}���X�����O����G��>-}�vs��_�=�� c�v|q�5�g7i�=X��C�&��f��h�N�
JG�p¾�'��K�t�vvZ��k�����D����E�o��`�#m}q*������תRf궾8�����Z��[_��Z��J��b*�UK����/�؜���[_��̈����hd�#
�ߊ�O�R*�s!���n����Op�oV��:{Ԝ&��f��{�j!���cj�|'�K�=�_�i��H�<�#����-�|@깵Gx���jw��\��~$�ܰ/�R��y�p	��Q�m_~�OAU�0t?��D�~*YM�~�аf����׌�k�M|\�m�� 7���4����7���ξ���,����Ͼ���|���7&�����cq��������u㧩7~��Q����hʆ�F#�8e����o,��M�=�z�H��\��0�Aj���5�kv�br5��Z���SO�|��DB���nHȦ��	�ug7$��z�4�ưu�H3�[��;�{�w�����-�b[�r<����Ⱥ6F�gC���g��g��c�C�]B&���� ���$k������L>��3鳠U|[�����|�	����N�����G�R���?�&�C���p�H-�B1�������ڃ��Kո���j�����_������'�
��n�t��1~�r��bnы�M���ǔ��J��X�[�F��.���ۗ��ʸ�ә�o1>e� �����O�*�O�+�u|J=7{?��c<|m0vV�oƻNݠ#Ž��<����|�h\�s��s
x�?�M^�W�{]o����x׈�.�o�����L��8�Ɋ���}ՠ������{������~��}2XL��:��<�d�=���`�$ޒ��/��.�h��Vo>�99��yQ��|��"ﾌ���EV_Ƌ���/^{�[�eߩ}z/R�2^���m����4^|������RO�=�~d�G����vG���߲s��_1-�F����!Ž�!q�^Wo(o���W������Xu؊�=�.���l]�WR�o�p0�}��}x�ḭ�����>H?�}H�}x�4n�5���?�\�=��`2�o��3k���/��������_�'ӾRy(�?������'[~���Ћ?�l�����k_\�5�/�����/���ƿ����a�R�b�=�~���ʿi��������i��X�c��������b��y*Ԫ'%H~*��cu�9�[V����>����N��v��3�|���W��}��U}�w��^D��Od@l'�{*�u�y�Z��=}���C����q�Ἶ����r���۬_��C���}��g�k��s��|�����\C��h�̼����ʸ�޾��f�̳����{�o_�f&�ӆ4)��O?գ��2c���GP��m���*����?��k��~�������_&�x��2W�_f��n�e�_��XO�eޱw�o�	�o�����'?{g��aJ���=��������CB{��pUy�N��˾��'�n{'�x��{���7��ៜ���D�m�Z�!F_�!�7"7�|�F䆘�oDn�9�F䆘?��ӆh����[��{�t�=�������������ߧ�/w���r����A���}��rW��/w��|�?���/Z�}��/Gc�9{�����_�����	���	���I��������;�������uk���_"��^6��Y�}�Ԉ0��"7�t�� �v$rLӑ�0G�Dn��w$r��#�l�AC�r�uH��ت��-w��J�g����>t���?���#[O�Q�����İ�=�H#�����
������+�h���/� f�v�����w�ջ�{2��>|�b����<^��PF!��3��vH�e^��i�w��`@{�Ž�0�Pz�c����o�*0*y�����˭?���{�[ŗ Xn=��� �������l�a�_��$���Y�K���xx��⃐l��e��k0i���s����"��|�T��eH�C����$��$�B%{�%��#�*�p�� �}�aL��v�}��e�&#X~ �` !���`�����~�&y���מ/��Rf�af��P�P�x]�o.�@�_s��0�����OY2�r���-���F�2�A'{u��zA�>IȨͶ�f�����ut��Jn+��ʋ�������FuЫ(�kl�*/��W����{f�4�5C߻���c/���(v&L�{����M�u����_��$��c��'�i~����=��S��{���` �=�����N_$�!�ǣ�3"�j��&!��W.^���dk���*�)����8O��"���>�p����pZ䃩��O�<�}n��,�6�2�}����Ƅ�-�ԄA���C�����: �D��Zh��Vc��Hs14�6hXYaR�`'|��[���@&���1�^F<�o���[XaU���'������<'�~�`([myނf�i�*����ݶ���!��v��>۝��k���jN�k���d&�X��YӺu(�I IQ=ƊSk�OA�3'���އ�$֌î%�NO��8U4�c�b��Ԓ�K�O��6Z�I�j��Zj�<��]��g�ca��z-p<F�/h��D���aT*÷T� ��q8��$�-�a3�.[�_o�䯆�\�4�� oqMb .� �n��j�f��>B�*|�~{]�a�հ����y�I0�>��֘��#H�����&i�xa,����Ǆ��;������Ck�ۓ�*�(�8�P���}���$A����r��r��\~��$�5� %�3�M�[ c4d������O���[q�L P�d����� ʫ��Y���)uPm�j{����� �5��!B��J�`\־���J��d^��HX0ٕ����^�����4�5N��H�����cB)$x��!���P�KS|�ȱο!�	uys��K	U� �{n����jo��ʅ�`8�km�P�FAm��J�w�}���1?*A�?B����F�K9��]P[��pH,�;�/1�T��b����)Ӟ�����5�d1�t�X�z��]�*;��V��_��!�]r�|���ɾg|�#q�?2��e0.���L%�T�X�א�:?��y�+��k��SGU{o�jIT��s�	$^��0�u7��Ԩ:~]���ů�����5b��Q��s�L�Ƽkp,�m�0+�Ä�͙�E�/v��X��5�*�;\���p(P2��~�BG�i���-��Zۋ/�b�X&�t]�q0�3���/��zX �+�9���F����;oy�;sA�<y�uN�2�v'��d���/����5��/�y��|f��ܥ�`�̵��a����b"{�(��d�/�!{)j������,p������L�K�3W*�Fu,vA����V�w�;���G+�J:�9�6f�� ��3���o�&��y/�r�8�dW�A9h��67����*��{.+�qj�>4�� ���w'�,�٣#%�t�l��'���P��#�(f�����^;��셱�ٵ�9#��Z�#Oy钌���N�C�HQ��J�j�z,�x��N�#�A�뿒�r�<#k��"��ʟ��͙g�,��,]��h�ӵ}�խz���+��K�|>��%�F�lRk_�\p�V��愄�@Z���%�杇�pm��M.8m�c/�Я���Y���uf�o��z�P�\K؏�{o�������Z=B�&D��!�\����p�pG*68,p���zԜ�Z�����������mpm�k;\;���N�vµ�]^������NQ�@���c-��A��k6!��9�"h���C�������%!-�I�|�|��|�=}$�� ��W�M&`���P� ���Ȃcì��U^� F������0�H��	��g I�P�)�Bm�Y��9�l~��:�f�l��98v±�}p�㭃�6) ����j���V�Z���&���j����"ۆ˨Νp_�,)���ͬ�:�-�>���"ڮ��<���uWB/D���gL���๮�����ۻ�B����[�@����V�"y~�� ���ނ�B�tL�[ɳ�9���#r��hK�;��v���@j�{���)ʜ�Ԭ>P�Q�6���?��������Ј�c�l���8?9�H��D�7��<66z
�1�p��j�c2V�2 ?�3DbP�2�h�S�P��!rSqʣ�%����-���m��Ӓi���\�1`83�<}�j}�^�%l]��5��Bր`,�j1 �2|Kx���N3�-�0D]�f)?�o����S��4�X7����{D9:���>ϗK.����C�V�Á���[��1I�A��3��mCq@���{��օK7h�5��M�Z���|���f����ҌooX�f:} {�{����_��{��t�+y��S�V-R�ThLx/�������>�{�V"Jx�XX���3^�G��ه����xC>`X���ӭw7�7v�W��#�[-��?��������o�٥x���]pͪC����(ьS����2yF��E=H�Qh}"��r]����b(:�j�%:V5UC�t�u�i�"l,��k79����IW��I+��El�d����԰+�☘�U�*�\�䢞G�{Q�����dH�_�ȭ��Z�I�^��m&'w�A�1�}f"��Ȑ ��P5��u����� �5o�V���TX�i��I�x��_�c7[4����l8��[�޹�H��s��s�v�$m������?�D��7ض<�_��F�L?F�H�y+G?(��eZ�ݥ�s �pF ��sŴ����@^��8�Փ�&�0��Z<�2 f@�1	:H�Dȭ�C�?7�"Â��!���l�C���p1�bA�'��
��P8��yhp����m�l��`:Z���L�%�!`5X��Kp�Z����gU�_�_�����v���4-	7����af�;Q>��L���yiƢ¹��4��r|/���g��-�]NY$����:O�,��9�}��HsY6�k(�a
�t
�J�\��χ|(�0N|alH��C�����6ըp汊��.*�Q~����rU�KM:h�2T�ݾk�(1͂�m_���(I��<ϣ��y��3fùxc��$�M�ѹtI̡˅Yt�l:\��,qE:ΈKۗ�հ�W�ݸݍ��]��w��8�U��}9��&·� ��M\D�bH�h�"U��	~��F��@�BW�`�HvA��H^NcH#�E�$/�q2��.���b��N�Y�0�����~in�l/U_���8���J��o0�D��&�"�LlƳ�	�[��t��Z��W�¹x�N�x���t]*��y]��.�~V�No�5x�Z�	E�T0�'���o��%�F��X��R��Z	Ĕ\T^"�Ʌ�g�1�X�g硬FD�
b
�(F�1� 9���X����	��P��X|q�A��VBW��ۈS�\��܌��2_s��y�3�G�� �K�Is���Vc��!LR=��/=�ʑ�����g]]�N���e���r$����@1���W�,�Bm�(��� �Q;T<OK,bW�-$�@�e�ƙ<1���.w<G���\)"�	J��\ \����WM.��|Ĵ �J�f7����:[`�&��:�5o���U��8�'��IvӨ�u�R���s_�Y��ɼ���z+����5�%j�<25�hsp� j����}���z�zQ���U͗��V�z�J���{T`J%���|v9@�9�����d!d&B��$a�6���N��&'�֭@è1G���"G�߿�=m��28������Y2�+�DK�:9
�PE��OޣH��Wz_|ݡGo���jg����%1�(�V��n@����L���# ��ɤ̺�1V�BQ�Xu7��vN+���u&pP����z��f�yܡ/,�v�N�8�'	�����`��1����m%F���K�= ��/ 5��d����8P1[���c,���BO
rJ�.'J��E e.ǯ[��`Tu�w���:+��y��d~���M�w��,~w���w�.��]�����Ą�0�����5ԇ]�y�����l17�X�yo%���4Z�}�n({A�(��f`s���+���$_+��r�3��Ơ3�^�t{(M��P�ب�෉�`�d�j�M���{�5��=��-��*�)GwQS��Z���=�p�{�bҗ����W��Kp{
�k3��tU�u{9�qo���M%�q��F��g �Ŋ�cwu�g ��N���K�B�E���D,�H��
BQY�N/X0���n.�(s�߱k<5S�8{�H@��-tO���T�=�&z��k�xel�pt�ݷ�V�,�_�4�kF(W�KU_���Ⱦ��k�/�¾����~��?K;�n��%���b8��vѴ�V--��<C�X��eh���%b���Ԇ�aQC�����y�~�'�!�y��JcV�կ������5��N8��ϰ�����e<��g�~���k@f�cث�F�G������ES�o!�H�1��i"ƽV��q²H-�d�q�{�lu������-=S<�끀����ځ��:?��Z0�O������3P`��T�VVAf��쀣e�@��\i؛�Cp��\�T!:�ؐ�c~��2f&�v�ߜᛶ��X�y���i_n.4��0Q��%O��g%����F.��~qX���Lj]��	o�}��d����=M�e,R�� ����"g!{`)�/�M�aE�ef(W�{�,7��2���sL��k��PP.6HJ�%jM�Q"�#=����|*���Ǟ�e���Zk!��f���ӍF��z�J)��֠�����:���(�M���V>Ne���Ȝ��O�����S!0�6սD�Ne�dw!��%��q<[)�"հK�5���ݗO+0z�8ٍH�yL  ��J��j����{c�'a��	je��i��<#�z�	]`�B�UR��١4�fď�T{<��`�ʇI׳��_�Ӕ�)	k�_�f�J�,z���q�1���� �'zB�cGq�w����ƌS�g�)�'�#�$��t�(��D�Rc%����|Z0�[p2�T��h�h.��T��h��j�ݨ�6#M5������-@�ǘ�%�V]��=�,nCN�z��N�{@f�{�ܙ�y~$��Zj�^v�
�V%�_�[�����X�p�X�,�*d������c�/6}y ���)���$6xgYK�K���yAZ��d� ~����zʎ����9&��>�?,%�sL��6e�Q�,1Ds?n��~6Q��IV�PQK�Kphۋ���~��J����cN������vT*�@U��P!�f�"2KΛ��&����?��P1���T�v�ʖ���������E���D�P��#����O�V�O5�G}7Bc�اW�����2&@�.��W�~�+��2��n�iX��5�C;��+�_�Ӡ��>W:��J��-y�M�$��24�C�0����'l߈�i-.�,N�;��Z����n��+^$T�8Ϭ^9vUh[�� �oB50J�5Sq^�,���(e���D"����x�T"
WW�6�d����\�ƒ� ~.� zs�
��`�c��JE�������1�Y]%N�iޠQ�(�fk3
4��T(�xL�|����r�9�Q|I��$��` YģJ��e[_����>��ՠT�w�
1����"��Q�C)  fߖ��!l:h��]�Н�z6"�K�n�6�Y�]X9@-12�`27FV�������z��!�c\پ$l������,���� s�`L+�4yƓ�u�F���&.�!�@���;B,6�EpN�U!a8���z~4�g@��I�SkH�� ��\Čy���=ʅ?؛9^S�T��Y'L���8hsIG�P���Zy�2޾n�躉�4�2gI7�-��.��m�O�{:���C�N��b�5�)���%�+�&^=��g��yze[Y����77�b��q��"P�-�4�R�)�!8Ӵ�O�4{�{0ٍ�&%�A-m��ʵ���D,��ʵ����gâ��4�Z$�x�X����6{�%�����l+f԰Fhӓ @֐�U��x�/��ǈ���\ȤQ�[���p�XN�o�s*�K#f�9�xa38V�>C<i�Q���&���_��<5���p�d�<��
�9n��߻N�<F�g�<���æ�qIf�����6LA��hHOu���:B��b�|fк��d��D�`B��|8�p,�P��aQ�Pk{h �Ƣ�Hb�����'�b
��CF����Fff�t��sO�u����a9���?��>�e��q?�W�'����s���#�Ux�cT'��_7/��ɥ�:s9>C ���6�-2|$���0�&�qV��=��1���3J�y��hP�_�,��劣����QC e����Ň)�f�5o�Ls4��TM ]�h��3��7��f��58|&���^>7Pм�?$�J��FP�L�Ak(/��!�]���j�W�_��c%��۬s���;�<����Fs�cP�+}/Z�J�R����P|����[�&��o�V�:X�oo����f��.
u[D�xb3%2�x>$.��>��o���x��d)�O�T�<m4���w2Wƥx�������)w:X�����::�JL^G[^��xW N�;t��0��J�iU-�$'��q��B�"�)U�gs�3~�i�ϋ��)�&�P�[��`|�}� �i�xb�1�/��X��He�S��E[�b
D��ǰ�E¨A��I�!x,V��g�5�nZ=�-C���o��;+w���p+��{���ƒ���w�^���
��?���(=`U�|�ȟ �/i+Cf����5m�qUb�ݴ�O�q7g?��x��pC�:����o(V��p���_�l�<�Hb	�:�c�i��~`��qFC@�n��5�~/�$:]X��V���{˗j����� �w�2߀X�����P��`,!<�v�|�C�&������ѵ���	��.OǴ�.w3����/,V�	��,�|�}9f����U)�Y!��� ���!�+n��'BgK���tv~+� ���	�V��Bn�����.��<�.6e��>z"��G>	M\@Q�"�8w�v�����r�������n�|��f�����)�=s�;Ks��%�R?���!��k,�F���������Xg�6��b�f���5���x_��X��W1H&Ď�ߠ)�6͝8s�M�S������͜9kVqf�;������
��(D���+�"���z����N`u�X���h�{!��\;F�J��I�*�c�rN�ag<]�$��� E)�39;>���%�_n3B$�x:q�Z)�_V�����>�;y�����c�N��pZ2�ؼ�?7CҺ"HZ���+΂ӽN8�Z��W@����>H[��֭[��S�����7x��Pgi�x�@nKQJ;�!o�'�Mj�V�mǑ	G���x٪vf|=B63^�c����2T�)��Nq�����M�o�\'��ֶL�g8x���Ÿ&�pb�1��-�q�Ieq��iSK���Y���|�3��I���B-��0&�L	��e��ř��fk��z��U���*Л@HU�Y���0��B���$�^l_-����,������1/	��_�:㞢��4{#)4��2|s�~*���9w�|�n
�6Χ��2�{l��>�1w1~�Jq��O�T e:��'��lQ ��݉8�	#
�B���g��ͫ���^�y��%����F����ԣ_��n�H=��XE89:m*F�3p/�����K�Ņ�-X�U]��4���
�E�Y�ˤ�k��D(s�Bm{�&����vEѴyƩt��?���z�x�����g!�L�km��
@��,�l��㴋�FN#H���Us�ћw�~L+R���~���A�N*
�(b��B�C��gs��M��b��IpN��?^�0��&���Zx��u��A��^>-
���X��vz�O�vz�����;��6�mPk����X��d���__m���A��@�@��x�IE칛� <#���qd]�����?H��߿�=��h�:7�I��l|h�8+�r��k$�2�gƒ!�,�W���f<�����y�:lM��;:�iZ��*�r��fV��c 4ނ�Wʹ��4ɇ��?7�o�y؀�l���ڟ�]|ȧ�u��1כr�:��V؅O�@�0�:�󸫿6�(}��koQo2d�d�d��E��u�#�#'���z�����9;�s0n�?�{cs0g�ރP 2�a�Z��Fu!>����Pn1�#xp�7*s���۱�Zw���抟�	`5wV�1�\�xL7-�|w�^}7���KA��7!���������oȼ����O4�I}`��ډ�N�9���N0�׍��罩��wsj1���@X��e�mPo0*s� dFW��ǘ�osy=���5S �QYbP z��pΜc�,� B�t��VW��e�f�3X=Bb=�J���$ݜ�9l�K�b�Z`�����So9�= ��T�)9��T{{�h���s'����4����Qq��z���\����������=�i�[5��3��*�2IK=�{��k){�:�3@^f8K)�p�o��i�)�&%VX"w�
5�<Ps5�}B�w���<o�5��C�n�A%@����� �c�R��>i*=��ӕH�¥K�TM�_`R�Ă���,�,w��Nn4�42�22k=�`�9KYx����NY�up&N�h�pש2
�kK.Y$v̢@�x������U�j�[�S�c@�Fy�H�*�Y�@�G��yԉ�aR����'$����~����^\>	{1追�%˨d�����������c�L�%�@�Q�D��,��	H6%�a�Ā>"MS�b���@p�6�a+�j��Ū}��ʇ�@�؄�E����F�zץJL	���sg7�@�}�}~��2;w�=s�~�{�9��sn�x��]+�gh�	}&�W;h1�de{�\�?�,"P���ze��7��P��霮�E�����}pӜp�h^Q_>z��|H���R���u4	U��;�2A�.o���M��O��~�iė����=���誦9Ŋ=u�@(C���C�{E�u@ZSO885C6f�z����
�h�>���C(Z�~{��i�,�I�M��h�N �ҏ*!��Ȝ�#�S��n+Y'�N@���i+�k�͇��Hp/�bN�N�.��Y48�Jn#��9���:��8���.Bn}���F&(���쓥=���rG�nξ�O5��-ҫ��9g4�����Nm���& E�M�_�|Q�j��Td$R�A5r��4ԏD*�f"	�l,�ߌ�R�3x���H����8GNZ&Xrc�&j��}@�*�R�6�O+�1�b�3\ 7)�-l�jǵ���v[_�.�t�P�0f�P��J{@ޕD�>L�%@�o�O(�8���''��;c`B�CJ�y&h�DlW��+�[8,`ݝ�>X�t��WcSjP����9�A�&ǈs���1���]�D_b�R���f%�<�3!qu�Y�$4�ǩٵ��>b�<�" �"�${1~��ɲ���7p�_U���7��B-��a�v�^�����8M#�w�������^���ښ�U���u�}XY��ƌ���9�,�8�DK]��曩�Ҏ@�%�m�M#!&p��S��`�Qc@�ͩY�b�Z`��FS!���H���!g����5K�,��\K.���J��X93O��H#�����gHm���7���+�+#̌!���E@7;f:�n��=-���&:�p_��J�VD�[���r�%�����7q��� �i�'����D��_R\z�	��/O������6Дȡ/��_�7�t\!,?q�m��(D�;�����Z�����Aj���[E *@��r-䘙��D䬿��>ݢ�����2՝��}�k�J�i �a�� �\�ךL%��/RoB�`������h��e?���n�aݭgW[�[ʥ��8�Bs�E����^�QHV518C $�7�7�-zI�S[����P���'�v3������4�lq3���R�i}E�d!&������k�Y�'�y<���N5�/����Q�>h�}]�T���[���)�H��hrp+����84��O�g��E�Y���@��Pf��!����-PNh�L�/�X�ł~[-k���ē�W����E�ӓa�Y?a2����m:� ��a}�˿�	�cj.Y������5��+��I�Xk�kda<�A)w�ue�;Z8�!���-򖾇=ȣ�w�2��"��5�H���X&B���?`��R�\���c�!)�[��� ���C�;�,�wr*�m0�]\��H�J+��{� �	��8�GL��KD���(���R�tTcd;��?�s>�./`\��mZn�8��!Z�![��ߙ�[閶��� �gdm���5 ��36ܮ��[�����*����6�b)"#�?��/���Z���]�������=��,��zx1&�,"6WO���UQ�*�pxB�lh( �
t� ��3�j��9U���q�l�����6�cj-AO��x�3nbZ��7���'Q�G&4��'x��Y��Ηܕ1f�+�`��k�ͭW6��*v������I���y���K��:�\.�e��&ܒ�<D���<�%�K�D�~8�)�ɑil�E�C���o6v���Q$�p�����O?�����{]��]dK�v�7]mq�"%�*�+zoVE\�)R;������͌�ɭ�M�-�?��i<.bN�ʂ�c�QoG_�>Z�͏��o�}a?�2n�l�i���a7| �֒"
������nh�0�[� ��9�����RhEu���X+�>�� ��@��$��!���fk�Bd�>M[+��0���s��ș-*Z`�D�K��E�WP�
�/�1���8ܚ\�mQ���KD��5�~������w�[��z�R-C/�A8�=��GG��6��l��sq�^*���9	�u ]d���^*@lO�2����-��G��4]���Ll[XM��P��"G���E�ԋ�/�b۾j :.q��$5èn5����3����4� ��k����{�eݧ����t�&�~D�Y]\�P]krd���n��^����W���e%���\�8k�Aҽ��m��@\��	Y�$D�ΤCq��`p�T�8��O����7J�o�o7������0��Z��܁�*.f���R9_��bg�ah��
�[�4=�Ի��EI��4���+wH�.ruh;:)����>��w��/R�z���-���eѶ��i�w >8�s���R���v6XvZ�j��8&�l��cmJ(*����;��ïRA~�d�Y��5���o�6�����k�� �u�/�WT�+ߪ2�|��D���v9���S��^?�@<l���z
�����Tj��Tt���u�8�U�ݠ/�Ӟ²�J�i9�Rdx<��T�ﶤI��K�����<��N�e|����͌?1cj��{"f�=$K|�y壳�*5Z#��ѥr�])�c��@(����e�r��׌����,�J�U�^��쓡+oR�,Q��&*�j�`����2��8Ѝ�yB(h$Z,5���w�F#�B?���!Ej���*��#�'5�%�qZ�znp"];� �k�,~�7)f{,���g<J�����%�תl������.�D��ݹ�jdqD�[�H�f	n���i[��pHH���N]���xw/!�l� J���5Kb��<^�/�0R�vas:�TnV�'�F�
RS�3TG`���	j*T��~�0�ɍ-R�E�DD���Ƣs����T�B�k�#@�T���Fi|LCRc�l��6����)�o���x~�M�7Π�~իӭ-�g,��үp�to0�G�%�{�钤^Ҷ�G��%�q^Gm3\����h��L��`�]�U˥]-���#~��{ 9�V���i�����@z��ӠevD�e��_�*E�����>i�~�����0Z�E�#߯F�/�E���xs4�mPwW����Y���Ef��c���	I��re�=�����"j��D��!!�BE�iq<�(5�����t�U�|� ,�V��xI�aU�^����z�9���N�����ڊs���8 @�_��l��`�L�����x�����ol�%��ml��	Ğ |Ï�M0ѳ�{�z@
+�����$�����S��,�Ƥ'�z?�u��J��'J�A5�2^nv	T���`X�G��m����5����R����Q�g�+�s���2�˝$d��[;a��lU[*�y��� ��uN$�<0��(�m%'K���"�����g���4hf��3�Hq(3Z8���5 �-�{X=d�}o���'7B��G��ٲ���T%��KTn0����J��4���A5P�7h�
��KFy�N�^�GV����t���F�#���6�N�ܔ1'�#����J��!m%���GFR���o(� �1hP���f�P����:��H��K���\T0�S��|0�?������"9�l+Y���l�{~$y�Mά͍�j;5 ���\�2���ԱxO8���-�q(�js�O�"9�؂P����`se��U�eq�<��eD��v�c<��;��z�ޯ�഑Q?��d7Fo�.Wy�S��j���ak�5�<I�F������m���0?��u���AL4"#y���"�u�M�oM�Yh������,9��<�؂��qꢸ�:g��k	�~�ĩ^�����PV��]���}.�Ѹ�k~�V��Y�cV�s'��.��-V���K���YH�N��j�Yªt}x�Ͱ��qH;q
�^iZ�(��d"d��z���#�������yD�I��E��f� �7Y=
�2���-$�͗�1T�!���a�-Qz��X�h\���O0�i��BZ��N�]����v�4�-��l��Gz�I��7C�3w�6e��Κ��������zJE�B?�)n�� �p�Q�ht��G�h���O
}�lwlA{��M��3=o���]�p� �9&t:)ԙl�&��)�mTo�p�Q��y�$�� ׃G-��Ǿ���CR�(O1�,���K�!�y���)�V��i@8q�D��9W@y�,P~��E Ė���H�LM����-��[�1�+P<�9T<)+3œ* ^��i�5�"��$��œl�l7�x�.�~�������<-�s�}
��,�A�%v��%�!ZL%�pH��^=4[F�����6?N�!R.P.��ʆ�k䒆�A2i�$�{�X}H2���K����H�K����;�������n�O�I���u�rqq�Ն��� 	Lq���<(�p�� ��w��ȟ��ȟ�b�������:��Q�m��啶���Nf�BҬo �͗�Ѓ8��[���f{1�,r�ϡMr"ă���pDAх�:&���X�|_ y��%��I�+ـ��Ƴ|j�������3�Zrp���4�7Q?��� $�<O��ȥ�',��I�$&+iI:�zd�WI�i8�Q*�?�����2p�����}��	��a�Y��D��	���A�:?���~B� m��筱��T�2H�����1�D�G�<��ɴr�4#���T�I(r��ǀ�Mv����/O�ߎ�-g��q0�P�.;bQ���ǩDס������q�:�����ZL���̱�d���1��J�e���efK�s��[_#�AÇdD<S� �<�0�_
��V�?�2�N�!.u���S�^%��b��:�7��qG'j���F&��x��1M'�\߆B��	;`�ڢ�q6&t�nAL���{�Ճ}bG&��c���4�&����s
#�o�bb�g;�ر�b�g$v��A����3���;b��,*��	@$t�$�&����$����I�`g�B�ٸб��лQ�	[��q6&t$�9:��� T���kBS��g���c>�9B\޸snzB�r6o��P�3IΘ	r�HhP�4e�8�(��(_���X���0H���|G�/�L�"5b�:���ӉAD%Q���s�"g܀pA.�Ƅ�)�,bc´��B����o����$�[f-�x�����|B��X"X�!+�2���$������;p,A��E�$����ʻj|$��!?���p��˻�85�?�I��р��Ah�"��,&f ��c 1�Lي�b/s1�����A���11I��������з$Lے� ���AO7��'��[�^q�TV[H�r��剁r�w��(���-�-(]`
I�9������1nkbe����&ăq��lL���ߒ`A��4�6ۛhVnl��#�R� R7D��9�,'�q��_���qa�չ�au>���*fu����vH�����M��)�a=Oz���nPj�js�1^�����R#�Ux�[m�~�M8�D&�	U4ڊ�ҴUb[Q���誴���ᱠ�h"�LՇ�{�C��;T�ƒ���Rc�����q�M/���[��I��klz�����,��6nH(���Π��mͪ&a�r��D�%�H�[�4ܝ�+�zw�%V���wݻ���©����"�:���:-c���#�ٯ��+��0n�,*��-�c��t�mhf��Ч���ܪ^�h�Й���K^V�Ǘ4����Q*§�U�q���s�O\G�S��$� ŋt/�����Ra}਒T�3/�����բ�|�5wF�*�oq���U��6Q��*lX���ER�q� Aq�T�^i.��%��!\{r?Iwg��`�p#빗p�#2��I7D)6�C��>K���*}C������(�g:���Ouk/J���}l��n�UL�ZXߏ��kv�.�T/�(I�6�SLBozU.��Qz�5�2U����ס�h9يK�����*��rH5_��u�y���H�n�7�2u�|C��ǔ-�W�)�A����Y~���D�`?�p�Eyՠ���"�_�A�z��=���;Ts��_ �0&���� ��j ��\-~-E�;Á:�B�(���G�� -7�r��D����_!=�R
Q�)FJ��,��.���|���HZŷ���H#�N�I���Ɇ��d-%�7g�Q���,����IgR��CNB��l�fRc�����T%�4rjN�J�#h�5U��N��:Z���J�7�r�|K{uOȪ��#JP����
Eл"�\-��P���`8�!��E��5*ԡ�ĺ@ʕTF�p۔Tyf�<U����+���y%�5'C�x匔��F��Y&� ��QF��zJ�͂-�/8�dN!.\��j�Űhe����ш�����X���*����5�^3�jZ<��I۹�^
ԭ [�kJ�^هZ
>_������б�T����V��h��z4��-(H@o�_���ָO�ך������A��Xe�>y=~q��h�Ao&�v�4@���0d^��U���w�r��.�Ȏ�$��V'�%�]�����=�	�$�C�*�Z�WI����%�c䌢�%���i~��>i;d�����}�E�*�O�t�j�(�ʷ�썗�qG<]��J�k(� �Ɠh��Ǯ݌h��T������|�T�A#�%rI�>%5�A\&�AS������"/|���2|(��od�
�{��)Q�b���	�荚Ϳ}�^�s'�TAMۖKz�i�.���N�ֲ{#B5~TL����^�N���R���w=��Uh(��WX(g臿{ԡ�������n�þ۽g�XX�%�{�hS���AL��38��$)�ր�?�����ʜ�Q��ܡ͹�>��؎�d�O%c��������ڻ�Ņ�E�Jɣ1y��C(���5��E_�x�,�%��t1z��,��1����3���3j/Fn����s ����=?�ϗM}8��>gL�1>��s3Ή+׊�[󵵋#)X�
�-@��Z�݀��N��ŀP*���&R��J81����(Q5_ծ9������.�ʩ��E?����8Ȍ�7!�>�5���D��=B��u�=] �B'5u�<]�.4��y;�I�RR��t�wi�����6	?�p��z��f�O2����s���G��A0m]��k�
��
�>y��R��V��n�=�~d���R��zت��{B��=�7'����Ca��|�E�8��}�p��E��+��d�n�������v�s�=��8F�)c�ڟ������_����q�-w�'5E���]=��F��\�����mܫ���u�;��`�\+���pxד�����g"j�q���pH����7��C��`[�0D�.�J��]~V��dI�:��N�'�F�
4��9�J�7�Z��a''s���}�ZgM��8x�I�7����9�{��bŁ�l}lݳ�@x���O��3r�݌�~c{y�}l8U�Ӊ�{�*�>��SoƸ�$4���g���2^������lz���q��RTA�%/��g{ɭ��(�>I�>������j�!�;4�4��P:�Qf��n��&�N�rC��p��7`���hY-B�/� s���C
�N��W�����f_�Gg?5�}��N�[Ǌ'G�HrX��$���O%9� C�N�'�Y��<zcş���L۞{|� ��oC��G *��������x��w����]o�J���F��V�<����2�{5�CxZD,���N�����bx�es���V|��_�̶��+� n ��X��c��g<C��K��"�!Tp�oA���m��?���ȶ6���ޣ����03|��6�O��N<�RO���0��ŅO`���^����6�7�k��W\ׯ�֠'��z
!���e
.�G�3�����;�rQi����q�k,�&�qg�*`.~��E̋�^I|hx.��^�T�n���!�[,Ğ[��V8	��؁�`1���=O��V���-�n��f�s��	�^yl�V�B8�z�Q~�];�|EZ�O�-S�l>�H��a$cH��� ��/"R?CZ����+ԵK-r���-%����^���6�DB�`׷a��,]��'M�RY��l\��� ��?�������-ȟ	��*&;�Ȅy� X,��GЯ ��p�u��+�`iN��}Eo Ҷ=zH[+���ZG�#gz(����/���@�Rp��]�bs���Yt��|h4r��!n���5["'i��cU0��ƅ���u z{�����M�IX�"w{]ws���Q/#rA4�>�ԗ_���i�ݽg�E��"o��a�^�;��!���f{1��Ѷ���[�����^��Ö�EB�x�=�;߱�*x��V��d%&@_" m���������K�h��<�ټ!	��G�}Y��Q�Qӆdl����HVug��[�=p��9m]^Ka�1�6f`��@��\��%+�3�+v�F$��KVf`D.D|�����,���7�v���Mݶצ 7-�l�HT�r�7g.�G�� 7/�W֘h��+-?؏h9����DK є��I��{��K�	.c���X?{����f����;�MBL�`0|��q[f�"A�˻�`W�ћQ.��W.kO�l�PF�aȨ��O���Q��eg#S���ʈD��� ��߇�v�E�@b�u|7�:\�k���=w���6����G���J0.��pĄ�B#!師�p{�=`=�_�W[&L�`�g�vWᗡ����b����\�1j9�q.Z8z��w��r�A��`q��˦}<4]�= h���Lz7�Y���Rʗ��R#z�����`���2(�(��R~��n�M�����uͥVgc����24YgsC#$�%�ѐ�u�;��s ٥��s���t����dP�ۡh��")Z~���d��,v��ϝK��/�&L/*�U9��b��m�
��"whE�W�'��~�e��$� �E���@��Tf)vh>1bז�&����T�ͅ������~Z"�/Жid��� [��w�_r�T�����@3����.��*�\<�O���Á�\�|�	g�5��SϫW"'2�Y���&�Zh�+��ϵ9B��5S���=�<���>G���e6)��eO�L�x`td�Ć_�����h�&>��϶L��<�!�T�\��.v.��_AtQ�Q�TD��aͳ�s��V�aB�' �������!�>5h�Ƌ=�Fr����q>�/��	P�Gv�P�\�0����|��b?�S���X�V�_wQ{���[�7��g�����g����O�^꘿�A�bVJY�sr������"y˧�+�k� M�l�/�
�a���$wQ���2�R�L��R�c�0��W��@��XۯLS���𫘙
�����I��Z�{K��U��~���,�j�����,�m��vt�_mM�\S,W���Wqyr5|�`N�LH��~���c�ᒴ�ez��\9����U�ǀk�r7�t}|��\l#���UA�H��#�9t��j�S���R��q����sx�`��h_`�_qs��~'�o����0�]�6��f3O��y�ߛ����QݙLG*Ջz{(�4�퓹3P{{�<��g�-c!�����߆36\/�*�rg�A\⼚-�/@�&�[�|��?.��P#G�����<�9�U�_�Ƨ k�䞒�AjD5mV�t_���QX��@	�GC^=٘��s��^)���n�8���F�^��:Q0z�Z�2������qJ�@������,֯(ŷ�{Jש֮���i�T�luhuU-y'6Uv7��{)�6�S��&�y�q���d=����g/zP��#=�<�ö`�诸��j.2�4�+�*HdT��ǁ��$&(p��ڤ`ywE�5D�
���e�mdm7O,��ЫL�j��c� VJ�@�q1l�kQc�^փ�H�P�)�\�\҆,�,؁����ϖ�<�	��y���� jD�@H���M<D>���o�)VY�bS.���\K�~h�Pq�J��i[�~��M��űGpi��I
��w(S�YN���a���Ń��T�*�F�8�{҃�Q��H�3�Gr��;��z�V"�3�_��ʀ��Y�(�� �p���]�]�v���1Ib��<~ʒO�����ܹ�Pl
��GLo�:Mq��Y��v��	�n<�s�?��2{��c�(�T^��R�ܭ҆��ͧ��aL<�N�¹����!/�V�ܖX��Ҕ�U�T�Ry_J�FL��D�j]�R�l��,Ѳ��T��ͼ-ќEE�	g��~[���������i��vB��a���f�� ȹ�qZv�0b]��@%�[0`�OU��u��Yi��_�����`3���]h$ZS9;�"0^�A�7?D�G^=��� j����Ɵ�������y������`�a߂����8���|��+��|@S���4�F_��C?Ę�6�7��<fe���_݁qe���`��Ii�*�ljc�`�F��"���;�}��`"��"Y�c���R���cgU|?�O��\�3t�T�|B�E蔠���Ab'�5E�Nօ��h�2�u��.���KL�(x���M��u��M ����p|�w�O�mo��ޫ�9�ۮw�n=]�9�A��*��_n��b�)�  w3p���\/r�2�	�OEo�C�J��Lr>劸�b��t����<վ�x�g�]/B�R�wck,n���H����V�?���n��¥�q �t�A�o� ����՗��T�6/;���j�)=%�P��D�\2I�b�a<&�@;ص�����K�����,u�x�i�w�Mr�僎�vq�*_�Y�/5V��m ���38}�גј�T�-Ҁ-2w�
���Z��W�n[�}�V�鞊�����Ч6r�no+̖K̃$/�}9 o�v�+��5c�����p��7 Hf7��M��s�gF�Z�����]\ܮ��R5�Q>�8*�e��X�q~���Wz'O����ł�VV����'x��./��5���v{���N���b�c�ꋂ3�[D�{�X����78�	�����b!�������&�����2�i~��U�P��&>��'�=F�N9t�GI�͞��U�Ĥ�=;�5�|�;åo��s���e���H��t�� P����2~V��n[5�L�#�9�~�[�b�`z����N�eI!0�S6}�=������KסWӭ�X�-=�[ߝ`�n��@o�eS�{�m�3}~i��ɮCU�1;гb�-*s�Oץ��D�����j�X��u�t4����j�kZ���}�w�3\�TO�3��?y��14�6�P\Nvy_ą�J(�x���/����֋�BlL���s���c�;��'�Y]���"U}�!�Q+�tb����4"f�*��Eԏ")��c���'`[k~�מ�	�����y�g�LL���ۃ�#�`�~x�c(C���L��-Ӂ$�����Se�(�����N|V�Z�5ę䃐���7�_=$�t~�p����WgO��Yə��'�q�X���Up�S�Wc�>����ϯ6�8�dpu�u�p큫��p�{ίƏ�V:��pM�����7M��ί�N���󫟻���7���pY��ϯ����'ί�|���ͼ��]p-�k)\2\k�j��Ӭ���y�����ױi����	�ͯ��e��(c��yN<����øo�.��w1�����n?�	� � �`��у�<�ޡt��һ * J򜽟��e�n�X'�vE�|HuG^��(�D9z��=��g���o�G�;w;-P. ��,Q&�,�r����f�tk��_�y]�lkWa�N� �ǹ.ї9��~��w�MT����W\��"x��z�V�P,��(��,y���*��C6<D^Z�0��ま��w��<�w���k��Vva��2ѵ�}�� �Y���9�e���`��m;bwk%G�_kܟcܟm�?�e���K��ʧ�zj�C���8��΂�\?���]��R:������S�ˬ��7�]*�; q�|W�/��Vr^&{�<wa�hIt���Q�������7�BW�'��
��]C\���	��1td?=��
�ӌ�#W�"��f��Ary?q�+|ٷg�?�?�>��+�� rg��w1o���~�Ę+�a�s\��s�ߵ�W�XMvx�?�
ݔ�)��ǳmZ1�x�'�c^Χ�NA͎��(�Tfܮ����Mi3J'�85��_1��{���4D>~�j�3���KB�s ~ӭ����s��jHx�\�0}z�yc�q9��-��pWG�E��n�W�C�������x���)ԯH�9%&d HU\ �a)q��$������4f�s��Pg����*��E��\�+�д�J
�DF37���?��+�����N����+��R��I��Z�%�����ܜ����\���n�Mjd�-|�<�2z��@FO�(t��Y�ƟSF�2z4!��!�:'#\	��킞��$�T��?�1������'R�^���N0��F��ͳ�v7�z���:]ˈd@N��{��|�c��g���ḱ%�V<W-�W�3�۽fU�m�a�6����?��Hb[J���'�%6>�� gV;eg�e��(�a�u�����_n%�g��2�1(e��5��%�#�^���5��P네�z��l��ֵW�;��V��c��B�T�kS�e���$��ǿ�M���,�ʣ�|��I���N�����;U��zO����ĜӗZ�����:�kR �"0O�X�x���s o!�����G��]���P�m����~�5�S̢u��s�ji{:G��>���[զe�Zh�?�UѠC׭ņ�:�#��I�]m֖X/I�'!���Wq�d�;��&�i	��^��g�BS�����c����x�*�c.N�7A��)����:��j��C����d^��v x�]� s	;*|U�Zk�<�§U;�Op�^�,�vH���Ѣ{��C�F^�)!����,P���g������]�V������f���>�L�S��
�)H2�͕��wXG+��9I#����pkT?ow���_��>�!����#���eKD4��F󔄙xJ�L<%a&�0OD��'"��f.���p � '�;,>� `(S���uZe�{�<"o��-�"/
�݁C���q���@�n��P�S�������q�����.t>\���?0��RA~�̃xq@��E�3��$W���xNa�2����&*_1�]�/��bڠ��虘d�/bj�r���O�"���_�@>�����b��u�6v��V�f����~�i��{��ފz1{qw��ޡ�����N�'�g�t�f[�~�=�_�=�=M���q��c?����'��t�a+�^��O�)l�jl�"cE[@Q%�G�2v�g�b�{���w0��|��Ů���l���t�a�t_��t_��੯+dv��X��k�'�x���nE�l����-�vQ��b�Pp#_� zSbOSM��O(�d�5Qp�)��(���-���O��p���N"M�/+YEG@�$ٌ��bV��I�2��N.��d�^�p'�1��_I�8�If�	��Nj4c��1��&3f��q'm0c��\w�F3�9�Y����Y��L(� #T&�/x�}��e�#@��4�?�-��-��m�^�"'�Nj���6'SR�UzV�[��R_�]�( ��"��b�����&[��ᥫ'�cU�J;.�F���m�%9|�=v�	\��[H;��aܶn�r�Sm����&�)�ن�'��gP x�X�nԛ��[�C�b�0�?A�;Ԑ-�d�6�y�t+���w�ݪLFMzWO�����N�^��k�02q��I777�&s�r�J���Q��	r{Zu��:��t����'9���:�H�@�p�������d�"5��k��7�`�]91X2M�j,��#ٓx���0崃�|�p/k^A��ʩ��V�ED�;Aa����ce�0V�����e��3�6��ZV�`a��������)�����<9�jb(9�����3��ɖ/�����
4l�O���]  �|}L��.3A��1�,/���P��I4x�	\��"���D�МO�
b� h(��K�q��"�Ks�̂C��	��BlG�OK��q��	�����Q����C�¢�4|F�#�JS$���J�I��[X���
�<S�8gd�b�{���إ�P�ۓYo-�<��Dc�++Ǹ�&ơ�?a\.T ��)w ���2	��ø�!bmqm��м�^ȿ��D��:�\�˔�b���������n����1�n�9�s�\���I�&> |xWߣ�G����]�ǁ����IC�<Gz�P��>O|3�3�{�Z/�I,~a�$�,�E�����݀g���X|�M�\�es��3n��0 N'���o���
����E�c����r�'���v��=�5K���5�Zu���w`H���
yA��yN�B��˱�=�R�Q��C���]6�֖�͡o�DjP:��l�^�lz�ې�LU��+���V�p@�����﷧P��S�L�;�U��*��ʯ@e}U,��ۿ+�*����_\=����t�E�����	�=�\�� A��`Tϕ�:[|7�/2��űB:�W���m�g�O��Q��-���3N2�[|�ѶI�X"y�c�8��������#����BY�Mh�ve8s�[�����Dn%ᴯ�l�����H>��t%� c��$�k�0g�5,� 4�E��}h2V�YS�,l%��~wU:�5���b�K޴8^�6����s��W/�m�E�o�߹�����mr�jV�3�lH��Խ��;��˞��L�$���W�sL��\���R?|/�R?F*�1��,�<���N��3�6�Ƕ�62w�L��k�+����Sg9���٘Bpz&$A[}���#X4��V��0�Mz	��թ���ٯ$�{�-�g���&_"Y��B��r�:{
�,��:_�)���75���MB�+����dd�L�"��0���!�����E�
#+���:��&v݃Hޞ�Y�"�'�[E���j�=p����,�B��ԥ����M�k�m�D±�U��{��j��0Ė�>���O�Hz�����zt�1!�|t�>�9Kg)#}���W�U���1�rp����d`�"Y��Ļ�oԲ��o��U�lv���[�I�x�-�]��y�y���!,���6�C�+��x���l�e!?�V��@�MUJ�w�'�|;���rSm{�'\� �/�B0�su#�R1��hV�2���NYK
�I踋���(�r�W�q�d�V5Xbu>�<vJ���p�YX}7wCm��f�L�Oo���)u���~�Z=��~�}�<&��}�Z�I���M��"�Q�h�Ӽ���X�9�Z�C�׀���)T?�ҵ��uoL��Y4X�>�<����*;03�zrh���s)�O�㉺d���p�@��Z�S�5��_�B���kG�_���T�ߩ7�	���M(S;��Q|�I��z.mN\e`�5���u3�%}��J�B�\@ǧ��@'�c�C�|n��>�v���|��w�\ݛ7�e�^�xΖnd��9+���59��_y�%y�3 ����;W�<Y]�7ΐ��r޸�W��k���u����E���]��^d�,f -Y#۰ئ‹y�jY������Aq�}���BT��j���?� 9����u���w��y��/�-X���Џ��V1=�K���D=t"��1M�g���m���K���,���!���kmj��[!:��^�v@}��A��͟�S@y�etZ����6S=�6G1m�IGL]������Jk���6z�q��%G#��>�[-.Ѳ#�Qg�?�����>��p컨��o�H��z��AlA�x��w?'%Z\�E�r�6H�8v�]�IG�2>����W�ÇQ�>��Lۚ��[ת���5_��x�Z�W�(�8�9ᕶ�֊^�N��|$>B�[[ap�P;q�Nj33��pf����g�"Ig�;D�rÆ�L9�q���M�����V=��;-2�9e�*yؔy���"�C �xE�ԨS	�JA	S�)�L���X����=gJ[�I�szB�,J;���	�Q�!;����y_C���ӗ@�J��UC����@��BO_�5��޻�rx���+uO��E%�o�z�13�@��~[�i?��U�w��fA�٪LU;mr��z�jX�
��/T�V\͞��0z<�V>dh�>#"A���2������e�i/�{��u�8���0�o<�p{�d�
��**)5^ ����x�\�~c��b��#�Ց���E�Y36%{Gol5<��U��Ɏ;1`ȸ��������bd�qf+	g�4Lf�1�D)��y	R��D#�^"�a@)��9�[��?�&O����S���qH��h��Ȃ�-eG�y�ZϬ�<44æ�e��(ʣ+��=o#5��v���cR�+u��]���Vs|���L�[l?:Vy�_�)W���z^E�Y4���O��0�r{�& <Q�F��������A�&��3�NjL?�e�]�W���P���!D�xPH�[�������o+�H�PTy�������fZP�| � ���Y�Ҥ�IW�r�^~@�b�!Y�3x_K\r�܏}F�v�G�����T'�V�Y�[���"_�mD��쑟i��@��*?C�ƴK�}���~���ӀK�V%]�)9=E%V�"`.���V=���+�>L��3?����#n\I�=���whx�07�D K��U�Q��G���ikb2P��&(=������Du��+ͽ�'a��`alC�?��|���[19-��>S�3"���ߤ��xԔŨY�9��"����[�4n��{g���ϋ(Z��EB1�)/���������6U�Ʊ>?���h���yN[�CN���2�e΄t��y����w��n�h]��E2�m��+=���nb�����V��Q���?��,��,�C/g��,K��$���b����J��V:�k�4�	�a������'��X�E��q��C����l��"�=}Gloۤ��s6�&B�2Zk�[��~h"̕��z=��~��ϭ���*m-?��C��d��C�	��`�.��%+��c�[�c,0׷������WN�ۦ��έ���zu�������J�ͪ�['V�<���6ۧ��!�
��ɝ0�V堫cr�����F����Z0D׌��=���L߃����az?���z?2���e�y�#�[ ɸ�k|����� M�8:ɵ��1�%��!3Z^�+E}��l�_��E���IQ^�W��<QS�7�
�NY� ��>we��Z�����
�z�u&�<*��R�xdD�����WS� /f��W�׈K�r�s�����A5�g�Sn!
��f��f��as�]ze����*�˦ࡍ����UZ%����V~B�c�4hw�+r�h^1��C���c={\�<���֦gR8�G7�X!�~@YǑ<˟�&FV��T��b���9M��"�ldM�Ͽݲq���_,���S$w;6R�C�p�^B��<؝�G��}��yzm-9a:~s,� �o��3�+���N\��\���=O�Nd ��2hb�S���S�N�)Y��j�Z�����S4���f��q��ܕ��	��G���X�w���"�"���-��ӊ���UvG.������+�3�- tx)Ltc�`|� ӭp��[pY�����mt����oqb�f��ݰr6��q^�p��厌��	X�LjګHh��Zm�!�p�����.�E�?�Yt��M���!�2�?�T߾vO�W�+����T�h�VمV�K��a�U0�����K}��ؑQ��(� J5�F^�Ec�/2�����Xv���j�A7X1l�c�s���Q���R��Xz��O�ip�-������q��)K�Y hu�6#}ϕG�45Ì�(�|����W=�H����V<��m��{��x�(L��|��P岕.�~�����U�'wd�	hEc�@��[��	�s�q\�~�41' �Ő	���]��������Bk�ّP��<�"Vܟ�:��Z�f�}gS'�Tg,��/15����R�IH�.��=�s\�p]�,��c��?�?N�?[��a)��W\������l�o���e��&�
�����Pd\M�v�\_;y��U:�Ʀ�i�6��S �C��s:�0���fJ�Bh8 �M�n�m"
��A�L�>'?�Lx��~u���ˆ�)�?��}�z��/�[_8rN��ׇ#�Np�2%�2��U1 �ǃ@5q��U8�M�����p�0����ߜn;'y�SC6*��&�$�d}�������������(����Z{<�q��m������ƹ�Ubz���1��H�i�e(�r�n������m���b�NMp�S$
�Y�8�`�Zߝ���9#/謳"� ��)��%��DK��']��83\& 
�g�h��^�nG�A�W����ou�����a�c�;p��CH	4�{}}7௼�h �]uD4��!ьN ����F́@<xi8�@��W�:����""WC�s�\@`�/�F�T���(4<��.��}p}��V¥��c�����z��#��.$��o�Y,����_r��H_�7��̹�?eC;*ر�Ń��?���E������v��/GJ5Á��~��l�2��c��d�
ABJ`E�lo_b���������"�΀S�Ι@���ߺ@����uƿ��o��Z�]���=s�Px1~���?�_�_��������\���^ϟ��5��`���2t_��������^�0�e0��i2�R>��8v�P���s�
��:��7c�C�_�.�Д @�;��I���|���_�|(_�7������c���\����~����(_��o._��o,ߵg�-�����X
=g�8!3����.d��.�$����m�������;.��@����] ���EH/�@���O<7�I�;�V��	�!ڻ:��ㆾ�����9y	�5;�a����Ƞ�<Lc��y����Ϲ@����K�d&`�����!�C�w\����������du>�N$ړ�����1�B�S�BߦP�����S�7a£:�Cx��
�iTG뭦���=�u~�ĳ��6���^N�X�~/c���Y�s�'K��~��U?�ji�h�[��Z\�Z߈��A=D��4N��h��WOG���[�v�[�F��op�z��Hˑ;�?\���p)YQg�r��A8ph�e�7���'q�a}7�� �TY"��T�ǿg���1V�~䮼l��(���ͺu��+��3����7�8Jɬn�1<?j�r�_��6�V)��R�U�Ej=�9�9�)��9�)�9ԜQ�ء�ZXP>`w�'�h{�Yԕ��9K���<b�^9��Y�<�j� �Hz���dG�iO,�K�@YC��k�G����ɗ,P�e�iE3��U�-��/�ǲ?��y}�&�Z���WT`�s�F��bJ�^"YG=�L�G?&��l����3��.������0�L?[��ay��^?�>1p΅�v{��'���?%F�)n�B�YG=��s��{&���"ҋ�
X�S����L/��s\��+*��IP|ܳT[R=��T6�"��l�|�^��j8��-�u�x�����Cl��g���맔�6���r+��6;Xj�3C�eB��:��liJv�x��G[�����PH-)�{�X�\��Ŏ�7�:�:��
�����964��%{���R�����B����m��K���5i?�]��װ$��9���gK��'I�!m�3
'(R�=8��`�"��VJ��VO�KT0@/0z������`��`��hD8�夣*!�}F�f�F�j��1���k���J&���fB&4l��ز�!W����s`��9�
/�%��I�v��
6�k�[e�iL���~ۇ6z;-'{�X����n�+L F��6}d��+�Įc�����aTvd�����z�V��+w/ ݉��@�v����6�5�q�:8촣B�s�`fԖ��dK��	����	���/E�tC��{B��?)��ʽ���R ��G� y��������˴���ep��β��d��?~>"5>���ʏ��n��G��/m�JU@����u���u
���K�lAr�$��xh(@@��w4|��Z�$��-�!m\�{d�N���������GGU?�\���ҵz��ס��r9 C����#Ð,���U���6�G�����z[��qVf*B�3"����6�ILx_+��ݻ���@�V�M+��>Ӳ�\�����)Ү�+=��?�7�'�CKԖ	Ҷ��
W�쭸X��>-i��_�Ba��(�\�;_�7��_�Ú����0�W�,5�ņ�K䤆ӥ@,�"_�=9������Mّ��P���TT�W���g+��Ƥ]���P`Qlz���c��
�gf��Q�8�B|��|�	��QW9�	�ֺ����HvO��o���~K_��*�6�P�%���^�o��qw#����8��uI@V�.���.�& �&@�A���l�J��3J���R�eИHTĊQ�L���\�Oa��N��s�3}��"v�W��<t��p�Z��TD�v+e$`�ɇ�����Vd�@��]�2>�Ҫ.cf�e�0���;m��h��%Y|��n)��@ D����(~II*�v��k�����F�U؋/���CYw'%R�5�����e�Ӥ�1Ґ�@Uu��x�B/?lߟ@Q��^�'�,4iB�$T��ͭ�Dt�	Zg��a̽U��̢�ċ~J�B7Ɗ^�ZJy��Ï�*�ӽo����2t�E<�EN��G�[���� ��̊*61�ؗE��k��N�ɐ�[3m��N�'�5��llQN7-�� *�e��q�h�{"��X
Mm|^`���>��!^s�����Ej�#ߩF�(���M��t��wW��ȗ����%	691�- �p����>��ϓ��h�4Uk9צ��I@q[5�=�Y-�?�L"q�*�=bٴ���0�$�~�v`Aޯ�z?�%
��=��u���������#�XuY�$bQ�����i���FY5-d�Q���jQ:��H�oе3tq���ߨ!k��Kk��q�ڭ)��e����qm�`�%b�g=0��ؾ���"^U�o{�e����*��fVT�k�	����� 	^�t�EV��={Q0QI���������y);�������(^**3+*bY�?3�,�"��������Ǚw晙gf�y���w^c%w�GL4=����R���Q�{b덗�=�x�[�S��hf���!�;�=[�F�V#�s��y�ѣ����cHИh��>!�t��g���c|Z7Kpr�}�3�+�}ձCZ���7��Vj��+]g���_r���.j.ǩ�]��R]7����=��Н0~���D4F_����׆�N\7Js|A
F1�d��OP�|Q���N
�"O������K���W��FW��U���0�����0#��4�c�o߸��) ;��w�������j��c���Z�Y�m�/ܑ�eD�"vg�8}�!����v�}Z3!�S�TX�����Eo��;PVs{YUTԾ�d��ʾ�����/>�����F�N�+��u<|�^�ݛ�,>��F��h�wD�#���i�)�q^c;��\���p*�S,���x�|�֬�ZS���~+��%��7<z��7!�����W��{�?�)��zb�uu}Է��´�T��q����F�w�)g��7�w3�T^9����^���1��Ǜ�z".�4]������?-��V�(��4Gk��fG���\����ɎF�	���4�;-���=��h쐴�N7��6��6�ѩ������*�_���%9F�WTs�+�:�\W˕�>��])��Vw�-bj�^�;
�{Oj{;U�6����?�M��c�n�.�ww���B��է�	%��g1�Eo�%�wV1��n��ћ\���~M�����@HY�7���X]�+������,����<����]��֬a'���Wm�03lÄ�g��3G�q%����k֬�ɔ�a���|e/}�+|��{��^$��`��uUt�jhɼ⪙�$��;^���������ǿ�r�8����C�'�1�s��W���^�e9^���uH):\5��0�����_�$W�D�?y=�>����Uc#k�)����fD�o-q���~rv(�����ߩ2�>�r�wԛI�}�ǫz�m����n3�'R�쓔�����%�&E�}�t��ל���o�5ݰ��TF?w����s·Qk��Y�;Jk�Zg��a�̗Y�i�8�-����c�]9E�O~��'��
J�C���4�s�+�y�_h4F��p���㾺�ae�J��'8�����𺟥��lUTQ|,�۶;,�[h����H���ۢя9��UYmuU$�p8�U%�;4�;#4��~`�l�|ɑ���e��K���[ᰥ�"ߑy��C���[�"_7-j�T����4��0��	5�`vͽB*5��襛H`lm(L����
˯q|&����<��ї�{s���\Eov�W���Ô�A������T���9�q�B��/{i`~�>�m����U��]�@*��]��K�t��=��mRu��-�QS����y����#���v)�*�t�s�]S�N���R�&�uh��>�V���C������L7����P���������:4�u:��ҡ�Z������o2.�����5.C�y�,�zVx�l�NY睲�;e�w�J���)�US�zzU/����O[#��KZ�ґm�����D�V�����vqGh�y���E�D�Т�Qы���!�-y�U��}5����s:B�G�~�K����t�W��t��ab����E������VT]�/3�}{f�Ľƥt:�}�ȼ�����׳��~��#�|ޤ���r�U�v�M�~R����|mF��B�7G?K?�Ա�p�̨z�[�я�a�K��6z�ݠ��(�F��XӃ}p]��ZՂ�������h����%��Dn4nF[�w�uC>S��y�^q�4zw'���Y��Cm��d.���69���ՔsSl��ڏ܍$��ыm�dfD�+�76���ݛ�1��fv�Y�`�
м|ּ�$�f!�����qf��5q􃚝j�p��U��W��������m�t���ڏ���=�˷dT#
u�B��-�_�Yq����t8Z8f�ʸe6� �J�y���F�x�[h����>�8���QEW�Do���܁�%�k�B���w��QW�$�(��ڃ����]�Ⴧ{Paem�V��#�Yԏ�����-(gt���/��`���X�Z=�~�¸RB��Ʈ��Rnܬ��n�Q�]�	`쩣eE?u?��m������0�j�y�5��Մ�o�]����a���5:JJ���=�����oa�.��7��o/*K/���M^Ds�_!��/�Un�"��
w����$����K�l���P��>4�	�����{����������@��n	Jz�FX��X�fotQ�0z`��"z|���vҫSы��j�N�:9��{ح��~Ԭ>KS��5��{�~�ʳ��Wy�x�X���ҏVh{z���h�T�"<�U�-^�!�g�׳��64V��W�5�������u�����ǔ$v��5�.I��W��/yu��ΰ���w�|���Hy�1���)v{A��9���Y�����ÊrV�5&�,�_I|4|x�qEc�:*|�.�V
>���W���7��y*}�G�'ʪ{���GՕ��*�0D��b7x<�i�b�a�_2
o�P߮+��[��O�O���X6��}�+}ɕGsΕU�:�CT2/����ꨲo>�:�9��lvw�*J>�c}�ۗ�J>1��	�|�G��P�#iQ��F����FO�"��+]������󡵷d5?��l4�����6��Y�
gI�d�
�͸/zy:r$7w������C��,��d��eT(}T�����x �;�p�}������E�}d{�ׁ&,2�!^㡢��$�Xˎ�;�5y��S�{���_;d�q9{�>I=c�C��!��[#��h�ӛ2�z_��(��,ot�wx�q�wN�w|����W�7�����w�����g�K<~o`�,���X ���->��s��OdI~��F��`=�g_�W�Q�x�ƊC�ƣ�1�8p�+p8T��3���01+/yYL���	a�j#��繌�r�R\�PLW"}�������E���-I+O�'D�����5�E҃�.�.~��RqY�p���M�'���}�Wq�N�� �_�0-��B�]�RO��d7�Gx7�q90��%	3�H���v�7?�6�M�`�C���ʹ�i+��e5�D_>�;m��O�ҫ6�W^VS�0�4�dQd��_*k�Go�$F���)�+g���9���\��EG���E+���F�&h�AÂ��i��t���/;��^�?z�� �wO^�+�&o��S���[}u%�{֬�f��,��GoM�"ُi��7�>��%_��$��S�^϶����s�D�%z��;��?]���ɓ�EoP����ߣ?۬'�Ç��z�{=U5�y��<��5����IU����ʯ*/�lb����W�8U�Y��D���-�=�J<��K�rL^�[��;v34�ؒ�nU�e���^hM��譑P�P��qע��Wd^MJ"�hvA9�Q帚S���wS��0�rV@9n.����3n6�Ѹ�1��(��,x�p/��k����
<��˄�uG�u���R(Ǩ2�u��Pv�Wxi�.�}pcR-8@�K�����KudixC����ȍto����{4��j��~D�e_�:Zu`�y�t�q#ӑuA:���Ⱥ�u�OLG����3YБ�0��p�#�:���ȟ��!z�6�����5�gz��:=YM�E?�{S����!�����@�B*0�$��K^���e����3�[���HN��ק��kV������l�M
�yQ<�8骋^,�W�t��y�}�Lը��i�?E�oC���)^�W���B�7�b�8v;�O��������ɿ�X�ϽÚ�6������ә��&��PT2
D��l+��n�G�+�Ȧq�/��N�1q�*I��&o��]�K�i�A߹ȼS���k%=�h�@*OS���I�v�ꟲs����5&o�sʂR:a��rN ����&����H��]��a��v=����zc9'�uM¸�
c~�0�u5X�q�J��ƺ���:� �	��(���s���ϲ	�|�	�
RM���M�ŗ�#���G{.@�R���4.+�LQK������@j��6�>?|��S}�������n�Ç
���;����%�?j��=~6
��Ue��۽S�9O%:C|��������|.UN5��ji����D�T�'+K��J&Ex�`Hl).�~�=�vZ�<�o�����h���$�ol�����^�ǢN��J���VI�{�~���D])цi�M��OrLS��P�@o��+>������Jz�c�kN���ŋO>D���%R=�ҳ�K�CLx}A�з�D�-�J�r�[Ɲ/7�b���CO�?���߂T�X�Qy:���L)u����	Y����+jãw\2!�<���]���]T�z:<��UOS�v}
#�����α���hw���@�W�
v	������q��'�P�P�������t�틨�A����a�����QWpe7!��z�|?$X��90n�Fr��>A�Cs��9๭�
�k7������@��T�É�+�A��U^��Q�oq��O�np�������q�?����t�E������F}�����I9������w`c񰻗�;�SƦq��q�	�lCI�S�}���_���`n����'�m��E��vw����/�t:��7�Ar���L�$��Dr-y ��+ܰ����h�v,<@Y��z�W���R��Qw_v���N��;��Q�jo9��-\}�����1b1@+���Y�
"�����{�K�#T9v�ʷ�X���B��[1���ι�Z\�M���עO�;��������е�u�Ch]�U�خ�]��R��<zQ	M�m�pz��R��S�^�E�y��ѷ���|��_�[����b���{�	i��Ôw߾��,�9�~�@�=��1����~���?L�2�goQu���R�lz;*�Q�"��ĨQ!���>��+���������W^C~��3q*f�j�?s"j����آ��>����+t ^�F"��t ^�Nx�`���M=���MEI�uW�ݞ�������}��Ĺ�-��W�&�uW��j`����'I�e�z��φ*��]m1-$K'���X���B�#�눤;�F���}"�}^G����lm���D�'��L������cߕ"�%�;SV�����ԅ�C��*�އ|S#�#"ٍ�_�Iq�;�ԫTM�侻��k��~6L�uG�#}/|�咞�¤;��g@P?�;!���@}J�I�.�j�s����_|�w%=1oDF}���Fx'DF��^"�6��S����K���g�h:�+W���;"�ID�6&wew���������k�@�;Zv�O����~)��_�?�H�W�Bcu�k�^�#��׏�n*�����܈Bj��ۢ��hU�S�jT����=1"����"Fl�wD��<b�¾[�=�$�_���=�t���#��#T�p�.�~{ld�`�.ٗ:�]t�R'\R����͢~���,�I���m�F6T��B����~'N����X�#݁X@$��$ �V �C�9�"��?�#=�X@��@.��3P. �w�h�$`� O/��]�	�{��Y r �	�����R��9�=@��H�/�L 2����E`=�!p8��}�z�}ƻ���v��_�H�%�x��T��r�g���=K�7$��μ�1���ސ�<�#�;x��������!��B2��؉�"nh�qs1+�� �	���o!9Č�$��#�	��KRqmFzKcF
/�k������f��l���8�ge��X	v�$ ��Qd$I���4.��t��
�V�2I�@�Ð։xⳘ?�E����p��̓�a��3X}rpM9��]Z2ǧ���b��@�]P�	~+��L��R����z�f"}BsX}ܭp\��3�\�+�����P�%�Z���O���jic.���,�����}jj.��j/Ԟ�Do?L�����Z�3LV��<�Y�2��c�e��hq�3�vg��fw�9w�e�-v��8����mΤ���V{�,��4�d���[��0��l3�n;��� ����qf��fS&M�vK&�q���69gP6H�=�d�	�N��I��:��6���0�t�ly��6�Eӛ2�m�<AJ��\nsҌ��6Y-���y��W����,� ��4϶�֔���G�L���pZLh��CF2�6��n�f��6E3��r]��	P��A)ڂ���h9AfS�S�-(Ϟ��&V��ʙ���N���s-.�+���X�,�}Ns#5���L���"�fg��岰V�YX?в�6�gF6�N$��P��irZ��[Po�v�ȶX3`-��)XY�72ͮ�Ł�c�9C�ew����3P�;XVZ�Y`w��m���=n8M���0:�DR��$�&�5(/?k�k�rjz2��w��;h���#M@��{�9�n�e��!��1$�'	Cw'��Z��%�0�k��l�n��=�d�0�� �c��M�;��w��m�s4��i3J�ĸ��Cb?�x�-�>'���'�Ǻ����g�z#m\�#b<�&��rǣ�f�=���¸k.��M3�C���X��jy}���ۂa�J�&����ii\�$i#S�]�����#S�C�ȅi�.�6ƜՒ���Ʌ��i�G��rg�	�������<����v�5op�T���2�Qk�p�A�?��8 ̈1�r�D
r�N3�4�`�[�?I�.���lx�wr��$�^A�Ӟ�",�������6C`3��,6�ۂ�?�e�%�ң�)Kf��{fP]�����`�H�\4�C�j�eF�:NNeڳ�����R��A�d;S;$����< ��f�l.��CE��h�&C�n�1���:���Bj��h���]�^������ε�;L�1�n{4�&�eМ؜( �/V�x��L���m698n)���:αد��t��\��6��h:���mq�=��[h,FH�!�j�A߻����ܴ���E���f3�k��iZh����9ׁq��-<V)��:���ŝ�Ĕ�&���C��?Q��my7�˯�Nj��hATR��9*���F�c�o*���Ep��_8�Q�*d�6���F'oPSZeHڦY�ȗ��,(17�:/آYP��I0�K����Nga�L0 �I��ckP<�h1��p�j���p3?�Ŧ$F�M��tI����&�����g���<V��d�H�a��'�I�0~��h�@2!�OJ,P�N�IB���N��T��i���#$ב�_$(H'Io�D�N�~;�.���~���������D�d��� �� ��A�g��
�S�:v���%�k�[���v����w�s�������^���������p��A��Eb�T&W(Uj�V�7��MH4>b䨇��SF�><&-}��&Nzd�G�N3M��4g�ȶ̜eͱ�t�ܞ�sr��>6/����r<����OƦ�Hă����QP�xAa:$������=R\\��
R��ucP��/@{�SRS�[Ղ؂%HE�-��ّ��r�9����'��/6�wc܍#0R��[��_K� ?^;���/�k�_SZ�����~7�i��k	�5����Bx�a��k����f��=�|��*�����m���!��J��¢Eŏ/^�}·��ɧ�=�̟�?���+^x�/����^c���o�{k�����~g��˖��ߺ�?��񎝥e�v���|����𑊣ǎ����S��Ϝ=���_T}���翹�mu���K�}�Cݏ?�|�o�W�����~o��'��P�&�w���������#��uN���j!��$�'��<�Hr���!y��LM&$>�������� )���h�.�7��p7�{fx\nBFy�,�QX[P7�����&g���0�t��o�2٘���i�4O�͇�ty4����iH���qf�XÜ�K��8]����L�����|�vH��]�����(=��44��pq�PD��4�l�0��"8����2�%�N=6�/y���j�0��?x/� �P�<A���R3���qx�H�����9�L�iNu�]�MŇ�cR�I1M$��pJ|
uG�#����4>&-1�s��A�A������zG4<Ja�z�˙1��[`�LwIg�f�&s�[,f��h�Q��ި���pL��X3]y�ɳ]b��&�1�E��� �9ؑ9��Y�>/��	��t���{�*�sy���k;>{�����m�?x���g����ѕo�{!��:�����F{*��/w�����&�ߜi��������ſ�U��#.��b��|�e�Ҡ��1<��^��M�[�W\_~���������������]~E��(ێoP������������J:�S�Մ.ߨ��'k��o�Cm��m\�����v��Im��K/�|>�g�����=(�ӻ�/}���_��g�CB�/�m�����h�o�:��_�1t�6~����{��mo�Ko�����{]��]K��o��_,�Ǯ/_C�kB矹��^:�[o��7B��}��c^�>���B�OΫ��⫡�g�+�_�J���L�^]���H�2tz�K���K���"��b��Q/����+߼"t�1����C��9���\����Y��l���\N����?��G�)t����=:��ӄ?����?���y����$���m���K��>�o_��9�	�_�D���^�7t��K��%��_�8�[]�;�	?�8t����(t�~�6�{ >~a�����0tzo�_:����s~��?������g�G��y��=��X�����ٹ��/��m��o����B��%�I�����A��	ݿW�~�GC��E�3{�n�/�"�[��p�Ϗ	��v�O�=4o#�wnk#�V���2>��x�?X}��ja���ě����ݣ���Q��'��#`�x���o��/\
Okq�[X}��v%��L���s����-��l����A;d�*�wAL��;$���1�{�ɮқ��tI<�� �g�o��_s�r�r�l��X�#L�L�a�0�.���m M+���t��҈�N�ۜ�=�ON�<�Ƙ�<��hh�4w&�!k.�Ҥ�rh���0��e�2�so��	�K�t�sd&!vj��A�I�zPDz��������6�#�ڲ'�����>�l���hڐ�G�F���=3f��Mk��iV��AJ���@֜9Җ�4s����'�ᧉ��'��,��43{M�aIf�l�����(��{m�*k�4����]%�]n�=�� �f��}C���3��%\�� �o�Hr5�\��Zׯ&H��>H�'��l��Ѧ��>W<�I�1�<"�x27�i��ゔ��� =�a�ٙ�jv�Gz��M�[�3ݒ1�����"5�Ն�K���.&��G}*�"C��	���F�G���,$c�Y�@�a�"N>�x��]�i�K�aV�+��2ԓ�evB^�W��{���m��_�-3�a�qUz&|��:�6�b�$kY��!��i�U�� ����6��k���2,)!Y�0P||��/�$P�����䅠ڎf;�h\���@.�$�fOH�����R��om~:���;�k�,���Ȇ>>����\���C�2���u!�i�
&!�J�"XFoH��ʂ�A��)�L{���l�!<�uТ��W�G��@ݟq=x��#=�HG�<����w�n~y�ڗ�2x�?n�lB�w����нI`��� e.���z��%�4KA��˯�i��'.�͓A�+�s��x���\`>t;�a��m!D[l��{�H��4�\���I�r��>|z�.�P��Z��P�ҕ�+ =[|#�{<��<��Fڵ�C<�u�ϴ"�Q��(�����I\{��� ˹�V�A�\�I7,����H�fа
�G8��= R���2���
�n.�@E��T�� ����� n�T��_7�ң,�V��\`�%s�0x8�ox�`���.w^�� X� ~ z}�#)�\`-p���<�v���1`9���;��������z�Х�GT�#�"��[��%�]�	(�N]��0Xl�"��1�
��W�����U��xDLr�7���@�:�x�5�) �G�� V ہo�ȟ����@�	8�<�3�L�o����yDL
�-@����� O ��]�yD	���*�p�u�G��\��� �5� ��@"�00�\�|�<�l>���.�@ǫh`�U��P	'��Hw��Τ�"]I7r���+�Nn#=���r'�!w���=�'���Gz�M�'}H_ҏ��<@bI� @�Ad0B�DD�DB�DF�DA�DE�DC�DG��@�H<
-�H�dNF��dy�$�d�BF�T�0C�H:KƑ�d�H&A�N&Sȣd*���J�`�9d�$�X�L2�XI�]� �ʥo2x�b�`v�#s�cd�'��R@
�BRD�b�8YL�/y���RRB�$OA�>M�!"�ɳ�9(��{�Aԩ�RFNm��k�W�٦�v猩��EN��I����l{�+ݞд��'�/���3��N��ۙl%���馌Y!i�&�4Lԁ�9�9c�ݒ�T�8q�-����t;�k*%d!1���9�2�d�C�l&g}�$�۠n�O7Yǘ��&o6ͺ)iZ.-/g��:�淫���R�7N�zͳ`��,q�J7��4Y%���C�{C���mSE���O����e�T��F-��f	f�-� og;�~�&���t���k0!���X3���.5�K˽�����5q��ru��aʰ���"�{�[��6C!F"�ѽ���	+��������dK,Ih����%�e۝�fo�h:''�*2�l�R�B�����(B�fF����馊2-.�3��4g�#Mq[�d2)lI{�mA�n~�R��c������7�������[��7�o��d��%i'�􅰛��� �v3ʥi'�.� nN�^�	�ͬ?�͹�6��	5	�f��)sL��]��������`�x�e�-t=s�9��P$��q���h�#��X����,� &��-��f�]fw(�m�9�9j���CM[ 2:[/4����9�Yl�`m;�\��=!8lJr���6���O���Y)m�h�i;�I��7�mӷbR�H�
6)BWk&E���
�m�lR��3)�ʨ�Iq��Z�z7Mss�
2)�j��L�6JnähG�`�6��L����Ҥh���&����}�Iq���pʤ�Y�vr�L����I�F�!M���ig�s&E[uiiR�Qnh����Ѯn��r�3'�"6� �-;���{D�ЦZMn�d��&�r��2��pЇD��AT+k�@2�>n[�.�\��,�x����vfZ��iW��m')}[���s8���l�T�b�HxCdf���|���3~��&T�ϦJ΋I������|���]�9��e��৷U�R��D�I/�ʤ~�P�����l.�^5���%�{������-������ff���0�d�ǘ�?>��@�i�,��9vT�E����R����w������������%���@gB��%� ?z:s;��.�����;�i��ϗ������������	��T�1��4�;ޟ�D�V8=gE 8���=Fe�v���y.����E��E�|��Я��_���_ޛ��~���O��c:qm��f7;�����Y8�b�� DC2�+���K���C�\���ݻv&���� ���C�6`%�pӀ$ ���{<�y����V K 7��=��]��[�ہ��*`����w'�b � ��?Z�i�0~����ʩZa~9�k������k���G�?X�x׹ox����>T���GǗ�c��D�T����:�`;��c:\�#�¥z���Ή��஄{\7ܻ�j��7.���>�������;� � .�?b?��d��7.�B�w.��{���*�D�=v�� �;]���Sy��-78��9�������Na��5��ȫ�f~�O�o{�뻅�HO�;!2�-����C��xA���,_��~�_���C�\����_���.���rQ����
t�¼����k�����pn�UTu����]��7μ!�/�:���ﵓ>���#���n���կ?:���1��X(=|��32���3��W~^u��|.�s����%����G����Z@	H!0�@�"��}<~p����	�8�� ��v`���V ���K� ��� 	$J�/t�h�C�Aϳ�b����?:��<hZ�^o�:����GW�#��HMK�����&�s��� :�ߴ���`?�����j�h :2��<@��p����Krx\>4��p��9���E� ǁ� �xC�d�
��џ�4@T�Z^/s�x�p4_W̆\ B'�Y�rA��
�qp�@�v��������G�O��4�_���_F�R�U4����\���������f a����i��1����m�n����\�i���K��=��6;w����?Q��U��t���X2����0;(��*��
�S.9�l�����9���$.���q	Ԃ�[��J6��4�6��l3��g;�sؑ������B_1e�Jwңvc�'�B�!tg���2����_�!����j��Yɖ�QjA��FO4�QJ� �{�D0j\r�Q�����=	��wʯ�9c��<��ۑ��Fz��{��tUid6������r��&D�v���E��:�7�f��hb��$腦,H���N��iZ˃��*-i4���nU��O#��?qlZpZF��"�%�m����)Mke�䳺O"�������".���ӛ��z�=���!|$��Q�l�a�=jlj�a�y0���OX}	�t��$618�NӪ<��t��gmz+9(����0n�)��"�ޒ���n���%�N�����V���g���\�0�='��ʓj��$�\�?]p/XM.�qyޢ�e��gԍ	�n���88O�=�7#�i����Z�oJ�|$��6�ב�p�n�y�Ht���K�{b��iO�)X���w��� ���=�>���l0��Ս^;�v7;��{u.�?�ò]��Ŏ5�f��;�L�2<��lN��Yf�رM�i���-���,fk������co[
������h�=d�AD���:���6�n&
�5�}�.ń-t^AD�9��&|6��3��4�q��ۓ77��iΰ�h�fi��Z�,㑑�_(��k�K&�!�8D�Ȗ8͐[�4t���b��D��9���4g6����^O���ӶG�2͹m�Lx��ҩu4:++�p�f�%h�\�jzA��r�	C�@u��5�l3;-�����	ZϜ˛��1��u�V~�PA�����8`!ے�'!��qQ��O��-~,.������G�F�����w6=�-]ڂ��zNO1�3]�,���8t����<����:�P�����Π��n��u	]�$�=�L�n}����A���y소B�;>~L�Z�2:]�?f�����}3�������©���!��:dT�ȱp��r��H+�Hk���0*ƙ��S,is�%˒����r�/������^�ǌ=F-�s��6�ۙG��GK�f��0�r���s=�e��77�M��Y7��������ه�P�$�	}Ow=$;1��w�l����ը9�kM6�����!f�wH�'�'p׷3��J�t���6A���1l��Pt�{7~%�p�lI $p�@���6��}ܴD.��SF�-QM_�@��8eL�|��E��?KpØ�����g���jR�fẅɟ-gj��	؊��n0LGCy�V�\�`P��w��=\�ڲ�O.Ǧ�5%��I���Cճws8gz�L՞��Y��+m�[�?�/�3�Τ��B2 �&2H`_��҄�Yd�rY&��C�=Lش¾�C���#��)d���;�H]�,����G�'m�G�ob>M�_�q����F=��M����4�$(1~��C�49��v��qSS\�i6����T�~�gqU�7^�k���ARM���II��6̚x����Jڹ{�`n���_l�2�kj�Ͷg4�	��7��$�e+`0�Z���9>�Z��&��ڑ5Ȃ�Wn�A��n��67�,�
�* �Ȼ��H����mq@c8���������{@��[������%2��[�5�O����ܽ�_�܊;����;���;����_����{vO�Խ�c��M��l����[�o�~r�]�Eq|�Գ	�t(���+qWw�J����S�?�۩���#�#{��:g/�ZZS���Z��x��T%WU�n���ϯ��k���'�va�ׇ~�?dQ�c�w�ox���'{~I�}���Wj�5��#F�O߲��Uw}�ưn�;�z
���?"y���o�I��m��wi�o~3E����g&5NY[���4}�R���o�I��~S�W��X�l���|}ߔ�
lI�_z^�Dؘi{�yh�?=��!���ᏺ.��p���25_�.y�ֽ�o������j[��h���h�=�7~�������[��t�X�x�A��>t�7]��䷆]��vش��9�6�7Iz���=;�?{a��=iO�=v�����.W7���冾}ʿ���Fd��5��N,��nڼ�M5��~HI����k���aM�j��{А����3���l�>㱎����)j|�P��/��f�K�n���U.��6��)͹%"�y����׆k��vz����`��=��9+�~�I���w��?�f�������[��j�ĭ���F�$��N{��~OM�X]����_���{��%��?�ݙZtL�C��=�N������������lme�6�~b�9f�g��W��o��؞�n8���]����g�#���F&�a��?ڣ|-7�js��ǌ�ved�sL�A9M5�_)S�\9�g�L�d�]n���_4Xx��[�@��ž����$\:�t�3<N�;������R���P�3̮@dp4�J��j�$f1�Hw�ɅY�>�.�<��zj���,��e�_�"qs�CB��҂W�@�q��Ԟ������đ)�'L�{��k���~��^a��Wa7Q�(U\/�U�MR,yN��t�����|��9�y�xE���3E��7�8�#��yU��9�yu����M_�h�j�zm�n�.K?K���3|o��ݗ���Kq��-ɕ̓HI�H�J�I�KVHVJVIVK�I6J6K�HzK��N�m���?&?#�B�^Q�8��R�WT+.)���k
��PF*�*���eO�@9W�	)���DtN��H/�&!yV�D&-��U�[f�} �(-�)�&'�E�����衈Q�T}���
�B�P*�
��v�n�n�n�n�n�n�n�n�n�n�n�n��T�G�OwHW�;�K�2H�%�?�.~�Ր$���Q�󄛄�F�����Y"�h���WQ�x��Q�Y�T�C�����N� �X2Z�.�#)�<#y@:N:E�Ε>!}OZ&�ZZ-�"���dr�F'/�,3�f��ˊdkd�e�ȶ��*d����$�"�K~���<Vn�'�G��Y�Y��3���+��o�,��Z��計B;<�ڋ
E�"M�Q�U,P,R��X�X�ؠإث�Q|����6�K�K)Wj�S�ӕ3�Ve�r��D�'�z�;ʣʓʳ�*��5%O�Iu���ʨ��JW�R9T�c�gTϫ>P�P�V�S}9�Q��ꨎRR����������o������S��&�;5=5�5��4C5�5ɚL�EcӸ5>�2ͳ�5�j��|�)�Tj>�|���4j"����h�i��ʴIڇ�㴓�.m�6_�P����ڷ���O���o���?j��t�uR�J��%��Mәu3u��ź� kt�ue���#�*�7��:���>Z/���?���׏�Oӛ�3���������k���e���#�*�7��z���!� 0�3<h�77�6L3�3��ņ��k�e���#�*�7�%�^~8G����0Z(�>(��N��3����§���k��e½�#�*�7B���(Z$�=(��M�E3E��Ţ�D�DkD�Ee���#�*�7��"���8Z,�?(��O�l���������������ߊ�K�HzK�%?`t͐n��J�$���ղ��qr�|�|��nE�|�����j��H��v�n��1]�n���4B�éƉ&�"�(W4OT Z$Z"Z*Z&Z.Z���J�Z�N�Q�Y�E��肨Q#�(]$[)[����6�6C�ɶ�Je{d�d�0N�*e�dU���y��A�HE�b�b��h�p���x�������Էj��ѐ��FHN��7�X�~:zq�~��s�o�^�a�a��%Ç�ӆ�/n�Ν�d���4�S�4t����nҁ҇�3�^�:��R�����;��oP|�*�S��ܤ�zN��j���u��]��{4�4ԜԜ�|��}_���S탺�t/�6�~�6�r�BJ^���F�Z��Ǣ;ųŏ�K�ó$�$����T#M��-{\擽,3��Pޣ��S^P�B�kTkUT��/@�����/Y�]�ݠ�X�E?[���D�����r˅��	cE��|��EQ��>�<$�"��Ζ>&-�
d��ɧ�_�S�r�b��}�G�O�Z����[TY�Y�|���?h`D�����\{P��v��Ə��������+�9�KЧ����^4N�$s��{�� ��҃�Ϥ*�Z��ǲ��^�o��.�R�R�+F)�W~��T�G�0�C�)�����(�����~\wAW��M7KRV��^oXk�`����fB���.�٢�D%�g�=����	d�2��%�+{�]�[vM.�Ys���z�'�C���F�JuNՠ�G=X�H]��T�����Q��_+����t?�F�W�w���h����]%	'��~��,/�E4D<ct�x2�i&z�/��J�9����j�&u��b�$Q2B�$I��/)���|-��\��In�L�H��\�<i�t�t�t�t��Jzs�%�R6J���U��r��X�`y��-)PQ�S-V�WVU�����B_��_�������j~�\���q�Y��ީ�x�V�Uk�jGi�h���Z�N�<m�v�v��5�h���]�J���DwLwNW���G����#���О=�5EЕ.��ˆ7oc,1��f\B*��D[������kZ���˄�	_�+�*,��~�$�I�(�,�bE
�^���&*�%�� �K�K�����?��$$� ]�%�0�NH�K.J1�c���j�A:c+]:Ij��ٙ��-WH_�����Q�g�V���]ң�o�?I�H�d�d�ew����2��ə%[,��xP����|Ly@�����z�^�����QjF@;=���Q�f�
�A��>��c���\����~�]��n�H��B��������������c��[Ć$��<C���1�5�~U�b�LW��!����`�|)� ��'��������*D�}�%lŉ⩰#0�-�%QHt��1�d��#��l����h�NҾ�$e�r���U��]�
u%�/�;in�܋Y}0��$j�L�L�,�|�J�[s@�5���ڻ�:�1�O����q��f3<�k����/�.�f u�S�]#�#�
�ra��G�Ӆ����|�B�O�B��p�p?�1��/��Q�%+�}"[�xz�L�B����J��ޭ�E�]}�:^=J��z��E����K�=�j���S�f�����ރ���~��UH)]+I�����o�N�e�*nW߅�z��������U{5oj>���iѮ5�͛똾`����i���G�S��������'���B��CK[�aoQꕩ�ו딇�����?�Ue����OU�c�Y	zRT�)׈�Jm�v�ց���hܫ�C�V�[W�[�{K���[�4}�~��X?֐yy����5�&�Q̃��8>�����¾�7���;D�"�x�x�ۯ�$*�3�3��$��ҿI�eˠ[��K_�?������Q�ҪF��T&�L�[�N��M'UU��Uw�S�EXmt����Ҝ��kfi�h���ت�	�?�^�ަ멻_7@'�tY�^{G�>��E�O!�ɷ�t�菢�	���q8B�a������`���~�V���+�Q~�,WT�f���j��8������h���D7k�����M��V����m�.Zw'����u.��7�#~����w��1�B￡_�ߨ߬?��+
�Ai�������!��i]�����$�@�	,�h���n�9a�x��*v��^�
���7���&�.�v�$�'��F��a	|)������S�5�7h��h;�n��~�u��6�?����Z_�o�7��H*���:�U�hbD}E����h��DJ�<Q�d��>� Y"l�U�#���*�U���+�S�W�F�C
�b��0����.�]Y�y��R��a�����:��B����a6�����`���d�,g��\�jX"��E��G1Z�vX#K�� �*�U���$/K*ek�#�N)R>��R�Z�zSuME��H�1C��.:��R[4�r�
���Bm�v�
=u}t�:'ցoc�w1�c=���l�U�л��뉃��5� �{�c�=aG��b}��xtd�����"��^��O|H\!>�b�ަ\�]�}F��yl����[�@�wk��.9�=��K�/Z�.EG
xd ��~*� �
+�VyY)�H���WV������e<Bw��
'�~]��?,Ɇ�Ɠu���\��)�P|����Y�F�9�E�Ҧj_��z��&��;���>2�4����l1����'�a�}-��t��b ��[�^�V'J���&�$�$��G�"|�j%�a���N��h�4I�l�喡��aנ��f�}��]�]��۠A�S�&�r1��a�]���k������	�\�
�6�	}��2d���#(�zk�a�a�ax�4\���
���s�T��C/�!S�1/l��pBX)�,l���KEJV�>�k�-�m���ˢ�o�X)NGO�Ź��u[��h�^7�{Hb$R���	z�����"�[�RrY� �[B*U��,���H�IOH+�������B�l��-˕-��`��¹,k����ȥr�<]>A����[�t�?��}���w�EբK�:��5G�#�]��˪��C+�'B�$�SY�8�2:���7�e�J�S��R'�3��s���ɗʗ�W�W�7ʷȷ����=!?'?/�$���2M�OQ	�ڠ�TT*�Ze�2Q93V��@����+�-�̳4p�����T�F�ҝ�U�.��$\�}�������W�KH
������$}�>��Fo�~��@�H�D�T�L�+�i�L�*%�.⇑tz�W!��m�R�鉕x_Xa[P��¾H�&	S�$Mf�Ұ
L��	`�.�%J�k%V뫅�����muHX�d�����ja��kB"�E���V����6V4P$d2�4�R�tN�
?S�-�Vҭ��73��.�����LJZ��PҚ|K�h�el$���oofcb��T����=��������������PK
    +Q�HR��%�   $   org/bridj/lib/win64/bridj.dll   $     %�      �|��8>�"!�Xa�E#A��GpAv�FfaW�����XQ#�"��Ml�am|�j[+�������� 	�0���s�������9wfvv�����������f��{�9��{�������9�qf��2ǭ��?7w��zYۋ{���KV�[.�<����y�;��%w?��CAǏ�q�=��A�w�$�;�ꌌN�k�y��9��w.}�3����Y����|Niӟ)���g�s�3�����Azn������A<��r��'�q���ۓԸV�RG��;�-6 #,��m�c�`��S�F���.�䪍TiwMPn��I}t|g���8n����eF�$Td����1\n�^C���A�ڿj���u���{���"�e,�9��q���7����7���+�jD���W30n�j+�_ϖp5W�1@*#����Ǝ��͟Wa��������3�! ܊�[�ڂst��uM������
���&D;�������C.�b�_<��s1�t��D�g��3pBt�3W.ʭ�	^i_;(�0�FIȇ�~B4㶓N:�"��#"w�� vb�P�p�ViF%���B���H�5n���c!�b�A�JP:�J98D+P��~Ѳh0Ҷ�������&$5��<6̞�{:8o�\d�Os�@@����B�'n��iWQ�W���"�8|��ǻ)nTB�?j�KW��b�	�����N�\T��
��⤷|x+�n.x��d�5|��X_Կx�;��c�H�5���Q��)�J�*���� ��m&���l��	6���w����ޞX��m~�) n�Z1�4���.A�����t`�I��2�O��2�t	dvP�|A|Ϲ�F��+�c �/Ά��A�E���"A���-'���u�+j������X�?:�	"6���g��E�>�s�L�������πx0U>Kw-�cw!��s�s���w�|.F�\�ȧ��Mz�gӪ��B�OE�A>��9�>4P�EС�g@�cY>H:m�*�،!r+PA�ʧ/��Y��~�����׹|�OK��I�5�|�J��)�@Կ��'q�(� q��"n�;��m��Y� �7 ѻZ�c?
�VH�����t�|��NM�:l���	��21����d��`?��AC@�.!�󋯑�� C��LP�Q�Ҡy���"�HH�6��[����y���?��"ҏ@�����E��2,E+��/Dn�i�$N��b��	���j���T�����fB���Ί��2���J���:*&�^u5�*;j��Q�-���#���Q��M�0r!�R-����^_��P`(�u�x
�uh<��Jeh�R�Ռ���w�X�m � �[�H&�#T�Hu���;�'^�q�H�ɚ0��^=�_�q*7�&�������B8�b�AAr�a~���{�� o�"��攠i�/��
(��#|E+0�	�t���/������3@_Q�Ƕ�X+���I�W*��|���J�%z�,Kj]�¤+׏��=
�-��z������[g	�x�
��P�"i�9YFY��V�ݑ浝���Y�D����3D;�:D��{4�Z�]���	~+��T���,u�Ja�e�#�P�#�;��'�	�o�t�-P?�yG�f��A?�&/�Cz�u�,?(�2PaБ�����^�*�es��P��\�b��������L7�� ����}C5t��T^�&� �!���=}���
��r<K��ӱ��ϕ�60����\OPOV���2�Ɖ.|��5E�7��q��pd��AU��%��`~0(P� ���e}I���WUc�*ж�piU�a�W�Y���-�0�Vm(�����(Ŕ�1��d刦��	��G�Z1eu�]4�`1����rL��\�ߠ3�$�7
bL�Z�(ޚ�u�w0VՄl�Y�y�(Bۗeǡ�e�<Yz�db�,/���9<�b��=$��Ɩ�n�����8���!%DR/��ݓ�%�ˬh�v���^�T8gA��=^qI����������Sގ5\�@���_χ�bS%d0c����|E�H�E�J u�t�"5u)�6K_<�%둓i)��0"m���,�^	hp�F����@�/�çա�a�19:���T1�.��L���ԙ�j�=�!x�'|�j��t��Ro��rҝ�*��=c��@�4��ĭ�Yz�*��%��+�N�C��}_&;m���z�%a�/Aܔ�<��,�W���V�v�*N���g�=?RN\T��]X�E��k��%��D�5Ўd1�
� tA����mo��6O�+�_|�؋��)�y�^�*��;3�(= n�����) Ke��r�/�į���N�Z�/頗@�O�fc80NLo�l����G�ʽ��q
�6�
���6�R���ɖ	��h�
�8�i���9���gy�b=ﮙPߩ�MW��p��t�O��z,��i� �\C��&���5zp��i�pa^�;��2�t92�> ˥��RA�c0����)��� @I���g=��L��B�$�%�-R@�@:�Lv�;��``X~ϳ�zM�Z�¼���&�z���6+&��i�'����d���Kz����t�u�
�ANo�ݏ8�<!z+c��؝:� H��u(_����ꛂ��+�0�O�y�h�Q���z;��o�I�P
�C���$�\�/1O%���	�����p����I86r��q,��a���I8~Ʊ	�;������#n��qޚ��z�->F�rg��=�+@'J�5��^��"V��˯j���z2����Bq#�_���B=Pw�~���#o�̅������,�K�;#�8�kf�����<M�p�+F�3�M7ԩ�a�3�+�	{q�IC�^��&�~wť���&���`�W������bW�����k�<���'§�'6tOV�����;ZK%����>�U�^AO̴x�gTk�Y�:�d�?��jʘ�)���1��/�5�v�3&�4*�\(/�W��
Cl2�&��%��(�z-}�.��K)����\����*L�֨&o�%�����|f��N�A�L ����]:�l���Z���D2��`��!x��t44�d/�� �F����)aX�!D�&��\iL�o�X������(4����H� Q�X��!���,���#�E��N�a�W=:c��b���iV���Np�=��~�S�=��;ō+A0��/s4��G�[Ƅγ�⤥!l�؇��H�ik2-B�mU
V+��2�	��,�m���}8��ަ1�!����������q��Xs<IU(���8	#��b��QM�2�r��~�sr�7�8�㞅߇`3���`�{~� <����*����|��/���/�]瘒dZ�:A�>�+i����W�<���aJ��c����e頭��ú��%P�����p;X5�ӱ׀Q�8O5j�BD2�l"�64Uv�J&;���zCp6=<=�������43#����do|���;k�����ۡ)�?��	�8�e���HjzF���V=A쏢1���vK��6jZE5Q�8t����-�tc�`�"B(7�ڊ~R���P��P�Nޜ �׉c1#hJz����"53��D1$	E"�\���S��z5�^~�i*��|�Ӱ���<R��%��2�!D�d|���~�/�Q�����Jmb?e1jn#�u��@�$�L��x
v���`Im^%��#JiZ�b8i3j�ϻ�9�Q���5�4;T�%��F"g�1�|~>!K:e�

��S�?�G�����h=Ꮝ"o6��u�	���>�j�b�C��H�;V,�1Yvc&�17ƫ�߉䊪l>k�Dr�Ԡ���C�*���w`M�YP�c9���zD�CfD�}f�Qn���*�^|�F�G�rQQ�w�K�����H¥��1@�9�;�%-9�S����؃��S�`ԓ|LG�ݑ�WU�K�S%�#fF�>��"ލ	Ly��?JS:d{�&��E�On��XG�%�&	�hq�����,��z~U���lZu��,]��2��r�]���'A�����?�ChS�;S�m|E�7�'������bw�<qV�˴�����D���@�T�ZK�^�(��[Lv(��|���96K��	���ej�f��ݭ3rwkF���rh*V�t�9��ٔ[)2�'�w!%�&�����������5��~y��7����ૻ��R�U����.���b������;4�fM�|v���,���RQ��DN�o�#�[������3�,cM�1��u�BxR�C!0�l��������[�X�z�%k�f��u�?���ϒ��ӥ�w�LfF� �.Z[�8>���Rry�NKY�g�J:����I�o,W���=�z/|��W��/������S*�/�����B���0!��������k]��R�g&�W\i�HsfΨ��j�\�q9�8� <������s���/~�]�q_�s<�\�q��9n1�}!����&NT?�G|�$�{§3��G���ھd�����|� v�vZvŲE
9w�F3_�:䐊$Y��D�Z�z�&*:M�+l^2�a�v'�l|2�2 ;�g�p�"�'_�e�p��>���pC��z���U*�W� �AZ�@�iJ	S�H@�|!�A��I�D�L�Fsn%2�7�.��?�]��
��,��Й~g�1o'��4�-�b8����َ}�f�����Q��[�7��א���1b"?���4l�%��O�'1Ah���Z0�on�0.�锋��\8S�����S.��K�x�K=�wN�?���%��֝{�5�
���GĿWb��h���P}��UR���V�ρ�os� ��(�����Ȱ�sRmv�5Q��gw�#b���2d�g�F���֔�d4[�?PL�b�@���N��p����M]sk��R4�����>�i��;�9��vȻq�L�o��F��y��9�y�+��?9�	���P��~������o7��57&�7R�O�kc>\�9�?A+T�x��p���^���0.����|�B�D0�G'�c�oWA��,A`~V)�������?��p���L�H��Q/ i*T	:|�8�_���me� �9�~�:��m>�|��p� �g͓q�Ie[���z� N�t\�"�}O+��\/����W��rH��m��(�%�,��M�Z�>�1��2�߸��AQ.��h���qE7���g��;0�q�� ��V� �^�O��3��M,�����2��Ao�
�A_"�!q�����Il�U���t�a}dx�!iw ����Hxԡ��_��L6�����m��"P�xn��yj7���<t����� �>������Z}D,9A�6��o�&>�.�U,�K9�g�J�i�^�D�nb��zzW$����]��+fY��Ho�F�pW��2����>����8���J/�e�t�w�F����o��N=�_$�[��=�ѳ2z�;��ћ����3M:z7%ѻ�ѻN�w�e9�ԁ�WM*�3Ǻ���y����czzۏ�O���V�,�������,�o��~�D�QF�g�r�噎�������7�e��]�D�Fo�F��e��#���G��7�e���}|TO��(��qT�O��ב�-��vE/�e���D����j�l,�%����y����&�l�ӻ"�^���ql������ԁ޿6i�����Wy�_]�4k �v�A��:�Ů@Vi G�tb����D#�|���ϩ%Wj�W�jh�7?�	7���U�{(�&�c�B�����!���|�)tO&�2w���|�0�*׽K�
����p
�_�����!���5�c'�K�p%���pjy��dpwjpw�p�M�^��&3���d�!���Ĩ}�&�p���F�w�&]���a�q
__ǉ�r�P�`���^+N�"�=�#�o��?�Y�'S=&� +�Ō��)�J/���u��:Jg�1BW���pB?���#�W���D�o
!�����#������O
��CLh�.��	5ǈ���B��Nh���'	������B�p�v���ޑ��PS=jmL&�.]0��j:�%#4���O!��'d�z�#���Vu[S�x�~���:����g�6�����NO(ڑЏ��0Bo�
^8��:B	�����K!���	��;�b�����B�o_]0���u�~֑�Fh9#�F
��N�i=��;Z�%��-M!����'TԑP�z�z(�]8���u�n�H�/�PF��~t�&�	�Hh#4��B��/.�Сm:B���z3B9���Bs/��=�3��9���,�P�����w$�f�2�ީ���&���:B�R�EK�gew�P���@��,�JxTYL��������r��)�:��>q�]I��b���Y�]�M~<C�W=�sVͱ�F��pڦ-�B���3q����+�c\�2z���ˡ[S��F�N��$�ד�&�lGw$�O���l� �ka���8O���FA��0�����!jM.�m�F܉�(�FzŊ�K������:`�E���`j"���X0�NtxDw�/2��-�����s�����rl%� ��1�)3"�^���[��n�bWTa^�_��D'1s��o�d���t~��Y�V+r��a^������n��Ok#�\�3=a-}�k��8�ʩ�W���+{r9�Ci�\S�:R���x�6X�o��j�9���$T�����@a�M�?���X��ӾiVZ�7���s=��*�T��+�h����?yI{�հ3�������7�b�=��R�X܅,Pl7zo��sۡ��T�f���w���)�6�C��Gt�K��������A+�\�7C1?}7?-s)����0�	����n���b���ʹ��I��L_n|(�z/j����ŉ�xOH
	� �>y��5ۙ�/=}V�e{���9_��#S��x��]R�[Y�|��<c��l��\/�&���~�N�$v�Q��l`��c*0���X�tM-�g�l��k��l(�fA^���>�|o�p6��d0l�ɮ�,�-���Ғ�w��}�Q�8�+;���
�
�Q�č�&�q����H���g�xA90��\'�ѯd9�|�2�Zr��O���'�wv����QP*w3٥���R����v*80��%:� �4
�F��$���(��y;���r��.�F�+�_8d���8������u��&�IG!|����n�p~�(�.�e�v\%���!����l� �V��H��҇����]$�b��r=fDA�>�=�ь�u$�~�F�<�#]���������|b� �u�nV�"n�����W�1��ق�sH��ҋ�(��b�4����Q5P,��݈�cj=;�^�f���Ī��Ó��Sᚤ�o'�uL;�t�p
�w�O���X �{���3cF�rz��+�3�X��ǯu04Df;��T'����I��|�1	O�}NW�����$~�8	�ľk�+^����c��ⱚ�E{�qݬ�Rf@���s�z����:���x����H�&�7�&t���L^��k �W��j`��#|�Y>�Nk@�8�jb���8���q�wm^.��<�:_���s}��3���!�=6_�&�o�`�(������ܒ�_GU�.����1������nbt��(��k��۪���6$�=,i�>Քb������:�Au��k�*��E����,��"�2������	�n��#�#��:�V�r�խ�UT}��$�`**�~��|�6 ��\��37���>�����s��,U���g��,S+�,���t�;�Z�+0l��?�N�@v~}��/�������fx�Q�)0�_y%�A;�H!ׄ�E|�N/@�g{h*�ELe: k�:C��V�L��+d�)���)�r=���@��~���2~��MzD?�
S�<����&�h�9�I�c	��y�Iɳ��eYq1A�>|
w��$�H6`�O�ɺL�8��(G�+� �I5@�T�Vk�l��w�"w�F�f�̂��k�!�:�j������5z�9�X�_��8Po�(�G����t5n��9�i��l����� Z��"M>�+�F�����AJ�6�k���2�x��UGe��?���9,��^E�����zM���<l��z&���:j�G��dRw�l���}�o��6+�U��!�XJ��v���ʊ��P�{�ffu�C��� _v@��	�n����P�X��VO�w�Pf��O\-g�ucK����XO{��TS���QmY���י�I������)ͩPu���v�Q�i;tBW��Rޗ���NyoNy�Nyw�������K���ם�|_�C[צ�N25Hw
P�|��L縆��j�eC|��Jz;�$%�x�5(�)�`�f�:�Q<3<Ά�E�C�9pv=Z�{?�\���1���LA�`��V 	}���H�h�[5>�l����\9z6_k�R�b��z����L���h�;叔5H�>Ş�'�����#�ig{����rr<�H6nW����R_�_�I�>�9�Id�R��%����vEs����{R�9�ƙ�4��VU�<��%R��M���RZ�E��Ź�.�N�g+(���V�|b[��
�i>�BKMg
�fd໶�͂,�#������d�w��lfph�J#�GP���Y�Քm��T�A@�]�We�5�����F�e���AӍ.�r��%,���C����j�u�e^��|���R��ph���/�0�!���>1���qzq��kmt�n����_�껪`�)x�4�;�w���L�`#E�6L��v�2��@݇���j�V�1e�F����G�m�/��ۈ�qt���l��l𧋌����us��d=�Ы�M����;��3{�yE�r60��(�v�+�|�(�%�n����ņ~e��ʼS�9���P�Ժ
IEɁ��A�	������^GSNr�U�0&���(�Ӈɽ̪����*&�FW%�n�*�)����Bq�zb�&�K��_�]짛���qW��x"���R&e����Y�M���!��'$��{��ֳ�'RY�R���h'��&BE��"1Uj�sZ��Fvji�JIIqW�/���]q�nӱ��ʄΉ��мb�:@�yG:��s�>�ס�*�u��쬧���.�%DV���i��f��-�j��e�*��e`~^�kBt�*�X���A���VWJ����㨯�'H�}�2�*�B���>l�+����m�L����UĒ��f��4��nL���� ���Am�.��[쨯$VX��?����ʍ��h�C�Ëp8��oec�ۃ��ph�W��l�}7�?��K�G���ݚ2���e�`�p����cܤR�D�7fS&���\�$��]jH�H�]&�T��.�vi� ����k�v�v�z�Z^AA��ˬ@e��\]��Fm�(.��L+N�����%	�2�!�Rt�;�4�� �R�\�H�A8ay<ސ84�31J��b*�����e��o�Y7�ֺyeRZ�6ڣ�)z,���>iv��X�%���+gI���S[Sm�� L�vm��4�+X�i�բimB����6����C|�?��I��2Z
x^W�\se	ӥV�%��2"�m��^VX!��1�߯\˹M��)�VwU^a��4�tJpZIy�w���z�����L
/vΆ��mAw�u$�O�l_v9��B�Y�:����	�g��W�&�ق�~��6Wf�i�,{�:�>�S�/Բ{aѺ���L��A`��e�]��rM��D���R���kT}^�ZQ���a��ߥS��:�RvPӫ�*>Y���riqt+*�/�bR��4�E�hͭ(qh�Y���x�\�k�/�/j���wL�/Wt:;��εۙN�!N�Y�4�."U�?�>_���m���U�;p�����ËZ9\�Ig:~���o��`�f���T��W�Y)
����,��K;(���;W�ɫG�7�Kv���?M W��*�1i�Vl=tu��61��}��{�������]U���о�I��1%�j��Ū=Y���n�@3�b�����EY�H�b�~�:e곥�yH�Oi�~���k�В4%GYJBY��Z}zy��Wt�l`����#�J�%/Ғ�֥�I��'�<�@���R�[�6��~e��h!�T3CT�n�LO�$2E�a�Y�,�B��lp$���@�2{���h튪p��m�ق7t���.����]٪/�l�o0[��:���@�mF�}P��x�.)Uӕ+����XzUս�Q���~�r�de.�]�Ɋ����9�ʫ�T����iX-�+D`�rT�����9���JN�^�)nE��#k�.M�էF�@�-�u��ږܘPm#�}����/H�B�mNW������[b~�`n-�D�����I5I��#;;0HK��]H^	m��o`M��������uj�K�B�Qf���pr� 7"P2����6�Xz>|�����/�w�P-_>CGE{�z��۴�n�u�\�n�|@lV�`g�E��m�F]��un"kr}j�Y	<����g��D�u{���/�ܲ���"�?���Ad����e�����J��D�T�f!�AϥP|=���Iw��oa�Cˡ-W��t�:�̘9�W��p��l\�����r��n���+�;�
x5��Rw~N�w ]*�ȗμ�����T�Np�{|Z����`7",������$G&�݌�l�]�U[Q�I�:p��������4~��EA/>�¯��{� o�&��1��"����i�Jy��x��t�=� ����Z|3j!�R�ϵ��	�G�(��xyP��0bMj���B�������V~e30X��5�~f�H��!};�՞�������Dl���X�B@�Jٟ�&r�~s4��S�r�������/���%�iԬ^q������6r��,�o����ꮑ9�Y˰���4��������ڥ�^^�w��M�9��d_K*���)�r?�,*c�_�����ʗ:eTv�q�&^]dp�{l�P�U<�i��Z;�+�OA5A.n��K�s��>/���Z�I;?��d�����񋔏�,%�A*���qG�z��(�i�>q> \��ɷ,Rˋ�]��[���Ń���X�n�P�˫����@��5j�Kb�'~�#�}�k�������֛ޢ��Ӆ� �%S���02�R-�oYI��W����EPN(�|7�Q� 6�|����D��Q�k�@�e,5�)h��	�� ������hT����%q���䑟m'�zEl�#��G��lG�̦}"�yYV�Ĥ���B"X��M �ұﺍ��I6��:�J`z��.���;�W��D'��u��d�렏)��̲��G@�VH($�\3�%�Rҷ'"�R#�٩����S�Dh@�����M)�m�RU��ߖ�W�-K�o;^�a�۬T���+?�~[��ߊ���~�ϡ��t�V�q[uM��m�Q�bҿ��/�K7�K�҈���N��2U=���=UC��ݿ�!�G?�JяnlA�Ћ�����#�#���OՑ�T��St�z��Yv��#u�Q��-��h��-K�`"�!���(�����t�ˊZ��=j5�~~�z࿣_���#��4�ZK�W�	��_�����e��[Y.M��R�ci����7I
���Ư�-%ـ��q�P��R�QQ)T��c��W�y�Wu�����V�꯿����_�]�gnEw�F��6��J�g�U'L��Rͷ/]�����q�kuj������B�4K���x�,���>h���[7�}S�|ҷ_�N���J��]��,?�a��a~V����*����g�y�gyj������S�g毺�?L���wڟ������6f=����B'���۷��[�ھ���m_!�}�����~`�[�=�7��������_�G�6�w���[��������eaj��?l�O�/�g���p��=0�ʯ�����7��A�(�u��y�Yu�����3��Ez���8�����jY��l M?![fV��f�~��1�im,��jJ��:%��3��Iߎ~N���������w.?�|.O��u��a�sN�|���V�/����\�=����7��s�W������$��(�^���|�h�R�G�X�H���݉��*����ta�.lх���iJ�'똦�t����RP`�P]e+��*0���3�T�	QvG��|�X}����gǒ�Y@lP2�=�P?��@�j��������гF	���鵉���GjDvjD�.��P�?}�}6+!roH�����W�W?�HՏ�>���ǲT��y�Տ+�?�/]���ҫ#����ߜ�_Z��_J=!{�W����oj������[�;�8W���X���WS��)��wv^�V�#he{���^V��*���e��G{Y?�d/k�������5q&Z~�Ԛ"l�?�V�)g����s�ҳ����ɲ�����V!rt�E�I�r��@�çM|�@T����N�yZi���%��A^��)�ƻ��2i�;�ro�1�ǐ)o�l_	�h?�������)9����A�(KB�+(KN#W���N�'����R����V7'�&E�"�Ǚ)U�r�Z�c3�*�~�m��6Ōr�j�l��Ǖ/���Bx����������,��b��2�%�_?Eۡ6��<��Wģb� ��	��VK�W]�֍n��o�C��+M��Ͻ��4�u�?��S�q�l�����'y�S�����e_Xw�K�C��]R�4"�YS�]@�Gpy���^U6���|lKt�9(忩9&��j �Q�1��"�5�ar�%����lx�Ք���.��?�C�3�5�W.���`x�`j���<��R%�Y����~�X���L����Uꏰx]��cG�72�NgW+��FL�Ó���Y(��
፹B}m/��3ǅ?B��6�m����~1�_�g��_S����쑋��%�r�9-�:��S&���Əg��Blm��N���v����xy8�<
�^?D}����|MG-�Mo�yP�qY~q��/�����V��/��(�xX��B�`��s�.w9�k��F�/Y��ݶR���lJ�3�St�D����=z�	�a7�}P�����E�+� ��(���P�LB�ى'�~�ԟ@��b�]O��$]� r��'��S@�r!L�K���ӳC�
�/�<�����}"!��;�8� ��3a���+�6����te�4���2��Z[��ZY��	���X������������±���PibC5p��㰳6�E��#�1�%u��V���uw�ޅݥ���Z�&�Ǥ,)�EF�?:�s�%J:v1� �3�	�R�]�E�����ьo'c�1�F�VW�`�\�35�ۯ�w,�9n�|�����z��W#��S�<��5u�[k�����mh`�3��;\�,�klt#��E������tE7�DL�u2o �U��e
;b�G�l�V]��'bTu�_�4)�
D@���-p@5�"��}0G��I/%}Rt��etӃe"�[O;λ�y�O�q��	���ȣ���v_�:${�LR:Dz\����
IK!��A��;j�D�
��/��~��&Ϻ:�o�ҝ#��
�ܵ] ��K�_i�a.�
��}�y'^��Ym6�Rꍼ�$���������J���?a]�d�>���
�Ⱦ:��o�)��bפ���~�&Ko�R���,����/Z!9�x�w{��#!��tA���Rn���c���. ݇���[�~�Uj���J��
�݇;���Z�����,��}���U�[ϕ�ۧ��R^��\�·^3
r]�h��З>PZ9q!|����w���x�\�ie���iB�ʮꂩ�zSq��uŝ�U%>��Q��ti�����Ǐ)��a{����<�73���	�������4F�נY,���f�z�K�B�"��� =k�H�>�
�B^ΐ�?Q����I |[�[z,n�JR�Ot��1�s���n��؅O����]7�(i�U�~!�E�Y�� i��Ş�A�8���ۈ�-E��wEuc�渎œ]���6��n��נ[�?��R�6pm�����d�}��/�؟� E�u���'�-*�q�$��?/��OЕ�殀�㩤mGu%��
x$��c>�U��� =�w�Y/���Ҫ {V�v8i��0궛B}�B��`j��S2Chs��J�����8:�[�����5'�Kd����N�]�������fP��Z��`��}n��0�������}��k]�D�e	��Qr4���_�_|���"-�W�}ǝt/쉧=/�������!D�Y�Q�Y��t� *�'<x�Ӡi��ƾ���A��,��.Ñ}8j�m�淡����ntXs�]�]�o~���l��;`�n�λ��6-xc[�!�����On�2rm[�1ȗ��������j��e�s g1Kh"��Ns��>�1��H�;�������� B��Y����A������@[�����0��:���?2Ko�V�m��YO+D��v�!��������%��1��Q��Y�|���[XR�.0`㰰$���T?==?_�~�~��ÆQY��a\�90.�rc���0�1&7`l+ƶ���-���oI;>�02�Z����֜#vS��j��!���Qm#j Ou�Dqf���*J4P8f�:��3$(�5�#q����ю%n��@Y�6������x��Hfh5�|9���>���kh�r}3���յ�_���ێ�ۊq�a#�$�;�q-�|Qa�M�a<q��9���g-z0*�7Mb�n�b�({��`�b8�~�8�Z)��$�D�A���|[umt�i�§<��Cr�T6
|�)@��	��C��h�FU7#B2��b��8�8j�z$�G���z���g���IzyM�2�oI?F깞��č���#�p/���Ԩ��	})�(�7@Ȍ7�>e��\t��F�&���@j0���3����j�Y���0Pf�+L����J��<�p�)������{f�3��Q�%��-���Z0qדC0Rd�G� P�c�Teͥ���e�x���1佟6������z�A��D�.vK���"-�%��4f���
�r��0&������6Z���h1I �@l�*��P������$|?��)^��7y\��vɻlM�ݚD�����	�»8�x��ޑ����{�]��:�}�]��O%���X��F�0"#w��㟯�S�l	�6��7Iӆ������)��ޥ�!!���d�į��d��%��G�� l)@�GӤ�`�ś��>|_8Dn�@?��/�c�l�;d���̾_��*w�F���C��L���0��D�}�}�"�H�4��Z(=Y��@F:����OCwH#!bm��,�U�(_1Љ9���O~�IM ���vH�=�X?���x+��x?��w�;J"|��(��S��R�O�}t�e��Y�Ol?�	
ď�o�X�[Ж9mZ��\��q���y��̅w��U���n���,��x�ԣ�p}
ҎI����.��4���f)+��>�ːs�rqQ�LW<�G�j	g
ݤa=vV�O�l�l�x
k�Ym�Řkߦ��͌�X7&9`�X�[<�.E'��v��%�"M�cI����{�����;l�d�|�ϰ-7`[�	m�����}��@G�˙��ɕk{��X��%VZ&Ü%d�xw*.X\hi�(��we�*˸
��K��F識�F�!{�`��q�q�!�q�	��fW�	�V�׎]ܱС-1����lC�x0 Jҥ �x�����I�Bä�����(�����W��)p�Sa�������&��|b�穫�hin���4x«�$5<>�����-kq�G��Tv&=7���nA�4~�Y�B�Z�O���=��r�����U!Kx�1��9�n,��U��x n�+|,��1����ܠ������宅��rW1� ��=���R�`e!t�7BY *\��e�1 �7��v����<���B�w�������?����xN֘��ã��`������N	�6z\���o�z\��]2�6-ފ���r~�7��||�<9~�����)��y��	��o�b�o�fqc��1h]�Cu�#Pe�+\g\&퉣���?�k	o���6:�m-��Mg��}�`O����>`��=��Y�H�5�p� �{!}��ը�E�#���>H�
�ﻎm?�>�2�ew!���t�W��x% ��:��ô�����><�br�����bq�tπ�����8�i�0�s.��k���iU����!7;��,��#:��w��ӵ����4q��e��8iS^�#ϖS�,d�S"�:Z�Qo����z˯!������<!�Bf��fd�@x�.���s\�b�|lX�7�}���T��������!���`p�`B�")Al��3�Ӥ����
��JP�8�.9�g`�+��4�<�X�Spn9�Y���kM�K�;V!�G#Z��Y����9(��t�3L�PI�sl�:�w�Dh�
����}�HM쀺�C������?��|�ڴ�"�R�3H��D"�#����~d���}�>�{�pl�
Fi�d�b�^��V�>�-������F���[��F��OEKs����(5^��+��q�������'a����L����sl׉[9.d#���^�Q����9��8)�8o�2Hǿ��w;��"Y�5hQ�X�;��f��� �T�&��	v�Cx�s��L�MD��"���������L8ނ�K���'�#,��3p�6�>�x��+^�麸�<�����g]gC]}ĺ�qJ%�T��,���m�fL�������p��H����I?�0���c�x\gB5�j�q���k�h!�x`�S��&�W􁋡����} q�;����8pq��:��<\@��C���y��x/m���.��ak?b�����!ۛ %��:
�$.��&Lfyt�N��/j��^�d4s�g���%��1�q	v���KN����Z�&�\������0ƴ�9�����y�4J��K�O��)��k"	S�(�CZ 0����)<���{p�� (��.��}��8X,2��gU�ߌTl�q��mg4�e�՟$l�4�5����E�Y��-�$�`������7��T�� �m���M��F�[��|vy����/���[1{�fos�� �V��z������7�&���:Da�h`�D��� � ���Ǔ��Dfx�
����r�"Ȳ܃U�ѐ���2�fw�ڌ�3j3sp'�4���5*�'���/��5����8@�5���U�&�o�}u��v3<.&�N�/��l6w}"��-K�92ȠU��%`Y�����`�|���������ᜠ��g���&'׊�7+rria�7�4I�� �n-���	�E�u�Z�܀؂���؟!���X���oU����걟u���&t�z;�J>�
ey�2��:O��'��=���Δ������/�����^�D�	�to�7S�D�E���Ck*
?��L�N������iF%���]M�+�rȘ��Vw���0m�cx���U������LcH�6�]�K P��Zih�ƭQ3�\��^ȧ]��Not�����:,u�-�jX��ܪ,z2ے��I.��	�PJgY�UY�L��"`#�bZ���9��h�9u����,�j����.ҽ�tk2��͘ �4��xf ��;8%o���Zu3.��Bx������6�-����@I��d�ߴ](i�_��WR7N�k�i�`L�m�ɯ���Z����&��HR;�Z���$z�?H�.Ep�����(z�p`��4�4�F��d��^��9��*�ǯ�N����I6/L����4�U�ł���G�������xZx|�#�u�-\b�p]�ˑ���`Z���&݀k��`���N���%Y��۱'��N�e�����T��>dߊ�����6��zţ�y_�Eo3H�T�:O���z\�.����O�X�|���7.<R�?�j���d���@�=e&�g�l��=�6$��	�3��J#dZ�	���@�XS�~ dڤ,��{OҚ�h�-a�{��r=2{��R�9�9d9��-�b���|��R��ݢD%����H!1�$�x�.:f"ߚN����� ;�Ȇ�B�Ox�b�J����.}����/�;��t��U%�h!tΒ>4�ۤ1�Б�W6hO�y�6ɇ��V���0��S a�6��Lw=u���������-O�zpm�@v��6|�񇍡c��؋��Q������WA��B�v���8˷�Cc�>�s��|Q�9aX'O,�B��e�M-�:'�t�s����w�rܒ����m�<m���~�3�=�~�FBtΉ_�w}r�]�%J�.[�-�������ϲ���v Ad���:R��ZUlا���w�`�9O��8DKs���ۗc�������x�/��D,�ywaZ���>��!���՘���Jb����_��vc_�^��KzB8n��a���_���~9 F�Tp�~���j�-�C|�y�p#���_��L��炖 ���h0�l�Ӡ�^b���SMP�壖݃:�"=p��l�G_ ͎݃�~K�hF�uh�w3T��F�<r5n^]�֛�o���]8yH�=m�,��FG��6)�&~��Y|���+��f�}����c�c|��&������m4�*�[�܅kӼ���Go�p�#9�ڇ�x!g�����Tf~#@����̿ئ��x�����">�1@b�T�oh�d�Y���`�!!��6��r�5d'<hF�t 3�B�@3���nU�{tM�e�/��#^45Ѓ��C�r��f�Y����d�R����[�u{���;����΃�7I3�a#׃8�x4������������+[XI�CM/ڍ�d��J�Yl����D��
��M��`+1��G�j_X�ұ�F�U�I�hB�F�[g\��я�	pԞ��\���r��Qޮ�%��:R�Qw�}��`�t<���� �؊�ߌ�M�=ݶ�Oj?�Ez���Џ�=~��!���N-0�x�{uV��GЍ��tp
Ïr�5z�EF�~�CmePWV�_���Y��nP��'^�է��VТ�Q���gp�k�}7��y��6A�r/_��&��>��&^�+���
K\�����o2�a��g_W��+;��:7��4AG����0b� ��h��"��3���3�E���x-�׋���:��]R��%A�\���H����Z�QxH��d8j�%�z�ހ�j���`��˜��[6�b�ၮb��y�+$ۤ������_5�Z��0�1(���	44�!�>,ɼ�1��4���4�&����l&��d�,���m���<�q�;�=��LE����տh�؟k�4[0#s��٣{���>R
�j�`��r��B�ؠ� mW��&n2�ݡJ(�[�)P��)`�+~Ns0>�-8����Ԇ�K�IC��q6�oG�gt�w��3c<h����(mK����4K�������!i�آ���O��jr���%��`4q�9�Ժ�F�f���yR��|���ѻ�q�3>Ȯ�Idߘ�#+=t�_�����8\�;��L�A��x�
�+����l��҃������~<��v`�����1��0�x��W\����ĿK�,�PL!f4���ѽ!Zj!ljpml�P�I05
�˘�`��u8�3^��G����d����7=�!v��P����{�w�-x�i�k��m�C���@Ӽ⎭}��:���O�{�Q�<xL�_<*:�>(��#..�3��f���n3�47�{,������6+�%����|j��!N}�n�
�d�\59��%����i�VJ�DI~�%Ƿ��G�c�J��ql���Mg��/�?2h����S}`������q��13��%~�ؙ��r��a��*]Dt�a��H�fy7>�B�.9'����':�[@�wTZ�FC����=~`J���><�ij��xj��@�!=CI�-����i�@Č��@!?�$�xK@��@�K�e��e�Q��V���A�:�	s��)���!��O�����O�FGPl�P6,�Y�K�:ܣ�(��#ȵ~W�#=��m��~��t�=�̮s�
ڢ��ct��RO�xr?�!֟l�ç�/�V^75n����n��05F j����?� a��4P�M��S�H6����`ں�
����µF��Z�\[wOY�@߉'|�G�We���q��B3Ei�9e�/a���ɬ���m�^��qh`^M|��-Ȁ��~�P_!}��C���ɒ_��M9V���Rψ�`,6�����jr�]�3��uF,#����DP_Ư���A�D���6Cj>��+UO_:&�x�9h���{C�s��޸�ƥ�AR�������zc�p�%�����Z�e�Zм��2C{��]G.�/��:K�����|�S5�c�Z�x2�ޢu�����*��s�x4a{� 7$٨P~�����jE=��ˢ^�EJQKG����5�Q��n���@�*քl�)���}�@6��6���yh��I�u�؝]3���ڠQ��1��X�Y�e7�����ٜ/��q!���g�O�B�D7�����E2����eRSS��8����B�O9�k�Z��Z--k{������K��+�q2f�	ܼ��$v	�u�A�DIx�_�0$�LW.vf�Q�������
�O����]�`�\�����]4�(���;�NFG+�Z�E>G3���"2�����8�+~M�����}M�I�&Ŷ��]ҋ��7��i���h�|ʡ���S4�!ȵ�j'M{2�5����W��v��AB�� �;pa�#�
�x�J��i��]�y|��h��)�wr�K��u@Y�[�d ~�F
��␚�@K��"�L5D�F�4�+�5��>؂G�l�~�t=�ʖ�?|�q���h��p�d�`����J�G�&�2̸�]�������u@Z-������4S�k���u�<x���g��/�r����Yz�2��~Ͷ�d�\a�T�E��/DH�L�idG;���u� m]��2�N�&�Q0�/��r�n�K�Qm�_�)�0����<��IZ5���)��]����Vg���^��"3��3r��a�L���]>S=r�W�����{�<ƕ��@(���]8���!����˂�1��C�8��Q�j�mR�8L��-N2J���>��t҃>���u�C]n�.l���\���I����>�QG�_�<����X6q�	���[X���(�N��)���y�
͎�5a��r�/c�B,������t�B=L����tgs]=o1��ٹ>�~x����;m�w@�=��ZE�?낯�J��hq�krW}*��t)���1�1�24�ɂ,:CQ��axR���y��A�(��GS�38���:h�_�D�D
��k��O�y�������`�J_2>˘�(K՜�e���} ���\W~폳z
�'���N�̘%%Y2���%NP�����ƥ����dAM��A�S�xd.�OZ��M��9J]�!K8]�eu�x���������h�(�*�v���M�/A£堹r�_�~�>�ǔ����F�RA����X4d�G��*�$�:W�:|x�h�H�@5��ѴJ�@R�C�}��s.ع���5t��2n�v�t��mD߃3�9�J�^���8� (J��K�x�~��+مˡ;|�OBi�z�ӥ��F*-�+���e�����e�6:�������tp��_u�G<����B����*ZZ����8֝�����b����4x�w��z��uLP>^�/]�`^�/���@�?b5�D��?�[��q�G�$����G�6Q���?�k�=mFf��<�|��#��u`w%�U�yBܧ����4<�l�+�
+kf�d���E�Gf�	Wb=|��������B��]
��+�F�I|��ۋ���F�(xQ��n���QT��2��4_���s���o��~���U�:�?�!�ٽ;_��<oκ��^�5�;�����axcQR����#6IBZ��f�ܓr��!�']�C<ᳲG<��yo;��THl���%�{� ��uZ�?�����&�QT��pw�;�lT��&A�F#�KBØ
�Z	�4�8��@��1@bu4����љqƙ7���!�B:!{ � .A\�)Q@���snu��Y�{������#��޺��]�=�ܳ9#����!x!�R�T3͵�z�7�Spv���bh$5\ȝ�����dgc�e�k�/�<B�m�/3k<����N|�́������R�Y-��'��B����=%If�v�[8�p�{��n�*Kk�R�Cľx�~]����Jt}�eiG��e�\��E�����>�
�� %5�g_��O8I=h���R�I��]+8_ �^�+Y��=x�_��0䬓8�9�M�O�����-rR<�0�o���M���8�.Js��s��܊۟߈Iy���[*��%����S8�wj�x��{��k?r+��0��t���|���p ?��k����<����p���cz�p(z`F���LZ_�V�6�XT��y)���zC�v��� ?J�-(��ե��E���8wg��Nu�c��-.���<��οK�G�x���S�9*�9	�0����#��� ���ѵ�n޹c��ƣ�~��F�I���YrW��KS5���>��Ղn�q��hC<�7'�#���r�p�����;a��cBv�1Na��z�A�v�����.�bn�)�G���.�����9!����&�㫧��w"
V�W}9V�"�q�Ҧtj�����n����$�����rN,鈸{]Ԇ81���k��5�76�����j��V�|v]�W�M���Π$/�j�	T��4��:I����l31ۙ�����8�q8��.	@Sb��0����u�kցY�j3�� �	K�����%VAx���d�B<H�2�2��I�a�P䥉������]�ZU{�`�
إ1�zS(��,vfc�':��������Y^� �c@f HT�{�W��-i�Sp��dŎۀ�P�[�u�s�r�5�Z:��{t��<m��i�C����Ɋ��A�򋰩�X�Դަ� r�@V�gꂆ�<7n�b�ӂ}g/��8�Y���v��]n�#w-��۸��P4E�ʸ���=������\��x��T��Зx�v��  t�X@XU*_w�wD��&�*�m��ЛX�|]6{se��i.�<���c�47��)�?[���1���E`�RB	$�4
��Z���3�y/M�	�u 8��]���b��R^>w�7å\�;�z	��60���n��!t�73���X*����9�_C۱�T' Oq�:� ���N���ن�N���@RV�VJ�Ml�xg�t��5Q�ܘɦh���,��6x�w۵۠Rm��۬͂��yw�vk���e�(�G!> x�.n����
ٽ��7g�ѺRA��0��Ka
9OGpG��h4a"����A-S�v�H�1�~�ك���v}e���TL���5;�e��t)	�y���^ȫ1腼������Vd�D�"��7"�p��~-���ׯ_G<#h��A0 ��J[�v!�P�tZ!�d�����|���P�KKݶ=�Pp�N(���Ǆ��8�{����y�@���:W��d��^I��9)f�
�!w�H=%u����VZx�}��,�+*���O�1i	��A�5�K��Xz�X�**��g�Q�F\���my:��:�s*$^}p��}�˞���+͡�q(��ِWsE���E��ӎq�c��t�7��7��kD�@���}zQ�0��Ҙ�mYk?�[���z:����țy�p�A�T�I�+�-���p�p��X�����k[�{�'WiSc�6yaҦ�d�6S¤�$F�HY�9��I1d�B�� #�D�\�k.�M�'E�b�����r#IB���O�ND�I�ͦ�I�6��mDؠ�׉ne!��N^i��� ~�8�؍ь�	W�8��È"
�2���ޒ�倜t�Q�:�
���GbgTZD�p���>0�}F��7T`a@�.��1��w"x*��W����nAd0�$Lh�]x��r����d��x�����8M<e/��E�+������K�y���Pq\�P�t�Nq_�6FGd�P-Aor�J C���d�N BH��9���u��(fą�����ֹMB�') �
��P�6í���W[�{I���p�nK��+hLCKq�a�"���+�[�?I+
�դM�Y�:F��.F\���Ҁ�pq��x2v .�mvVqUl�� 9'
�j��N��;@ȿ )+6���}��W����q�6 qa�-͌�hE���"�H�~<�f8YD\T8�8_"���N^5Y�B�,�ɫ8��7�k4���A
`��|`K�X8�c@b!�߂Y���\=�L�	@�|4�0}W?BA�/t9��
Ao"�V��s���	"\P���ξ��>L'�����pN��ir�+2����E\�l#�̩8p�q�'�|ul3K�d��	�6Rc$ʒ������|<GgJ�Bf'�O���ٍp䦩�E�L=����j�.@��>�ԗ� T-d�����ή�?M@� �\K�_��]ߋB���v��J�i�޹_��;MXK�է:��s��'j�6�~�LB)CmT�EhW�נ�u֗�&A�}�y���D�菻E�}���'b|$hX��p��A���p�U�w�S|�����;���7:�{��D�{�@��4x.�2�TJ�g����ړ�-�&�)
�$� �#T�lyU��#X5H��5櫼C���I�9�zz6�_I��]����ɉ� r/�_ ��� �����q��]��	���-�S�y�^u�Y�&iB/E��:	(hu޴o8_��Ɯ�=�z{�w�K�Ҷ����d��z~g���-$�5��ޜ
y���tdT�|.p{��a>�Xޠ懦��iω�T�Q�.B�ui8�sU��{�3�
Ų�9ty!0�q���SRL��y���(��|"w\�g�v�7A����j�H���FhRӞ�u0]���2@�W�z��i�7�v���жn�"B��4�0��d�\ٺ���d�����U3Q�q�?��m�D`i[1�U���-'�|������$HȁHn<�aJ!�x�rC���F^ޠ$�8u���aLa�,�os>'1'[Œ,���f����'���s'@έ'p���f���T#�r���[{���l��^��;��oZ����|EIN��-w+֞�f7*�;�2X�Άr,�q�jqИ[�k��;?]�Z��KK��#-�;\&�t'��Qqr����3����|������K>�=�@,���d�W��a��^�ж�a�,���.I�Yz�d�/֚�γ叺�UG�vK��q�j��ԑ"t�H���ښ���J6�ސ��ka��.�W�Т���Qû�Y8�.�N{�%��kE6��͘amyZ<ZT�B�.fm}�0?g�g&i���y�f����6t.�n�\2�ã8A���,��`�3A�"í<�U���D���:�@�{ŉ��׊��qִq�$�� �8��c�/�s��ؤ�ή埈J��t=^FMD�� �0�4���>��r0yƪ|�M��8��
3�W����A���R�N�|2��b����_n0�N�XҢ�7D�m�_��1�7j�p��EX�
�+�3���L��M��w��\=�c��d��}<�~D�`�V�j�],i-mP����?Ma� %o��I�N!y�KLͶJ�	"���D����y�ҘI���(!_��dŞ�!K�3 ��f3��j��Ai�m���΋�C�몎筿�{�E�ry�EZ�q5��8XK��l|�G�e�����m��CSu������4)����a���t���gv��;j±NC#!�^�8I�;M(��dw���c�x=�&"{����`�s�ԁM�Ʒ�;��C"f�+r.�j�6-g������҆�����Mq�&Wm�j�<�9U^��4����L�k�--jr�����7P߰��M-�pX@�!��@o݆����=4���|.��rz:��?���F�ֆ��D\���:��'����W��ш��&ۗא(��_��X�6�3F�F�gA0��<���kQ<A}�J����+�/:O�X ��_
�[_1���s�r��'me;���	XO���|�Z�1㎩�`��:�?n6�	��(w�(l�a0�yJr<�Е��[��H�@;��^����E�0�Eۤ�fۑ����&���+ԅ>p��HPa�?���b�D��G�=eI�<�a���,��a���x;ÁoPa2Yb�Yq��h�9{;ތe��=eVZ��ί%�Fǻ$a����[��
����0E����|�7���ב��=Y�|�lZ��¹G���sU����p�i��IQ��_o��{"�A�KN`��Sc���C�b*�t2*E�]Z�_�����˩�fc������B�dv�>�"���>G�Lo%�^Et��ަr_�������)����SJ�ڳq��4"���&��O��!��i�p$��z����塈,?FWX!�ŭp;p��ds%�^�u�Vs�]6o�����MbIf��]@���7�G�e���\�J�H)�v(ɳ͈5�(Pv(z����L�^��s��<s�ƙQFr�X9�	��Nٌ4�7�Y�_d�kUN�c�.�V�i�TN�yT
>i7VN{**�
ӦUND��=.���iOF��Ԁ6�r�/0-���`��qYx��O�L��O:�C ��_gԢ$ �8�r��XD�:<˶�]����e�^��O'?�i"��$��f�� �/��1�8>��ǵ���)�>�^���s�	w=����x`�2x)���l�s�Nh���͂��;@H�
����J�m�����i��$km�WI��B�r��ٱ<��A�/���J���+u�Z<_c�\�Q���=%㠦M�j��d���]O��|�9�_3����ф8c�/����ۊ�d���j3V��_3̄���e�1 P�zg���5B�-MB��44yx�v)��V3����e#��V�V��2�oz#M�F\ݚ8��(�'��#$<���r�UPv2S��ȍ3��)�#�L�O�%���0�!'mdR &s� �u;��ߺb�"1���t}o�Z}>/R��������T����!?�#��O�(Z]�#��5U2cU0��bP�ֻU�m�8� 5��Qev�/���&� 6�
���G�����7#ςf({�z�otB�qm���1��z7�����|�b�Ef�	U��C��'�|ɧCHq�����C���A$���'d��	X��Ιz������M�s<N�ۛ&f�+���b4�� �B֤f��o4bɆ(%{�W�C]Q4n�_}�U]�'���l�wR�-v
;���i���c��Qk֎�Ϟ�k�}49�s=��ޓϞ�@�7��Vg�S��fVI3q��UȌH��wY�2��m����O�n���t9��x����z(�|)L~WGYQ��J#����|� �в�m��(�n��P����++�Z�(܅�1��)qO�R
����
���BԇO��&J�q,��"TQ�0�_m�ߙ$�6�=F�W��.�Y�~�49��,ep�s�����]����v4�"�궼����=�R=9��b��7�>���l�wʍ���`[Hr�*��Cɒɪ4h�k�� ?��L��Z��Sj�B�}��/�k��@��v �ۈ�G�o�v�qS.G�=L���=��	K��w4J��7�}A@8�~k��Tij�mf�rn�Pn=ov��!��q|������͘Z`��l}������u�u��G��y7��U~�}ÖJ��V)U�6YJB�W�7��mf}������vg������R��q�J��G}��q\�g�!���`?�+�xD.5�S��yKH	(�x+����0J�A&~��N٫n9�w�s���=���iȦ]�&iȢ�E3���g�6m�k)�_�u��?^٥2�!�O�)��X�Y��6"������>D}�?଎��'� ���嶘;#Ú\*�v�^�E�7�0P�,��2��ͺ��v��E�$�-��'`��{t��m�(�d�A���$>153��&�i����gp��� �����W�̅g��L(��V��_5Z,�[��g'�*>g6L�h���<K��t�P ���e���o�i�q�β�N��@&^�_#�$��T�W�}>�ԪٲaX��Q*��IU�U�D����<�S����<*힄g�m��g��B�ۤ�̠�:�x��b �;�t�A��(�!��-瘼DEI����H9����Y����S�%�o��Q9�L�X�����_RX�2>v~,^�`B%Q�򋐴��|�^u!K�+Q��ȢX����x	��&�g������]�gR[0�������%d��e]�'��S8�K�Ŧ�'k��$T�أ��7�i�[��dl?�o���_�	p�U�G��N�ʴ~��~�>� _Į]�@ʳ��-��A��@��(��6Rh�J�K#U2 �+��'�
3��hO�.����	�ߧ���ާ�,��/��'��S�?h�`N�A#)�#su1-�`�����?ݣ�8�KW����^@�x9ލ��J��>���nĽ[a7�!���db��W�N�.��\	%���3D���?�Q-��Z�҆�O�L�JJ̇z3]�24Z���s�0���>|s_bI�r�<N��Vu�� ��2�gq�����W�HQ���`}8�F�N���q�����X/���U�E7Wy����ɗ�4�I�2k�1����)U�A�g��x��
?�0k�J�b�5���~�Ҿ�#�1$�0b�V�6}��F@������eX����k�<�w ��=L��?��+�<n�~�F���ͽ���_(v���I��̠�w���| �_��b��,G���+�u�`gߣM��ꡆw��W�� �tE����9ׁ�������\�N�苢M{��������F���A��k>N��)��y��t2#��n�FV��H䷋�'�0^���|j �BZso�����ܫ�L�J9�׻�^����q��(�{�f=���v�w�<c��.�Bݲ��޵�7�-X��g�ĲH����|(*�h&+�d�ڏ�H_��g/�3�e3��F�H����n���{���.��ƍۉa�)�g�BH��	R��bpj�//��I'����K���zU��W�ы����6G���~;�����{�lݭ|$?b7{'�%Mt��7���
�4�&���џ�^4���dH�L���ތwQn;��p���GbI�h�s�������ryb`ܥ_'�C܃��r-9z����R
�x�q|�G��׸V.A��!:ϗ�gX�I���)e����Ώˏ�ǃ�[���y���'��1r/z��̒C$�!�3�h��{��V�����������Y���䅧�V�M�#30K�++���غ�9�ng��Jᱎ��^AӀK��ρ�ay��-ڡ9���MZ<��"��V�W�Fj/�1�q6��,��9� �9�H�Y���O�8�T_�q���[��i/���*l�掰.�_����=Rf��%':��=�$6:9th������I��Ϟ��>���G�(�#������i]�t�GzD��?;U��
���o�����$ź+�?�Qƃ���7{�a��=�:��KM��g'�:�	�L�L����Qf��-�o�3�G	J#���
�Vy{� tJ����D���?�ѻXJK:
��ۋDKR�(��k�'oO�.�ޯ��1����j��9߷d�y���O����m@F%!�Ҩ>��v��!':}��Mr߈�YhAr��ο�y���o��g�.4 �,؍y.��W�t杢�<��r��h�>��q�Qd$�[�q�,�
��&�M�`����?KI:AN���E|�����t���U���e���@g�+fi�!p0L�0L;i�F^L��^v0��I�ձOD[���=�^��>$�W� J���U�1����h�f6­$q��zʇ2��P
�|����=�f��nz �����8�+CM��y��\%B"�5��쎊��Z�.B����M<�t/�_Ph����O�'}!O���B�^�^a3hn�>:�@�Un �2ܖm"j�?��l�7��@���'�i����5hc�
�(�*�3�lf|��;�f��Y��E������菍�sƕ�]��p�88��Bv&�M.<�� 2=�~QX�zJ{%Q��V���, gr��{��xuI窂Q~�ԧּ�(���n���<B��=~#R���3���L����F�Y[����P��n���T�J@�',De��;U���(�W�~F��h�4J�]
;@P��_{W���!�����;�G�hsʜ�j��W�sU�\D��g(z��U-� -\uj���6@�k,TTo��xN��癥j�Hk����d�A+��3�,��Ȅ�	���w w��[���c+/,�s���,0%����t�v���`��5x/�8=��X=�)c6X���n���Vq�f�J��YM�z�����QH���0Oxw�)��Z�ڂ�ȍ��b	�Mp6qk�)��pA����B#��Y��ߡ�H�'��z/ܳ��gTj��M�6@���\h�b$/7ň���R,E+�{���w���t��j�&gA�����U<6B��N}B�����]0/ܙ)}:�T*0;"�?�?ì�Xy����[�w:�3�-t����f�_	nD>�����Q/�%�^���_�p{T�����%{��I�ۅg\���z��(d6��dM|��#�ٱ�]ͮ��]��	Q��X��y�[�<g���h�z�u�8:]�N�FzOOQ�*Q,4�p�I��=��=���T}�C����a�:�D�bz�h�7ުc��8��T�i�����H��y��*ƃ��x�6<<�*���ELĆ-6bK!s~���1Gݟ�����$��l��)��wr�����_T��N<4=��,9^\�Q4[�vr[<Yv��ٛ�.���ّZ�ۀ����} ��=�I��C�z�K��Vއ(C�L�j�ԣ�R��^�ډh�U�����>��s���!Y��Ȳ^K�a[
h�|f?S5�ј/�V[~�a��p��!s�%ݲ����X=���9���F�,�+�����z��N�t��,��in��=h*�$��۵�"K?2�3�{& ^E;��LH�o���O��#��'�)�&��}���ч�_��/�ޝ:��"�>Q�����"���9����*��!�"��q�ۡ^���8t�%�:�|��t��m�i�P2��g�Z!p��F�8��fӪ�=%@.ٲƒE�v�Q赓�j�z�E��y��U��gG�O�̖�t6�3K���QI�f%Q�O�W�O >[N?j��sړ�hu�)X�M}=����IRj�Y���#������!W9�ǐT�����Ţ$]�����n��I��όL�u�~�"3�$�b�S�I�<�D��ܙ�<��n���{�7(����p��O֍Dg��巊�V���y:_ ������Bܒ&:?X~=�;����+u�ۅ�&7�H�{v4ޣ^GQx;ۮf�W���S���5��GKO����@��mzK؆M��ɷ�ɴ�\+���GQ�D�����z5��p�܎ښvɒ]D�8]��d�U��PcSb����=]�]�.O	?8�_�ynC���(vV�cJu�v�P���q�_���vK�F���
?��r�\�~�1M�߇~y8��O}�G������
2�n�S�uf��S�҃���V���G�����j��X�]���4���O[?d9y^@��+����͆M*r�p���ON��0OO�)#�
��:z�()�H�!z�/�9��OԜ��cίzm<�5,��㫏a�C��<�����3�������ϟ'L�V�+�%�P6��^7���G^{�u��^�{�X�����������6'��\eb6_3�?O�if�x�j�x�v(�x<1�������������c����6���x���l<������x�o��?���xd�?���1ݻzp/����GE����/@�����V棉da".�4|��k5vu���K�u�ۻ�ׇ_��"���$�t]J���Kw����]��п���&�ɮG m����;�����'�TQ)�rs}�b�¹��O��,����n���)<{�y����y��g��MϮ���_�YM�������D�;�����;����&�u���h��n�ٞ�ٍ<�z3��ø����MV�\>ڵ������L~�������:�YE����"��r{�v���| T��W�2���Ddc���HJe4�Hed�Z����6�䪈i��P�������Cty�2�����x����#e`d&���+�����6�*TW�x@�
 �*���Hz�c�ffN���1�/�>�WM�Z�*ϟ�����>U9��4s��L���Y�S1�g��t���o�O�Y U�P��En��u���j�'��$��m���"�C�G#M����E�6me.@��׉�����`��#$3�%�[o'�0q�nKڐP{���Z���VX�z���7�*M�(޳r/�OՒ(�A%�~8F�b0K"� MQm��D@�,~�y8����//�>�F��H���0��QJ�˹�;^t�,��K�)&E�0n^xW��g������v>w��$���˭�FZ�r�����l���[�kR���F����h���������Y��dy��*�P+��:�Ҽ	W/]�ᡧ�,��Q���&�T�e��y9���J��p����׍dh"���?�{�|�^�l'f�v�v ��;"j����(�UO�� ��
u�?�B���C>dDD�a�7�`K\G�w����m�La��h,&<�덒��k��P*�iv�-̫�q�F���p4�;A������$�x��JZ�P��rP���?�'���h(=�U�:��VK��
-bq�r"]�:�yD�i��{��d��»�Ga�^(O���
�XQ�[�(�b$����PW�tuA�qR����?��hP��U��T�ci]7��T���6������`\���0e��	��g�����	�)P����\NG���qU������ߢ=�|	RM?�:�#?����<�Р�D:x_�v�BV���fF����<�������}��x�����qVQ�=�Wn�(�ȧE�ŉM���S%����hŅ< �}̘+9_-��߼��X%�`�D��B��-�� Bن��C�Q��R%�d7���+>��8�p�S���:$~�΃�9��mB92�v��/�K9��إx�#%������ᤍ�S�܏8y�o�HB������\8[�2��w�ռ�ݍ|��y9h������=)o�y%��3ygpU�͂�`�+(-~����-���A�7/м�UU���I��Sp~���[;�zf�eט���˟�y��z���Q>�Kp�o:^{l>��9~���R|�ü�v����官���u�sw�1�s�3Xf!	��ꎅ�(���UP�0f�q�v� ��VQd��jvP�:3��`�Gq9H�+D��Ӌq��p�~+7�H	��R`w){�J��ӂKN���o�y3.�,a�S��}�;�9�D���v�d���~�cy�:L�N�.Kt�̅�~�e?����Pg�4��B��NX�3��@��G�����,nLl�~�4��r�����Hױ�@s�$C���M��z#â%�{E����S�ZL��O�S�6u�jHs��k5rIB�	���(_	�NԊ�e�l���ڕwqyU��XHTVZy�+Ӈ��(��Wz�Hmc�J�F~����'P�LiU��g��m8�!-ڎ��Q��H=e�b\�-����s�7N9B�*���� ��rw{�m�'B��ƥZv����PYB�Z壀�4�S���9J�B���q�ի�W�Q�R`E��5��&���ſ|���B��j�,$�3P��5;��wY���f��6Y0V�&�� ��taU���|����uhJW�
�M��psm+m|K�y؎��}xa�l��@ܣV��'��h��dG��
HA�sA���[���E��
�C�a`QZ���0�/`��e��u:�>�+]jm%T�K���1�R��BN9
3�H�h�aS�t�2 ��kV> )�9gt �b�G	9-c.W�BN��^����� ߽"�v��ʦ0l�JrF����A��3%(3�B���L���X{��)��(�-��3N��_��$݋/�Q�A�=�?� ���w1[��o�rU���x;��ơUe��s�J����i�~������S����n�G4�ߥ%�X�5��Xe��F���ʾ:h"�8�7�E@n��<���D@��~�@.t0I�g ��,(A�9:���Fs��C������=�gg@�!%4N)��X@3����%��!� ɥ I�>L� �i��q������4��8�t��VWv�v��IJ�)�& ��j:ɩPGz�*qM�!����{	�9��ث��a��-��&X��6���pX8�E��M�wG�@s�������K�x%����!�?��1��܁2/��L�o�yZ������-*�+"_���k��mW��	r��d�Tu-��2d�?c�,��HT�g	yj1��,P���E�����,�X�f��2X�N`��j*�˯���8ݪ������e&�h*㸩�0٘iea�к�����,�0F�+�0�/�02$էY���,܎�rF�?u���,�jj#>�zXu�<&a�XEv�Fq^ulY����Wz���(�v=DaDqկ�a��E�����#>��-��;��3�wȍ�ߩ�l;�<�R^d)H	���HM�fpSG��Tȸ�e��M��{X���)E,eKH�|#K�d)9�"��Q,%R���8�"BJK9��������}eGG0NScί?��{c$�*v���r]/�oV`D|i�g:WZy��+�)*�Y��z�V��0{�c�/�'t�TͮwW5H�'���6�!���T}��K|�D�!8�F��p"Z}^o�����k/�.�(]Wc�fM�^�db!����C�x����$Cf��U��Ê�A��Z��w�
S.$ؽ:0��΀`*S�S�si(���-��7>"�.?&,��
�j2sGi�)ICE�E��a¾>��`��l�z'�:�Mtf�V�t#�٬��7Q��&���&���	{h(�L�1]A-I��}���X�}���c�z܀�/޽�(AQIn>�h��rߝ��G�y�a1�j��	�y�����_��nUH\H��f��R$�N:r0�p=��;H� �n/���vR|h ��[��c�@E�hŽv�y$�s~��_���G�!#��4��t�̈́��L�qw��9�yS?!�; y !��ՂR����t�[�{W��S���>R�"R�"vC�6R�hQDL��"�[dr�p��f�2�CJV�\4�'O��O*)��|u[�	��s�ЌEO0-���T���@+�I��v&��F��tw����[��7G8��� �
&'O*��5�<�v�x�ԓv��N`)@�n4��^P2E �&r���?k����I���^���'}��R���'��b؉@`�������ԘU{Xc��~���-����Ԇ6�~
$V�qbj"�������# ���L��j�����M�KH x��n�F���n#�>�p�� n�驺�'��Ns��R8%S�YJ����1��EK�xl��n��T"�I��V�D��3%$�c,Cb��G0�UR��,�:+RL[M��L���_*����<jz��Qص��-���.W3��L%�^�����f��6�"��r�<�rr�0���lE��Q:ryv�ɛ��>�_�ױ�(@O��E;��hi��3����D��ا�U�䘭x�@Tv�CO��(�S9J���DC��F�G]� ��p��$S�!��L���/��Sw���}� [Ol֮'a�i��J;��c
��?���=W��6�=��T+S+��,�0�%�F���i�$����Q���������+���.���I��ݩ&-U��c$�SM��n�3g4�&f�ވ�#tM5�(�?/�8�)̩/�om$դ"�ݪ����Znp��Z��0���8��o�;�;�V/�+��c�x��u �j>�]�S���4A9bH��~M�G����zG���hIz��!Dn;�Q�~JqD��=[�7d�����d��F�������-K_��+K�rT�ò��3�rò��Z3Z�>����jLa���H��VyG4!4}`a�GN��ox����h#����3k��T�icߥ��%�җ"�,����Q�=أy�"&;���OQl޷#gGM3OJ͛�p
5	�p�A6<P�5�1�f ���B�-�+��y}�A��v�+����\�,��6sz1�r�D�ӿ�D\p嘠t���v��7���oN�S��#��y�W���*)�w<zk�h��0^{��b�z�s�T�+�t���u����!:[�ǟbtt|�ױt0^ǒzy��n��n�e��S]�4kϸ�]��`$��#{nB����3�еH�����i6!'�$K�8�)�[��� �K^P���������\�@�<��G+pvJN��T��_,>�p���6d�'^ ��̚G6�-���#_�]e�^�[4�q�^��y�+�Hw�Xr�	�݉�
�5K�V��MX�����̞�(+ۉ2`�� +p��Ș��ő���1��j�d!O%�d#/{�X� ~"Zj�O����_�)�G���%�p�di)�F���<�5f�<<6l�		�(%�P���$!"%��)��D�K�^|p�)��=
�V�����n�Ͱ��D�Y����<_-Γ7���בWl�.PC���.v�6��N&Jw!���Izʒ��b����2��Ǣl�^�Z�� k��XQ�C�oF�Q1$	��Ew0ЈS���&f�,��3	UC�w��f���Ѣ��#��3��W�@ľ&�؇q�GOD!���(�����}04�槬�wC�gAO�Q�O���z�Q�{[F�|c'�����	4�6�'.�i�h*��`
���G��e0�āV�-�ufj`�=�2#ob�f*B�B��ܫ�7��k�z��^)���3�G�Eí�愐w�N��a+%͡#&C�$|,_�|K�{��Q�x�ze;��ϫ�k:�BT�4��0�x2m������:��.�l,[%1�d	��Zz��V�{���|6tei10������F%SŦp�+u�sr=+ %s�צ#�	���p�E�]3Ø/�˰�0�����h8�"Ӕ���=��>iK�!����Ʉ�<����X�y��X+Do��(ٯX�E���S��>���m=%�e��b��(�U�W_&*���mv��NC��J��e���#Mp�u��WL����3��츾�����荺Kv(�j�B������.����)�LX�������Pj�G���=փ��vB��� ���%��+O�© 9G ,��1ʬ4�_t(�ƲP�2+��Ҕ�T�f�;Je�������81�q�8�����;g�!(}��p�v��u�։�p(غI���:���%P&>��~�'Y~c���P�k�,��3b��~K��u���s� �{�<M�����ʙMt��	�Y��8���M��#����~�V�<��f�HDZ�̲X��?A��uU"����z�\{�����￈��w���<�ﲮ�D�U�����s���kࡌ	���?�?���	�p���$Q�7��ȟ�od�F17��H����k�Y�X?�� Cy;]���xG��١Y��&љ[�@��AFU�4������� ��J#� �E@�D-+%���J�S}_pHݪ_�����ie�'  50��[��i����b��E��`�ΧB	^,���8�yh���Ϸ�����|�,b��򧸡x��Ê06@M��LA��q@u*V��fEWG�}��٩��"���\�P�����F�����ï~a����U��$�̽R�8�?�j-<�O5�CW,�3��׷Њ�J��
$oF����؜��@�@c�bX�׀�G������ڌp+]h%���I���TE�zĞW6�\@��BLԾ&_OI=��/D��,6�#`�8G8�8g}F��<���\+��W������^CTQ��������tyt��~��ş�_�/^�/^�7^����������������y��9��Y����i���⎾����{{o��d�/�i�c�wroO�;g"y���|���{��F�}�G)@�O�a�W.M��"wM��,�8�-c��_[u�F��m٭�X�R?K��e�bJa��$)�(���"�zKӊ1���2��z3fi��H��ш�i���±�@QQ�S�h�������6g�΅�ܣ���L�+��Ys�΅E��E�W	O����\�������w U��	�/ƒ`�@�-�~��f{B|�=����M!�R�!D�|c6t�+���oP��x�%���e�?�D�+L��F+e��d��hfmc�a,��7H�"���Gެ�޾@׹-���SH=-�8� �>Q�=F6KN�#�n�׊V �[[3\T��m8s��:
�X��״�As��ڭ/�`�����/Ԍ�s6��;�*���9GM�0�Mº!��0j����/����PS��L��'���%uE��טs,^4
_�B��Ƽ��Gd�M,宰u�n2-��*�Lg��BTH�� /R[���:�R3���ц1�u�(� �f�0�"&��ߐ#��C�{���}RN �������f�K�v���C�@1��n�yo�Z��u>�pd�г�����z�!��+��4��:J�󋲫��H���H���:�V^i�ss�x�9��T]4d�C	�������ą�k�U��n�tZ��tV��6���K����r���K�+xyfѲG�w.�K���k��,n5�gW���7W�0����jLϭ��l��f2qOEˇ�吘y�-��;�m�ݜ��,F7��҈޾���s'�m�c\���p���ɒn��T��8���i�y2/w�[>�v|�6��T�glJ}Poi5͋Y��E�R �}����!&���ddL3����FT�fy9@~͌��.,����)ȮC9�B�]c	P�+`y>bx� ��<b������_G�ˀT`�x�$��HS�+�{�e�ZM&uu�$��~x�'�������6��C���C�J���d��0g��Cfkv]U�[�7B�z3��ގ�05��ʿ�E]�H����8�v%ʖ�����Mo��&R���<B��6	��W]��,,Ë��]��F�ȫm����Ձ=F�?��G	���UG'm� �B�ͭ�;x�7<������NS�\��nA��}7�͙�gM`�=bA{������p�a�H�~�.�J��KZP��S׺�[�aY�.�F�QիĉAo�@�;�G���5FPv����s���k%o�M�x�����7/U�zH�X3��;QoV�����M��q���6z{ő�����9@ωQ�a_�$G�a�ղj�P��B��'jM�_���e���qαr�uU�l\� ���w��o�[�m�*N���,�.;��y/��!pr�E�� v����ʯz,Ȑj�!f*�!��������`�%
���C�UM�c����"4�ylu6~����X��8���R�+�!K���������sU+|Aߍ�cW��\�AA���Еb��"�T�U�\��J���5���\o\E��j����k��<[q�  �w����N�����AW��,W�H z=|��u���e�*���`��#�lܙ{W&4�`�D3�Z"�&c�U+�U9^��/�k�v�;������!1x&hRXs׉�V>`.޿?�#s�b��vvycE����)bm�����H8�2�샲�����_0�<S$����c~P�#\���)��O�9��V�?���$�_H!��f%6�ӌsL�q[�rD��+�Z�l3��9j�3#_�����շ�
R� P�
2����V7Raؔ�;��*�����	�
�V7I�{Ge������b�N���&�9�I@��޼<@b�iM�/i 	3��x��������]"�[EKW���?Û�@�Yu��A8�)�;nC�ѭ�̫:��$k��gv7��4(;U��N:��E�G%;�������M�I�G�W&M�g��N&`�(X\u��_�����3���x��O$UL<���e�E�Լ����J����Mç��ζ��SO��^��
�&zI��^���{�M�S���A��t�eDN�4���yv�����G�q_�N5��o6�
v�s��;�Q����}�x��S���-������������d܃t��R�����c����B�ޢ�~�Y.�A�����&m5�����v�Š�u���l\u�o���:��2��H-l4p��h�ջ ��4F�F�3C^�>
5�q�j�������Eҏ���g)�����;U�g���-�ÓG������r.F?#�{��ގ���p >f[�l�(���c���U�v	�iu�Q��vn��9C������`�.l���e�>Y&+�)F��}#:�@�X(����6L�y������=xPiS��7!�����D�5���k���\n�]�&f-��hWu4��G:b��gWtm� ���8�K�:Y�"��M�]���t^/�w�`"�w��/���:L4�@��0��2T�sp��7 L�j�t ��UU��	7�N����eI��6��N��!o����LR<�mIp������Ё=@��cͧM&���uu9�Y�Lp�T��J�{LΩ�X^��( ��j���3�<sęa�?}e����r܆�b�v+ݣ����Rab�VDqJy���ʣ�L��Q�M�fD?yn��^�l�kM�!�`��&���C�:�M����'����x�Z��)���G�G�j
���M��y?o]~)����\�e��/�5`���f6��s�X���+��[��Z�E���v�Yֻj����gH+�N/c�r+'ԓ���Np�7��A57������@�P�^P��g��;S��0��vn��~�P����:b� ��s���A��]�D{��;�ŵ��	ه���p�"E��
��Gx���V~����N�c*�կ�H:��lw (���u��,�Ѧ���4���$�]���LCͪ�$�8�F�nk6����B�3:����df��.(GQ� (�����8WZ���<����%��̶|��V���|�ɒ�
��%��;[�hʨ��5V|N���%F�-���������z>�eS>�l)(i�W��i>$9�-˭�+,��ٔ���Ms�����Σ�E��t�U�� 8��g��b�b;О?Ax+�G��P^>cY��O�1��m���1�[��j���()�6�<�g�����k���h����g�'B,��D��7˥| �N��;��hW�G�]��Q��]?cSZ�.��Q!���<�����S�������L�#��<��qx���u�=n�t8n"&�^z؈��RnWb�0��տ`-�Q>f�;W�尬�����6��4��A�}��_���E���/L�O���=?�o���|�D膲3?0��l]n��V�({h��?��t�N)�1ߨ�Ɯ����5-2�3��t7�pݶbr8����`z�`~pX|A�>M,��j�'3�3<C03�#޿09ʧ��P�Զg��Ě圱���7���ĭ���zZ�ܦ��i�l4�Ul�h�Nh6�,�+�v���|e/���`\ۧ���.ُ �-.�:��-��B��~�j�;��QA�Ϯ:�$s�J�X�Q>,�Я��Dl�&��Ƴ�&X����P��	����G��Z�F�i��G��t��k��{����nj���a�VȜq��0u5{yX�̒Ș�IxD
�u��/�D����&��.����.w�y-�?��bG�J����Eg�So��g� @��΀��dg@ɛ��>|o���
π�_�_p|�Z����g����g�������3`����������Q>r��H�����k��)�Ma
H�z�?�g�]�� 	�0D�(g
�+������wW	��n%�;E����Q�Ūt9�ք�Z���D9�f��(D_c��&%M����$��d����T���r��{rR9Q$�C�� �3�0�2[��~
|Ny��*����v�Y�T-j�3OB�g��S���3�k����\ű,���W+��,�	�k�Gg2�+*�L�.�83�{b|��k���3%�<�qO���Ԅ~���3�12��Z^���"�K��5�5��[��Mk]��[���^}LspU�@d��<���N��߈���\��B�{��oI�c�-�)�'���.�	����кj �
-���b�/?h��`,8�x
L�|#)�%m}n�X��Öp�嬰4�l�o%��t �:��D��>������Zp����cY4�g�Ǐ�+6,g{�e;/�b9������C����J^�������H��u�~��7{U�,�Ȱ���q�ZBK�����ZldaH�+�M�8c���E�����$��;����hn����3��P~w|����͐�PH�N�MC�iJ�v?<���بf6q��Yخqi]����m�,[+��0��$������X��\H�8��=�8*�E^~*c1f�'85η؊�+�����q\�����`5�d�ۚ��j9�<�=v���xT���-:$c4g�t
��bX�࠺��)X�~ժ�Ώ-�h����t4��Y޸̿��U�	�ɭ���:��er�{��F~�7��JtZ�*_�����1&C59^��Q9��i#���f��h�����=%��K�s��E��Br���<10�R!����J99�f��D��L��*������0+Ai@Gk?��R~"z .,�U!<��5�!`�C���w9�i43�;�srn�M�"��Y�=�3�o��������C�����ץ.K���x������u��؛���qhe��M�&G�Ͻ��掖^%�P��b���[����̀����WyJZV��+�nHIŞ���{xnC����	�a�{�E���.�;UD�B�����<,YJ�SQ�*��㖿�2?�t�es՚�B���A�|	�[����"�����1����Jg�jY�<���+�\���c�]��LC㡹c�o���}X �a>��F� ��Y�Y^�����6nC+|�>�'����Qu=�/������i�#��6~�1!q;�x���T��><"�x]�l��C����&t�RH=�l���}��D�湩��W�u����6U�Mޅ��&�<lu��I��wn��Ÿ�n��-P|�Ӑ�o�	Նѝ7|�v-B��FS�X�&�[l��
g[ �Rp�D��RWb#v�k(�O�/EM���=ڨR���1u�m�
}��J`i�߽���6�\��b��=Jyz)l�W��xV�I�զ*;K���%ⅆASɦq���V�B�X
h��Rޟ�	~�_������o������AE5So���T(��H@j���dr���hV�*�,++{(�륽��M�V��v����v1�˽uo���]{�3/����~���ut�w?�^{��~��9{W��q4������鳥��hMx܅\��v����,`���R��m�]�gc]vX�3��m�0���� ~������~�����H?�O��i�&�t��nNϜx�l�Oи��F�����!im~t��ܫ�0�DhMFH�R<!3�`̚/��x4f�1��7b�{_�KB[�4�\F�ƚ�^ǇERo�)f�.���k�bI����X����;#r��zv"��g8���vv��E�\O��(�T
JE�҉4^�_�];�^Z���y���1��)�3qMF�d�������ِ����̺��ω���+�m�{����Q�=������&�Ҍrɴ4��2�6.+{����壖��Fz��EFΝ��Ɛ>_��b7�{��5��~���o�%���#M!}!غ��}�d����h�������jO�nh����Z�L#m_�j~���/�מSK��Ť�a��,zf�|3G&f�z�<V�$�&�գn�ƘI=t�a7u��g���>����'����,��gr��ܸ���t�\F���zTL*�bV5�������CK")Y��{�>>�TaPy�f	
���Xl ��u��k�A�0�ğ��q��	�/so5�}C���P��xm�yƺo�0�`��9gm��Ǒ9�_� ��e�{�.�Gq3�{��̺#��|�'o���2���1_g�ڇ���c�?��C/!�E�2���M!�Я���Nʩ劵�� �x��|��.��s1^����l�Tw��ڰi��!1����L�\N=���}vm�,-�C�6��j\��э�{B0�V�l9�Ϳa&�:�'�=�c����\�� �lH{���%Cɋy���Q,�#m�h��I>k�-%�^9���3N�D%�)��Q���.����MWh�Eז�+y�/�x��H3�ם�<Ɇ���u�Pm��F���T�$�H^��˨%T�J�΁�fZ q!�^Uf�:�w�^v�@ٷ�̂������CG�����|��!)'"�rɒ1�Q�o�勬������YRhfݏ4�<s#?��w'�:/�:�QX������;l�+m̪������U7z{�ʐ�u�/�P�Z��],�	�?{�qҦQ�m�'�\��vߋ�->Ͱԉ�e���u�[���F��������L_c�Z�M��V����޹��L;��eT�d��������k�����1'п��.C��i_���U��rjh_{1���x;�at-��{;�1��`{|���q},�t�����&���֊N��`E��Arfڏ�����`E�������e���}"z�����z�����������;���Nf��dbPGU9�a��!�Vl�'rx��4��#�c�7y����t�uD��(�E�e�������m��o����:*i'=[�c�s��o鮺hT�΁d��TiQ[�ֶ���Ym�=�CO��<��$�ۋ�85s��hacTV̡����������{.����4�wcvF�5��P�����vhH4c�#X�CDԛ`�����kmJ�ګ�i_�Խs}5���ml�ϥuJVmx�Aѵ3tT4Y��âd�� ��`���¸vT,��i�P7iq�fX��L<lH;@�8��B��5��Ys�,�5�m����3V���7�����e���S{Ѓ�4F5ս����ds�j�GTm��5�XcuUX��&$7�*yM$W��x�X���N9w��D��z�$O��!I�I{����F:t塙l���#���C�c^�k�)���0ګ�o��k�X=Ӧ����E�G'���~����{'Ic��'}K���T���6�+��UzfXUF?:�P���<�;/��5�cV�>�b7�E^�eR�Q�`��e��G�F�e�a��{Ӹ6�2T���������Zݫ���(���uXZD5C���jkÌ��a�+GAC�P:އ�H3���	����IFؚWܽ�y~m�Ȃ������ӄ`$�0��B�ok/
�U���:���W���d�:j�&�����7�#&��B]��Ô���0�#�>������Vmh&$���`{���\١_�z�T̚�?�:��*󌇲PϺ�u{�|K�JО�c��w����.CWz����D�ߌy�T�<��кft��=��d�������,��ȳ�~���&�1��z����H�.��?P��|+"��mE�w��o��؜ڸQ���.���.�3�97f�5�n��XzДv�5�c2k�]{k��ˡ�i˩CZ��Ϊ}�����¤����'�͟�ņ5�S�{{I^J���9uo��Zs]b3��g���{Wk��x~�����f���阡���%S�{���� )�x�&v �.7�5-- <I�緎LkW�U/�ꀹ#���֏W�K��js���J��U�R��>���"xEok�U��R�XaI$���?������'�g��za{Y����W����T_YAWn�Y���ڕFɜ�ފT:����%�)Y@E��t���H�魇'�VT"����,�Sx�-Umn~���a�;�{&HW�L�Ŕtwߩ�#�v��睈��^�'��������@y�x��}c�/��UGmnR��\.���V��H'�Ol�'�5�OG�`�ԟ6k����yIA��U=��Ϳ����VO��W��oj���_]_��H����&M�2�����o�o)/�[1�E@�b�9����u���z��d��86p��K�<܍�5�/�W\=u�W^g�љ<�o�6P8>$�9��J���/$~/Q���8��%�#q�ę�KtH\'q���$�(��O$~%�{����|%&I4J�+�-�V����xTb��6��5����%�H̑h�蔸R������$�O�I��D�A�z��%H�J\)�^�;$�,�}�����>�%�-1Ub��ym���(q�ė%�#�s�?JԽ!p�ĳ%�K̗x���}��Ƙ�E���`����i"|k�0�����G
	�N*�#
K�Wa�,����8�KCfa��3������F��y��Y��`c�O�
bC��U0��J��Z��;��ï"���Q����@;~�)��E<��K21�YyIL<;rҳ���,�+���KW�Ө�0�m������?i��� ���+d��r��R���;���T�O%�I��E9m����N��H�d���e��p��WǎujF�R�V���;(�n.�/�U�
���Ӯ^s�6����Ү�6�TFj�� ҍ�]����}9�iA���Ȉ �\����4B`�ժ.2Y�%Kݪޥ^�Qm��!���TK�v�R���֫���[��b��`K�êV�6�j�����V{�b��Ti�XM%VUڃŪ�L��m'�"�_���g��7�&3�DB����x��-R���T-���d��U��N]�Mw��6���,EHPa�-�[-��.�c2��۬K�e(�޵��V+���J��bF��Ų�.�	屪en=�iV+-��߿�6���;��=~���ns;�V�ݡ:M���r ���vu�G}ڕ�yH�Z���Y�Yk*�; ���)-׊Ͳ+�����A��^���ܮ`������K|��nB�f��������rY�flo;Q9T�ݳ�\�O+�W>��;MN��c����r�լGqK��Tϟ��Yu�:-�hn�Y������
��g���PU�;�����;jE�vx���7�_`6����8`��2��KMVk�\Yl�����5�fi��;�����t��`vgf�ŝ/Ţϻ0B����b�0�S.T5�9�پ��-lᗸT笒+�}�Mh
s�|��\n*T����7\�	q,�M����*��V����Md�(��\wzln�7����h1ű��Y��"�f�]��e�Y���<�i7�%ML��4���gVK��Y�Ʌ^cV�&��ɤ���ΰw����k�ZJ`lKѧJ�Nj��q��V��RyO5��y
?�g��t)bTSY����T!ë�qZ�|�#���bx ;�0;��eN{����+J`�f��b[���H���b��-��˸��"��H*u��"����u�>�/�a��[-�UH��8�pi/�6J�AST����
lҬO_ju��3f^N��P6���!�%��F�5�-�;�;��m��\]�M� ���kB���uWE�	}��Qh;�q=ׇ>I�I�s�7�,r*�c*�C�1�U�CH"����=��|���4��m�"ݹ���*-N��r����/�S��6����P@�*z�O�Xo>�P{ۭ�����/��V9�`9����J|��U�-�r'�\��OC���G&2��&����x�M!x0pҊ�E���Ώʹid���l!�n�y\��%��p(@}�&uZՆ���h��!��N�����=���V�A�M�a�������u�>�R괻�X�̶��f���K��/��ƍcS0q-r��|q��?��Z�Lj�����m�^�++M��Ě?��Z}�N����e��,<$6,33�]�&a-K	���s{���IIs�{�U�w���b��Q�K֛�t ���I���4��>N�?��G�-�:?�MA��������o���WBB�z���EDF���ۯ������':���G�1r��?��x��c�;n|҄�)�w~��iS�^0-�0=Ø9�¬�����ʿ�����s�^:��._Xl*)5�e��-W,�V��+�.��rI��eW-���k;���|�y]�\R�Y01y�1'G�_u�u�+�р��U_��:�W/���5k��������F♩�s��>h��|�k�>��������\��]�p,q8ڵ���K��_��_�����г������+��)=��~�߿���������p�o���iP|�zzX�����>�����?���?�\��,���i}}�Qk�^�r��5�]_S{Cݍko�y�-�޶��;��p����{��l|��a���-[�롇y��m��ɧ�����g�{~�/�nڳ��}�_��W^}���oj~��o���w���{���G-�鱿|���㟟��˯����|��?�������ǟ~>��'��'�MX�������߾`�<�?B�YY�+*&{�03�s�����X�����7��O~.c�\�oTKq��z����+��pGK�B���"�E����+�7�0���B�VrM��r�~�Z�����q�L��{�/�E�I6�$y$闒,�C�)+4�=N��˙�HcE����cl�j��~E�˵�x`�G��Mr(=�!>�x�/B	�R
^~	%CQN�F�QT5���ʘ�7뒢Q�-w�E�wӄ�-��,�w��oY j�:&)���0��<Cav�&�ȱ���hJ}�[��p���0~�������]������R�J��Ti�/�XT���P�L�C��:�K<�ٵ�5�ҕ����U��/P����_1�a.�rn�]JL8�1G���)�r(1
�Aℳ������`�(�m��ҧ9�I��]�����q���~	�,�d�#
�yX���P'P����x^B�)?%<��'��GԱ��H6���,�פ���0c�G� ���և����N3ǲӊb�i)}�i�&�nؤ�	a}�~L�e�.����H���`	fK(��R�YB���~�a,���p�E�z�i���"����;{\�Ӏ06 �7��Ms�3�mxƗ�Q��=�K���X���ơ�qO�:�Q���A��P.��h�׬�ܲ��/A�J6�#_`�{�1ah��,&9ʡ�i>��@��<C�ؐ�A���qIO������X���O�b�q���b������}�}�J��[yvCy����d��1l�5��6�%P�}nw��.��G������6�9��_KLst��'����jy�d���A�?�ٿ%��oSGT��i$t��]�Px{�XdA�C�)L7�ɮ�F	�vբ��0���a��z簶!-�̓��Jl8�u�f��_lr�&%"�E$�J}�}bC�}b{�ז��Sl-r�!����8��%�:�L3d��P�B�>���%0�;e��bz�?Kh�2��ׯ��/���M�#Q�#��#�#:vZ��#��G�#E���#v{,�="<�	>M��	�z���X��'Ye;�r�2:p�,�Qoo?�2������N�A�X�:}����|����|�F	��	���Y��&~밤�d��z��/륰+Awk6���b`71O�~|l�{�����~M�ڇy�{/RaC���&o�6�Q���	�۔+COS�B;j;�Pi!���F���lhJ4Z0�m`ˀ�~M1^]%Tإ�CZ����~)}X�����k���^򑭢\��WlA�xy�`��}������dQ�z��BvJ�G�),l�߸>Da�A���_��C�^�ŗ��7"l�p�@1���ɗ0B������/�w��M:L�3���o���[�����7����#��O~�=;�	c�3Ow�A��^�ـ��OD��ZÚBd����I?���F�	��tǲ�1�EYODi���D6뚴vM���m���W��792I�O�k�sa����<a t�W䑯�Ϥ��2?��1���%�7��ϼ��|����jv�����5���6�\�(��"�W`�h^�Q&:5+�̨̄�8̮�mQ-ͽ�z9C�4�:��N}%z����L��r>���*��"c���N?*�μ���Ӄ>���d�P��
��{�(�{��^�ۅ�����w���0���ǡ��x=�f�}áE�͠�;(/c�_�,C���1:6q#�D���^хb�
k)�z��Hք;�c����pư~a(K@���>����S"�h�j-�N���T��nG�;c43c�0�ND�ơ��Q>^��)���ѯ����-�D�!�{d��!�?$yPS�PZw�Uh�E6Q�����e�f�A
�=�t�ԡD��h���D���;��Ա�\������~�	�X|�0T3(~���*P�I>��B��d/��Z%.L�Hrl�q,fl�b�\r��$7 \�N�wkO�>?�_m�.e�]7��X�=+y��?L�;�E:���4��乁��aZ{o5�Q������6�rYc��y��|cP�o��t��IO�!���Amq-��c��E��8�S��:`F���7�5vLS��OqT�2�֮ ��0�X�o�J�m�س�;�9E��c��aT��0�o��o�Ԋ.��
���!I|��<�aO�_3[o��۠C����#�p� 6�ܟO�ǆ?!V��4�
ǈ��+}��u���C<a��Yw�n_��h6�V�������F�A��~�jofl nP8����|��� /��D"l��"=��E�vk{]�Y���6���;]������pp���dƉ:�®t1��:��`]츁���O��j�]����7�/K6�f���;�P=Պ�vU�j;T#�J؝^�]��]/�J؝^���_'�J\�O���:QV®�j�kDY	�e1�_#�2�����V������U��^%�"n�t�e�m���}^�V��ɢ,�����X/�z%�N�G���B�08�R�����]��o�2vz��+a��j�?x��a������
]̾�}�����ݍcS�f웫�8F؝.,G�\.�1������t��aW����W	]�*^�]&�!�`]$!��eB�.k����Q�R�����V��}U�.����%�=�D�ap�/U�l�B�]�b⯭� ���a,�R�kxe{]lD�f��apz3�*<"}��}�۰&mt����/D��H�����N�b]Bױ���D�~��O�nF�2�0��/N߳�����s;���J�~�R��o3���~+�ߋj<�1�j�	
ǈ�:j���A�qM���c��36��~<�^Ba+����J_6��@[?}[�p� ;�:d���m���	r�M�^�m c�
لJ�Pֻ�V1Z�8���>{�������q�kHK�k,cg���|�j����[�a,�� ��wz@8�WS��R���w�X��+c�[P�Ά}3���~qJ�ެ��|�E�I��;@�}H?*���c�y ������PĢ[��q���ү�ch>�����caH��б�@֧�?ep�*�Aΐ$��(����m�,/���yx֖�����y�}H�J�2�Y<��zcEBQ4��}X­��ЋE~�I��ot�Z8��y�����$�=Z��G��⪴{{���KƢ�T>j3g�:=)a={Գ�[lK��>M���b�|�����yN?O�Оe4kϓ�3���]+�;�u>���w_��K��w_Y���|�̀�J��g����B�߆��[�3����Bs�]��K�j�}�Ŭf���,5��ꂐ�&�Ge��W���#��j��2v>�����f�7z�o��|�
k/g~��Mf�ˤ������e���*��!�����E�y�9�Ǚ��uas���!^���!��G�R���(u��,�1�43�%�Eӝ�i1�m��(E���r|0$K59x�}�-��qgx�N��.���f��.�?�88�����Xlh�	aE���o�N��V�Kiά*U�#
�?�'�!�N�_�v�Z-R��P}Dsgh��*��m�ņ�����}�ǡ}ܔis�_�k)&��p{��H�Z�f��
���`b�6z�?���En;�M ?�4���F. W�Tr�v2�������
�R�����T����򕿝�}6�6�F����:��f�Y�h���gT]n�})�E��1��}����A�ʬb_PO&�a��7I����Pek`����nW����g�އ.tӷ.k���G��NR�aׄi]����lo�r���Ћ=�si��䊱��⣕ʨ�E��Ų>��@�,^K�eV�zq�~����꬐܆̱�Vf.�߂Φ/�2�80�M�
Ta�E�པ����9�f�a1W9�9�SV�:]��_ۣ����~��y��\��D���ȅ�p� ��~hj�hO��8�������!��5
�Cޘ��F��ZG`��Dv�_g�ﭨތ��߈��	�%Q��2�v��E�k�����#��j�Jڀ9`}���VX�d��uX�:�֤�bݙ��l�Ϛ�Om����p���m&�ف{�6�/����-ϯE�՘���iJRL�#/ƽ�ZxMp�/A�׀��w�5�W�¦��u������e�y����@8��30�7�q��p���{Mz9��-��B^���'y-(S5ʽ�[�W
��=,h#��Bg!w5���E��i������e@݊Q�b���ͨCաV`(y7�>m�Oҥ�K��O���n�ui��:�a;�Ӷ���D�����^�<�	y���c�d�z*�0ĭ�Փ��~��!<�v� :
9��sA@���}�|KacAE��@���}��'ār@Nн�W@���VX����7P�;
K]
r�6��@�AVX(t%�&��O@Q�*�lP>h%�Q�k�6Ј�vh�г��A?��x_a��@w�^�����RA���@@�A}��Pag�.����@/��

���@kAσZAZ6d�z����c����@����z}�z��@.�&���Aџ*l
�Z�z�3h�1�@Nн��f�I�9QX6���t��3��3��,���^,�� a,�E�>,��e1������,�d��`��6�c����t����l$�F�?�3Y";���ưs�X6��gIlKfY
;����g�l����6�]���tf`�1nY&��.dY,��d�����,��.ưSȊ�%l6���K�<v�����B�S�W���;�2���3��-fVV��w�+����a��0b.�`��]ͮa�-7Z���^8�F��i�4-�;-�)�;��r��Ud�Ж@���*�"Czz�/�^=H��d���S���胸BLJމ��\4�n1k��0�Q2���I�Ej͎�RwG|f���!߅V{��Z��u�2��.�ʠ�¥%vk�M�a蒍rr�b��p�L�//i-�c��$���g��P�Ѣ^�
�dw�0Ʈ��o��ڃ��w�+���t��f��:Kמ��Z�'|b��L�n���-�����P��j��X{TL��;��A_/�DD��Gl3g�vӽ����dSXnw��<'��V�.~��뜍ne���N@)=��*�'$��	f���4�N���Ï��fnG�DwW� �_�m�X�7�]�vW>����#NLs]�uW2KOs��c���������{����ulwe�g�y��qZ}���Dw1�U���Nc�<Vk������E�N�Ԋ�����pt��R����cЮ&W��E����D����%r�Ð)f�Nغ\n!��%�S-�a�㵟S|x��E��ޓ������@��p.��=��%sOfn�ڣ�W��l
vu3�z6����]=��]]M��L��<ݍ%��N����`W����\� ��v:�z2�c�y�=��d
vu?�~������j
v�`
��q�=b�t
v�d
n���<��t;�j�#ŒRW1޿�"�Y��&7����rMUb�59��ݹH<��,��i�˲L�U�qc�cr��fK��#�	���%b0j�X��p��'$U�\Z`ZB7����V���-��%v���~�����+��")T"��Cg+�<�1;-JGJҩ���Nb��H�7H�%��rceX?PI>B��+��ϐ�|��@�J�#�_*��pڋQ���8Ø��5Bփ��e�WH\)�W���R�~N�#�/���l��m�����!�ߖ��.4�u��'�:��p����I)��˝z���;E�9�\��ػ�0���Უ�N��%�%�$�� ��M7J���8Wb��x�Lb�R��wJ�*q���U�%�KL�/��@�-�_�N�%��X-�!qn��� �^�u[o�,q���P5;u����Ɖ!��v�e�^dSJ�\��!����������*��~�?FpW�����8!���!�'�~m�b���%J?��>��/���?@�7J���K���K���I�PM޽�?L��J�p鯑�ӥ_/�z�o�G�GH������K���J��/J��/��x��Q�c��;�J?�(���S��v�W_���|m��b;�D�������֫�ͦD|�!��������@����I$}'�)%$�O�0��\�R7?��f�+h�C`�5���Oû�N��Y`�ħ{�o������a�o���s��<�]���w/W��{Ż������a�w�M�F�L�,���\g���5�?w|>�J�ºօ>,���I�~m���/y�"��e�ZZͯ٥��������i���_����e�,��B͞�帱�a�7J���Zb����$:$�K,��/1]b��D��$�%�/1Nb��>u�$2�?>$��Hl��"�ă��'��$>%q�č�I��X%�-�\b��t�a�6����7V�;�c�V^�x�婕%��E�Cĵ�]���E�l�\��_�~�,w�D�g=�����DC��+D+�?��ї<��נ~��U(>��n2�:���;@O������x��Kb̪)t���l��Jb�E�KtHL��&ӭ���Z�,�N�:�/�E���ޞ��9��)��W�+Qn}���YRW3L�Ќ��U��
��/�ji��fqU�GHy��=l.���q�'�K�7�8��
S�i��d[4���i_�I<k6s8-�)��tq����I<+��4F/	�<.o}|Lr'��Q�˝Bչ��M��gN�g�lt��ɍ�������ٹڑ#"���W:���;���\4��h<}R��gr�?c�o���g���K��*�gV���𦨛��������,Gv7r8o�_=�d�E�f�J�bXb�CI޴������vX�@�4�M�@Q��~�	H,�O�y:�������O�OO<�����˷/�%ߵ��J� G�v�z��TJ�%���诉�����M���^��f������_?3��q�N�#^����4Aԟ��roZ���{����0g�<����UP?�+ӟL�gg��y̬��O\����N�L�m*?�k�`0�i���;�櫼}`�~�EDɴ��d5�\i`��o�/d�l� ��2ҘC8��R��e��{+��+�_�o���L�Wx\]�Ŧ.ɶa<��1y&�3f�/ h>Nl��+�[_�x�Zf�l�4X�]�"*���4$�ᴻ�);��@��v�d�g�$An�"��%����U�TZ�h{j���Pb>�YT�YF �t�N�Ab:��E>�R_.�ew��cǹt]���~u�����l�؀�&��J��������1vY���L˫G�t�G�^���j��D�*뢝;�ǁ�����J����;����Nf�u./����Δ�*�;���f�8�w.?8A'dK9�l�Y��R�?c2%[��f���k�Ww����}�����t7�h���D��u�jS��R�=�O��g�=��胣�t��B���3��"�)�`�TǾre�[=.����e��,.~�di�'�h�\�i�k��]N�u5>0v[�<U5��5��u*�]��ۛϧ.�R�S�A��\��fno4�m����Ώ�V�$�3���v�[O���)�/9�
�&��f鍆�9�y��,�����>з�LZx�¤���:~f^�%@W�HN|�u�T�lz�y�٪���-t���2Ki�w.�myු������XfA����z�ݲ~I�jӻ�K��=h��Mj���ȗ�3G��䪒�}��M�ϛ����%�h��O�#��MgNfaf�1�vW�3|����;aNy��~�5�f������=����%���t�޵p�Z�[O�y�r��,�Az��>M��dg�tޯ`y ��B�~oKz��d��m`�n���\�xϬ�5����}�q��T��?�Z�K�Z�J���-�ީ:�4&)Z�*�K���]����@a�էOٹ�d�zn��NDuu�W��B�VG-a�s��GtV��p�
N�s=u��v�ÿ��%�����Bn�*)E0�JP?��
NB�,~R����H�ʏc�鋟�L��O�?=�c�ȓ������ʷ��'�2�Ҏ���9OG���*onŹ�Bp�q_�%�<f�wf�_b����i+<.nj%v�%�[�&-��Tɏ�@�����e���
�5����U��y�����Jy���8��zx+k�S�\u7Ol�7�<O_�-�J{�������k���/�O+�uy��3kt�25�w���J��K��
-��,W�1ϳ�2!����S���fz/8t*T����ԩS�� �gb/�v�Ɛt��@/��{�ם~o�;���{�7�5w�in���;l�+CoJ!��_|c��#y�����v������,��~��!7�J8�*��;޾=�o��gm�?����_���Ϧ��V�S٧W�=�n����կ\��m[��,���Ik�u�,��냛>��N\���~V����5~��?c?t��O����xb�ѯ�=���e��T�񖾍�mL��aF�:��g�u��W�r�N?��Ii��|����-Y0u�����o�wjAcۃ����7�oz�yu�^P��{�����g�?���j[�+�ܩ�!��x�hU�����Ӯ��v��~NN�gN�h��;m�W�s�KG�Q>�;��7�>�9f���^���-_MKo�a�n����ם�6q���������봽?��iu�%>6m|�e��{q�퟽2��}�i��q/޽mڇ��[?)���Z?m�ȗ?��\�Sݲi�K.�s����?�p��_�_��k�`�6j���6����[Ϟv�#�e^>���K.(�*��Ȣ%�Nݲb�-�ONXV::cB�#SFԾ����;w���N{�f�n�㭟^�������w��9��q�'^9�������^7oR��/6�yw������?)�ߖ���>{���cc�K�U���G�|iئ��^�C�����kͼ9�Lٝ�����Ԓ�Vݼ-|��������7�������~���W,cw�g,�%�m�X<�z��A���n໠�g��� �1p��M�6�g��%`XA8�y	"<�h;d� ��b@�;��~���0�G^�Ӡ��
�;j�i�-'9�m�+B�������p�g2���MA'�Je��j��I�!���t� ��,����@��"�	_�n.�i�τ l%�M�(n���ы�
7}�2�y��e��7;R d��}�C���-.��}�� %���KЄ�I����f�(�i/���B�6a�p�7��9B��ڋ���a	�ǝ
ǧ@_��L��t܄��3���gm�:�6�.�	o�\��`¹&�n�?�R����.AٞR�"&\�;�0�	o}Cv�w&���!��2�n�:P5܄kio9���J&,Z����P=���%��YQ~�	i���	m�Q$�o/g�Tc5p^������sYS����7���p��M���\)tE�Ž��mОk	�K���v�n�#��v�i��wA����΢}��}�<�g9ܴ���?9��g����{܄��p�����?�P��;���=�A��&ґ}׀b��1���I�{��D��}�m�����'h5��Bħ�"�i_�W���i?�yKa'O+|߽�e�-��ۭ�=�N���M���� 7�i��
nګ���'�}�F\Yp���]#���m��
�o1��i���p�>9��n�#�v�n��϶��/T��y)+1&��+�|���U���w�<�A�iO�/��i?�sW���}_]-�'�a��A)pӾ�ø7�g���.����� �i�ę5B��#�ᴇ`&�n�W��Z�C�Ҟ�Y'��7�U�����G����
�[�/�]pӞ�Gn�~�������M{3λI�8�f�
�W�4nګ��u(�ڏq�n�˰�-�y�i��so�~��/�v7���mB>�A��z16n�]�/=�t��C��w�3�h|�?s��L.B�{�&���n�ɠ�pߍ>rl��q��1/�(݄�������c��)[�r��������m.�/����8�!�Gp�<D��	��5�`<B8��GD��+<n࿶a� ��m�q�I���q�O�/>���M�����࣠*��ہÞ���&�o�~Z���O��;�g�~>
�u�h;D����L�����"��/���=+ʰ��s�#���{N��G���?�~�����:���K�����r������"�>����w��)/`c�H�x�I�o��#����c���	�H�[�+��OA������O���6`�K­�b�_\���;���	w:���h�g�,�.~y ��ۀ�^Ř7��D����J{ �y��s�����!�n^|H�������m��(/`�fQ�X็ѷ�
��_�qX���\��(�>x�Ǿ���$�
��r�o���;(	�o�K�$l�
��c�p� },���#>������M��/Q~�o.m�~Ho���	ݶ�C�*�ׯQG�?�e��(��aM�z�����a�
����"�w��<)�p��w����O:p�H�8����p:~�/����
lQ`w�ԅ(\>��P����0��p��Z�����ѿ�~���.�)�}��G��I��@M�����r��Gal{\�j՗�_4��	���q@������V�� ���׃P'�3X�����O/����	(���D}Ӂ�	�������\�E^���C���7AI?
<0L�}����>�$������z�(s��:����3���Qm~+�'��������r�m����i��L��1��W��v���t�:.�%Ap���h!̜ �wNT��E^,Ea���l :��f���nGS��ږ����:R��A�P��2I��A���h��ߘ,��\8c�O�N��p�4��ip(~?��=M�Qpy�(3�z��i�a(�������F���	*��7p��ܙ
����	x����%�z��Y;���5p��u�@5�v�Q�	�n��	��ø��A��8o�����B?V`���=
Xv���j�ۅ@��+���})��<2��}��e��w��_��D�m �Z �|����ܭ��
���ŢM �7�N�X\�6�/��}n3p�M�ˁ�%@
��z�� ��հM*��偪�N�t�z������
|H����W���M��r:c�܄c�����&���'\!�	��OJ7�!�&�L�����n:�� ݄��M�\�	�Y�C��t�yd?��X���Zy5�M�O��i�|�c5���캠V���d7I7��u�V���R�ni�(�t�yO�H7��Y�����S�'�t��C�����{��_�O/�,N�e$uNߑd�5��0T�c"�M1�\jE�u����jsM=��Mv���&��
K���ǖ�+&�\�*'���0�,e��-_�zƄqIg\��Oq;=.~>F�M�ҥ�z��R�G�S�҃\Ts��Ri���T�7�?:�
I�D9�����S�0��m�������b(��&��Qf���3.�2��ľ��w����e�2�[i�����yA�!�`4f�]8w�t�?�Em�����@}K}k�����[ԍ�8S�a���~�c<���6?����Y��>�>�^_�X�T�Z�^�U�_?������Q_U_]_S��~C����������wxm�'�Y��!�!�AߐؐԐڐސ�P��hHܒ�e��-U[j�lزu��-����u��-���[��n��:wk�֪�5[7lݺu�֝[�-~��1ݶ�mY�ʷm�ִ����m�lk�ֶ��PCX��[�0�a.JY�rV5T7�4�k�а�ak����M��ihihmhk�m�oJܔ�)uS���M���n*�T��jS����-�[7�m>��5�c�����I����Y���s���U�Ս5����������� PK
    +Q�H�^���  
  &  org/bridj/objc/FoundationLibrary.class  
      �      �U]SU~N�d�4�� Z+"Z �-�6i,l�S�M�Z�q6�i8�2����Wz鍷�δ���eg��߳��Фh.����}ޏ�7������0������T�kf�iɺ�GEյ�#�at�~j�M[6���}^�5DR}��J�a���jKi�����v����i������'����e_�rw!}�Ζ|W�F��k8�0֧�a��v�(���|HoʚS�s�d
�΁a�O�t�$'5\ꗗ�k��@xq��<�*��]���&���\VH���s�SxOG�3��=�1���)T��Nh���	o���d��+���`mv��)����+��a�Pv�Kad��s��d���`��b��/��[��,>����4'-����0�	A)��g��M+<5,0hOw�>�v.��]�mK:�XfH�@� �i����w�A1p+:.�3��#���A����l��C����jDFܯ�MQo7�Fh��M�R��퇘���m�8I��(Hpx���&E�f�_�}{ ;�ɑ�p��lt��j��k�Ӟչ'\^?�T�m��k�kt|�-��F٠"ywyCx���m�(�p��`�R��T�P�I̢�Tp��ݬخP�VV�Z�o���ߐ/���\��˒]�hv������}��]���3V��lvl����֥t�`ǩ2��@h�کo���;;������(H�ݠ[j��N�ד>�����F�^�Q���-Q$���C�}��N�N�,�z����(3x&���W��<P-���� W�,#|��%W�MZ�
љ��1�.��1��I�"�B��Tcc��&�a����>C"���čǯ��7K�_"��d*z�ܽPa�Ga�7�қ=�Kܡs�X'�ֆp[t��6��s�8
D
*ӛdq�`dH�%��`c�'�� Ɠ�����د�E��1v�h��A&i��5��
Q���!|O�NZ�$�L��$���G���R��/PK
    +Q�H�k`�A  (    org/bridj/objc/IMP.class  (      A      uPMO�@}C�@EP�*z0�(~�.&&4$�-lp	�d-&�,O$��(��B��&3��y3ۯ�O �8##5�J�&�(����4�������u#�B�a2,����>�n�P�-B���9�H;H"�@�,_�����s!��<��G��Xy�W�`�c�ۺf��f�<�.	~`'�Ӂ��LE_B�#C�B�wS�O^ٞ�~�P\Wv��W��-�P�˩���� �O8��ւ��k�Kd�����(�.9�s�˵c�*R��W��ګ��t�.�8�^�?^�(q�1�9�+���~���81�T�95U�PK
    +Q�H��E}    &  org/bridj/objc/NSAutoreleasePool.class        }      �QMK�@}kS���U?�g� m�bT� �+��&]ꖸ�Mş�I���G��TTPp!3��{o^f��_^`�������=C��=I�6"<����/�e0�- ǰ���?�#N,��ƕ�|n��#%��=׉�s+�b�lI%�1C���Q�����coḛ��畔%�o��莖�
��.iV�F��f�q�/
X��FdL�2�R�X&�3�'�_�<�q#y��4��/�h'w�0��RW�����/;����,�]��P��T�z�(+�DOƒ��(�m��;��u��K�Gq��<ʌr����#�R,�����5z&��+asT�g���y��|��0>�3VRM�)��ȡI�f��c��!R�B��PK
    +Q�H�c%��  �    org/bridj/objc/NSCalendar.class  �      �      �R]kA=�l�6i��Zcjߚ�m(K�F�>�;�7�30;[�g��������M�	���c�s��a~����]���� �����`<ʅ҉�����|ȦbWAQ������+)��R� ��J��@�J.2%��L�GF��ɝ
{�j�}x�x�3�����e3άU��>�9�m0>�N��V���KO�\ċ���5���
qݪ�ܠ��\�c<aaC����p˩�$����;��V��2RvuR��LK�YΏ��6�ǀ�,���&Β�-)��d6V#���3��RM)%V�Vk�o��
���� �g��w'�R�_9)�;q{�-ls|��s%�F�EM<`Dg����pc�U��\����c7�/6��Q�K����8�Qf���� PK
    +Q�H�ܞ��    !  org/bridj/objc/NSDictionary.class        �      �W�We���e`wLW��� ��&����\TK�]�ep��vR��Vv�����/~�/y���s����;�,��hvN��3�>�s�=����ׯ�x
?
�Z�T<�5Ƨ�Vb*:l$m�2��EB`S�`bJO�
|�ٛ��YM�F��3����k��#�-5֔l(�8��6�4�v_�~XEj~��ۓFN`K�
n�j����ө-+b?n��g�{�T�	fQ2��fL�q�G�:��n��1�']��R�eoX`�x��Þ촸cڹ��.#��(�^45�8���ҶJ�=�F2��)�8gu��<� θ��؂HUx���q)�*�NK���f�y"3�+o!���xgZ��}T�;B؆:�J]Đθ���<$��Ob�t#VRL�R�@Y��4��
l,���ө�Ma�F3�-�W�G@��r��FU<��a��>��t�u;q��Q�~�H�,f�T�*I
��uKCv�0S
�غ�����&�3Y�1E ���R�=�S�:Bx�''��+�[�g@G�%A9��2�a�`*zܐz��%k�yV_}!
�]h*��bֻx<�Ai���(�'����c����|T�͵�n�RBz�����U3Lܴ�a�Jޯ�˺�1��q�(�b�t��me�r;�R�w�w��0h����+̀�9���%"D�G�U��"���䴭~��Ү�:Ul@DJ����v0Ul�&�&�,i��r��i�!'O�H�׳\S���̲\mk�OJ{5������K#3æ8+׸�.yoʉ�U��'H� �{"�
8h�V����Z
ƥ_VN�ʶd:�]���W�����)#Gu*�ʳ�#|̒���xu�~zX�Z"���Y�L'8�\JՐ�25{&��sG�J�z��s�J��6p�VիA��e$��l�����$`�Ľ��XZ�3�u������@��}h&�n������T�!k&�����c�zֹ��9N�
���_B^������|����/���g|�.k���k���.���Nqʣ��;�_p]S���k����\(пUx���k�yM(���,�!�/:&iI!=۰�'x�W�k米�}���I�X@\�5,��8$����5��_��&���8<���<�$���$^������D�C?Ӫ��B���	�0� v�#x�Y�W8��|+8���2cx�8�W�}�k�_>F;�W~\'o߮������ە+H�Q��ⳋ6�������x�:�p��yݚ� =8����`�ڜRʅ6�0��9wP��p8���h�C9�W�WS4���A=��g�0] �r�ihl�ë��;sv�߷?	���#M���9�v�Z��K�J�:�Ysx=��E�D8�84���a�r� ݎ��"8I�-؃w�� :Q�����n'��L����L5��3�W��}�v��[��>���\���QJ�|53{`����'����N+�)�B�:�%��4&�y��q|P�ǭp����D��(j�8-���G.��^
	{(X�PK
    +Q�H�L   ^  !  org/bridj/objc/NSInvocation.class  ^             �S]OA=��)�" 
(��1�F��$�J�jf��:M;���6��x����G���Rꊛ��{g�=s�ɝ���� ����v뎖�A�s��E�L��7�S0��� ��@�LI��Y�ဏ9%�n3�R��t4�_��c>C��T?�aXhH%M�!Y�v��!�G
���$}���=i�C*���Ju���"L��3��U�P�.�b�v�aX�����2BQ���'�r%bYJ:�n0�|��L���[���C��`mc�*�q,��}%L�U7�rѝ��6zÉ�K���i=��)�k�J�./b�j�;���קܕ�:�r-�3�v!��T�"9BOvr�*Nw��6N�����43'��5��w1b�'�*��VkF2�^�ȑ�J_R�m��H�X)τ�BӴ�K��x��Si{\��6C�$hB��K�s��d�t�+�7�$���b��X$�G�B�S�ǵ����l+�-���s_Q���4��ǈ��Eq5��-Tn��q����>�Ofcd�5meї��ݛ�a/lײ ����yi�!lW��PK
    +Q�HIU!  <  &  org/bridj/objc/NSMethodSignature.class  <      !      �S[o�0=.P�[o+]w����]�=��h�JCY�JŤ=L2���L�Ӎ���M{�؏��9P���)����>������;�b���k�9�~<�����ît�Q �`[7P��Xt)����1?��r.i\)ۑ���:C�{�`(��r-}ŰܐJ�&Cʪ�JȣP@E��ɐ���V+)�Ë��#���t�E۲���Ri�k	c��X�D��2t�M+���I_��V�F�t��fظ��cm�9v��ʧ1���
}�5K��{5�h�j'/Y<�D8B�zD���7�m��Om;�G4W��,�1�1�����6�����x y���!G*q�j>�_���9�ņc����r����f����O�I��M2:a��Hi9=J������v�y�2ի2�ܸK�+z��q(=�,ѵ4_��Rjw(�)2���(}���Ԗf�����ѿ��X+X���������K�7p���9g�)�����&�k�F1��׉T��E�̾�OTL�,.�@B�k���z{�p&�(��dC��PK
    +Q�H�]&�  �    org/bridj/objc/NSNumber.class  �      �      �T[OA��{�P@�
^�u�wQ��@JUJj�۴]�4ˎnwI�+�^|Q��W��̴쒰�a��9ߙ9�u����@oƤ�4j�h�YkՍr����L'6���2�nQ��c�|�p"�6�m�$jw�,2������w��.,	[����T5��i���s�D�a�t�Ψ������[��b��N�࿓�v5�?`nخ"n�bAz5�T�B8���%i7s3���EKr��b85�ޓ�[�t�zRaH�\�`HY�\٤���l*2�5���X�!Q�������������vd��gQw��LE�;ɕ����FG�0t*/�)�l�t��a�d�2���<��l3�Mcs�Ž4"0�d>���M
K.խ�ƲA�U7xL��m���S��'xF�[�SU�unU�#8�r�kAdK�6;��FRѴ����C5�t���UN�{�ɲWN�@{�)�W��2��ΝCKW���͢P�0��ٮ�7��-�VVl[���ic�t���`ꍡ�!�,#����7r"X�1�	�d��wAG�X�
��Rs�	a�ǯ_�%�&<�Q��e���:�+Po�U\��:nh{�N▶�q��[#L��q����u�)%;6����Gg~#�5={���X8�9ѡu���<P���C#��ús[H�L���F��N��Ŏ�\���,��h�<y�z�8�d���ڙh#�PK
    +Q�H�Q,N|  �    org/bridj/objc/NSObject.class  �      |      }P�N�@=�*�Pw ��HH���F���2�!0C�ք�bE��𣌷��d�sϽo�/� �8d�����lw�u|�y�u�,�1$)u5K'��������R�+=�����z��P0��u��<�Z1�u�d�`(��4�i�a.ʭV�N#�U�T�$$��C.�H��0�o�z�϶5�LgH�&
r��<�_�6m�s�ϻ-n$���!2����?K��R����	3��4��Ahȯ-��_�����C�k��CȞhɁ$�K�t_w�#$Hx�%��Kn��a��>�����D�laEkq��ulR���Id��]��quj(�3��)9�єS¨�:ck>���9�I='o?��p@�J�6���? PK
    +Q�H�~���  $    org/bridj/objc/NSString.class  $      �      �T]S�@=K)�|ʧ"���E��(�R�Zc+��ei�S6L�2��A} ��g���$�v�2v����9g��n�����s2�Yv����lX�r��d��-dQk�y�/�!��[�.�����:ڔ�H��mڗ�f���=�*OLWX�a��>��t�=���.Ϲ�n����R���*\�C(?`�N2�X��ˏ�`�Q>��V}�H,�nQ�(�6���9�b#:�e�%�0L�oIՆ�L�$S�`5~�0�D�' Ȏ�{d��"g�$��)��;����1���6 �ˌ�򐁑��Ve��kՎ�� ����H�a�����<��n�xJ寺��,2�{�RXF�d�w��?kxƠ�Zv�<��.�u�N[²N�����ݚ�t��4Fy�b���+Q�R�J�SJY'<�'�Si�4S4lE��~�xM��kpxʰ��6�W�<5�ſ�U
oTTo�zV��Vm���M�l6�w/]��M�a�Cu�U0+Ǧ-�|����П�g�gyjNE�ZU����z�H��T�t�nȧ�t�?� pRJ������(���w��Pߗz3���n������L3��3q����=�Q㘠��U�'-L���IZW;݉�L_�Q]d��D��,�.����r�yG$����!�+WX���@Ch]������R�+B:�W���ď��(�$v�J��I��+��FGs=��F�}
>�:��3I�$t��2�yH�A�PK
    +Q�H9�I  �    org/bridj/objc/ObjCBlock.class  �            }O�NA���DPP��d��H�����l��}fq�eǌ���'~�e�]T>]�S]������
��M�ƁtfVF*��Q�,�j�[�t9�J}�	;�v_ıjr����
�}T��qǑx��������kkrc�p�����,��ص�5�I{������%�k�L��;�@���'��3ND�9���qj�V�x(�2�79��I�e6��}2��͜��&��.J��O� Q��U	5�(����LP����3O���X��hb���l��z��? PK
    +Q�H��^�  �    org/bridj/objc/ObjCClass.class  �      �      uR]OSA=�ojE�"QP��<��km$�$��������Ͳk����œ��?�xn[�`�dgvf�Ι�ٟ��� �
�ΏۑףI�E���1��zF&IB�� ʭ�PF^`��?��R���V��|�5���rT
�\'����u���5[�N��Ay�V}yΚn�(Â\)^J�*�*P�6	��*9U�ggGgN`����w�N���5�H�s7:t^`o1�����	�+��������C�{5�	������6�UύXq��bi��ku�	f�k��ӋH��gi��V����z�;u��ld���8Mm�j�͌o�uA�,�S����P���qr�*Ad��ܢզ�Ž�X��!�ǔ��Uܡ~2��0��]�����˴s�6��;�{%�*u�G��`��
ް�`�
��(#S�*/��Kz�MPK
    +Q�HR�o3�   �   !  org/bridj/objc/ObjCDelegate.class  �       �       ;�o�>CNF���t���̔,����d}��,g�Ԝ��ĒTvFF��ĲD��ļt�\jr	;3#�<B�_bIfY*D�3�$�(-1����A�0=�9�\���Eɩn�9�l�L,�l ���$��PK
    +Q�H�@�|  �    org/bridj/objc/ObjCJNI.class  �      |      �QMO�@}C ��B ��pI@������R��
�3
�.ڬ�Y=U�?�?�b�X��`igv�{������ G�L�[7B�����(�
G��ˋ�P�'��S�#_B�P�%�)K(�����Ph4�Q*c��y�Ǆ���
-B-r�<�@���=fG�"2A����Ym<;�S�N=�GǑd�;-p���V����D^[��K��N�C�4d�*�OTu�OSM���N�	�]����Va��SCX�j×�C�.G���K7zh�O���7u�`�|��ֱ��}�����Z*5�z��$+)���E|�c��ɺ�o�nO솼�����S.s�[��(cY|]N1C��)��1K��Elc'W� ��*��_��:j�˿��/PK
    +Q�Hv=�w  c    org/bridj/objc/ObjCObject.class  c      w      �V[S�V�dcL�	�PJ/$M[cizť.�$撘�$�ie�`�%W���������δ�>u�?��]IHF��0�tv��{�ݳ�?���'�Y<S0fZ�BՒ�݂Y��k����ICQp5�^��'���
C��]mOS0Z�5�(<h�l�9�=��
��O�#.��=��َ�����H�Q0���0[7�����mǒF}��_�nɖ#M�\w4{GA2;�� -�ş�Z�Κ�A�|��O���Q[�V����hV���б���l{Uk���+�E�:c	�e5{�$��ѣU�n�M�옵%�R����*�W��閰�M��`�\��%����t��b�k+�h�;�|ȵn!���[��ϟU�M��ͨ����/��[�-!���w3��{܋;ҦWK*��i�b�G��)���#P�A�8�M��3)�͌��4��ۺcZ��P
�n�f�)��g�ZǬ�w�z�.Ih�i�T\��A���V�QO�F�2�'��GR1�/2�_�A"�^�x��XP�>Π��(�V<��V9vw��|Mm��1\���P�>���ٳ��U*������2���UJ���P�3]��1�8�>�9%�&T�� eQo��<�/��n�Ҿ%��&t��Y�GDE��i[4�n�M��R������c�Ή�?�+��s� t�#|өn�V1�	-t9V��L�G� ��=\j�S���%�jCl����I%}�����4�j�?�f�<�#��_�b�-],I󿪛Җ�x�0LG㯠M�%A�P��2��~?T�|GRߓ<�!?%�bD�f�P�[� y8"_��#��C#"��5w���q��k$����J�ۘd�V�p�V5�7��������? )	Aϫ����y5�<yo�Zu�aM�Vuw��ebkŏ��F��'G�����a��5P������x`��J�;��:�l1ᩃ<Ӹ�F��m|HV!�z��h������;c�C|Z���>Z̕���C,�!d����-� ��|�2�6�c�>!R��9���7t/�Mh��h�/$~E*������������7�o�ȹ�^7�D���y���K@'j�@�v�"�I/�BP�C<�������&���s�_�l�%$9G	sZ��La���d�8i}�PK
    +Q�H(��,  �    org/bridj/objc/ObjCProxy.class  �      ,      �X	x�y~?;��J�%KxmL�`�j����W����.,��׻ci�jw�];mBh iZz$!i M�҂ۦM�"�9�aH��дM��mz�-=Җ������v�ӧ�x5������w�s�_>�z�
�e�������Jt���2'NjA�c���D^C��٥^;?�9s"��XFN�h@-v���T�`<�#8Q��;0��莁��5�n$nZU�C��F~2�-��q8���n�8����I�V�/Xl��g�I�ŭ	#/h);�E������o����6::>�mpG%�h�2�$np���Iк:��������ŏ���@	|�f��oԆ;�	��e�d�tްz:���:�T������$���]����Ak@���G����h��*%,#�7\=G�t��;�%���P-���.+�em��dW���� a�z�����ea��!�K�_d�,s��HVt��D�-mn+�w�ee,kut+g4@WҮ�z�I�<�/l c���
Kc<�$M>�Ȥ�QB��B�t��wff��'FV��FƯ�=btF�y��9,^r<�ۋ�t�0
U[G#��F�ޙtޜ64�����8]2*�<Oi�ѧcn\1_��3f*�,کc�1�B~�!��٬�&��xڶ ;ʼ�� Jg�cʱ�U~1�L�eK��Lx�6�U�GU�lֱ���W��C�~��m8� %��xE�;����C�a��b��J��eP����7Y	B�L��Bْ���b�e[��1���KǧZ�u5��Z��./��J^m"����SU�*=�V��ӕeug�5T1�X���k/�0y(ũ���%v��w��}ti�i���q��N����aJ��|EE���(��t��GO�ޤ��	�T�:7g0,K��Q�&Q:�����YO_�C�Sc�V�^�}4�/h��>@�l\�U��xl���Df:;�7�C���`�ٓDp����~J	�i��R�D��Z��/��V(W�*3�g��iյ磪z|LP#��s�)yz;�5����P�G�(m1���#xT�'�)��O�zrȨF��_h��KB ��J�g����׹|<�`^�wzT�ʞ@����m���4���NhY8V�;/� ~����uG�R�X^��g��<~S)u�bTpv5<�nb�3W�̳oӻ_�_�,�P�9��S�]�8:3�95�|OV-�&�	�Y�C7�:���i���3},���@����R�~��SW����Y�\�������c'���%Մ_��*	�T��;Wzf��a�fM�L�|Ξ+�x�(�W���WS1<U�B÷�JøEh��D��[�a�y�w�m����ǓE�\�6s��|b�>�˄�]g(���b��U?�p�ȳpi��漢�Ǭo�f.�x$;��TuP3�v�?�T���_ҫ��nӰ�Vb��;?\�2����)V����1��飫߹�mi���O�L����(���s��q�Z-X�6�G���&�pܪ1�Pc�=��.�r;��o
�^��`����C���Ȓ8�e��L��d+�L��+��
��a�^#BƉ<�EP���2�p�	�Q	��	����*ꪻ[#��[�ҠD�W�����b�9��W�_5	�EZuY"��5�E2�I'�nO*ru*9n~���e9�QVT�F�Aeϰ&+�[ނ~�8�ڃ�K����<<�R�v�����j��UJV;sg�@��٪��	��^v?3]���)^�r<�HLw�E"=|HD�KY��O������:r��fY+݊ݺ
��5��i壀�W�|]n4���˘IM6R���#;�Yd��h�����Ae?!��w�ݾxj��n���v����B���cVf�b�!Y?(���c<����Tޭd;Ua���-��E�Z�mn\v�YE����a�>0�̟IKQ�
� f����>WW�bo��*%�.�WM����hs��n��c1TXk̖��z/~o��6k�,��m�	K6�A[�L���Ilz� Z=0K��&R��F�I#gZF���1�g�q�����娪�,eW����=�m�QX_&i�Y�8�/n�*�cq;��ic�+
+�dԷ����[���+�e\{���˿��/R=J�;!B}��G33V����*Nu��X}�����.��� ���Ј ׏��͋��/c|V�����;|ˡ¿#rm�s���Y�`E$2�Ugp��xK#�X�R�ϡ��.D"g����7�߀�7`�V|^N���z���Tg#���O�I��o�'�@��{[u=W&��Bv�sޑm?)H���=Ԣ�DM�R�Mԥ���;t�r瑮9�<����p�9l9x�(swK�,����e�?�;�}Z��pphMtw>��9����"uB�4�$/(�km�#�<W�#0l/�q �pmZO�'�T+S+��	wo�{�ʫ ���v��C;H��v��8���6Pص��Cj���|SQ��|	�O�e}Y(}�� �F��i*Q˿���*wir
M�Y�\Ľs��Ӯ�!�е4��{�̇V��'é�Xg�>��6PU\G�z�nI��HTx�|���������5�K��U)����g��ދ>�����S�v���8z��|X�h�~~�4iA]���PE)����mʰk�p��f:��g�h�u�$p;W����� ��!J��r� �;1�#3���ᢙ�
�7q�M��K�s85���|��o��u�7��n������`]�o}L[�f�?�g@�>���_�5<�gA���]m<���Ԡ��5�sxn��N��f�͋x!��Y��R�flnloT�~���?��r��e�GE�蟃u0���������[��3V��_����h�������:�C�ނѷ������?����C���bͻ���殟��,���09��4��FO.�Y�;~@|����?��
ěnD�,D��T*!k(��'���j������c�1��&�������pcw?2�)���=��*�"i_Ž�tҍ�_]�
���B>�E��Y�S��m�|�-5��QSu�U|����q� ԙSo��Ur��y}�K���[%`�S�i��8��^;���������*YĜ��X�9�o�u)@Ȓ�謴E�ì¡��/���$�.���/蛕+cZP;��������Mz�����Z��>�l��U�@00'�ƚ���6��ȃ��l��Xs��M6�>�0�}�&�S!��zb�26(6Oʖ'�n7�hP�nQ)!�DK�~J���O�7����U��|�U��}����;h�ge7K��$.�n�������7����= ��>(�,�MĆ&�tr3�O��}:ΠMn��F���b�Ƹ��c�,���^��>V ]���W�d?O����CDQ1�0\Kmސ�f����3�a|��	������ٱ�1w~@=xI�q4�ul+�+n-Z!C��h|kQcU�Ii"��#�>���:�<3��SMD�R��U����o�3�z��}w��BI_ev}���:3�<���=O�\�?^ħ�>�o�����
�^�η�׸�;����ɱ4�rĝu:�>,i������N�����P]Y�Z]�o{l��PK
    +Q�H�́��  �  (  org/bridj/objc/ObjectiveCRuntime$1.class  �      �      �R�OA���n{�-V�_�U
$���Mh* }��n�-�.ٻ���E��Q���5�afvg�������s��.�	k���Ȫ�00�0~DCgj,['#���� ��0�A�~�"P �ܡ��ҙ����0�V`�P���v<���dʄ�z�P��A(}TZe���F��C<�P���TJht��A�)#O��̈lt��/�c�4Y���1��	Cf%Z�C�g�����$&>�ɚm7�s�𰂗�$���ʭ-�㙪�I7�*�y�a���<]D���Ԍl,��I����*��.����C��m%a��;��E��#̱�����OG�8�y�ūIy��?Mb	U�o�J.C�װ��?s��+o������ק��N���(���A�>
hL0�8Qa����3;d��*PK
    +Q�H_�Q�7  4  *  org/bridj/objc/ObjectiveCRuntime$2$1.class  4      7      �Smo�P~ ��^Da�t�Y`2�ݲ2�#��f�懶ܰ�]KJ!�e��?�e<��L��֤�����y�s����� �xF�=�S�|��V<�kW�Y]ar(j{7��B_ӫ���C��ng�%N�w=�����#̾�5\"�&Wa�|aS��te MG~�y�q��4|Է^l���e��!WS'���t��mf�uB<8�}��ߦq�G��P7	/��4�����`6�r)d1��넨�*s($�<!���. �Wٙ�^��`�GvA��q���
��X���]�r��'�j�掆�|*�j���٥QW�E��0P&P�9&�7J��1V��lp��٦�2}iZ�x�B�!]�Z�����}�@������<��*�b��Ӿ7�m�-C�W��x}�vފ��kR;�+��c�����<�xd�j. G��=��p��Ξ�s�c�T>µ���o��%>�5�@.�&n����wh�ׅPH�|�	i�"���1��cY�DC�ܨ<�Q�
�"��%��UΔDZy�mh�iz����G��8�4<�C�{�rV�J�+2�qf�� PK
    +Q�Hx��r  �  (  org/bridj/objc/ObjectiveCRuntime$2.class  �      r      �W�_W�.,;�]%m�%���k�<H�h�d�R�l�;;;����:;$}����~����o�6mR5V��+�	����X ���ܽ��s�s�wν����~@�#p��LG�������Y=:��5tל3b9�5��~B��ъ`y)���1�֔=�Hس�����zf�9M@��E��i�-�����ѴfMGc*�Q�<�^��#%4�̓A4! ���p���@�F�|H�)Vt�6V���R�S�����"v�6-�p�F�в��`�����I%!�;cfýL��v^2w�!�2݃F��4؍=M����H�l��.����$x�g[,�~��[��wn�Y  }3��y��]kL��
Z	A`Ǻ�(� 3Ӳ�iMW�ǭX�q�M�8�����?D��Dm;���'���h�tRӟ��<Ni:��OԚ�Y���҉�I���D�1����� q�DΔ��)�q<�Ķ1 ��O�dty$�!<@װ����X\�!�Pg�\��3�;3���m�0���b�Q��0�a쓴��@K� ���R$���VPq%�	�����J��PR��� �1&��3���l�Q��M0��'%��J��d�'?X�����M�'pJf���e�eF3zR�㎡-�%��?��U�����3�Ѵ��f�,�zN��]S�2������v���Z6� Y	koo���t]��O�j���M����YU�P+���1��sV�؂nd$�0*M���:���-$�yX��v�~I��?XC.h�M��N�~[eCQG֜�������w$g�S����#�� pQ�}X3�FJum��A-�뎩�D�Nَ*�W�i�e2��~�]}���&�	�<+->�.��_/�Ҙv�̺-�Q����x�#]�0�+rr_����W��k<g4���MF����,�2`D�U�>A|ߐb�$�,c>,q���m|' ���yA��שGwA|Oʿ��쫘=ees���Fj<c8��xU�Hj$Ə��3��J�n�\����NV�ۈpYF����e-�Y��EƦʑ��J^��J4Xb8*N�\3=��s��-.v5��
~�/�+�Y��߬cV�P�d��$	�t� A��z{^K�K��?Hf�% t6�]��F�S�ú7F�n�k[��MdzorW�5cA^��V�l�J|��*⤕�L��;k4A.��+�u�ֵ�i�1e���j5-c,w>�C�0�k�S[\h:iN[��s8�Gx@����MZ~�\۬/N�9G7�M�1KO�Y&�����t*�,��b`d���6���hi��X�|�܅C�/B=��`G�U��]˸�
���|��k�#�7��8�7��� 1�'�Y�Im��-���
��c��]�]¡���v^��|�8�}]W1ؕ�C+8ƥ�W0:ֽ�����䘷�{g���ѹ��%4zo���C�A;!��Q<@۽���Hzr���,��q���ʵ��ce�O���3��>���t~���!��a�1^l���/j��y�9�3b�"�����bD��~	;<g�V0��&/�3/Ԃdq[���g7����Z	g���8�_�g��q�L����l�x�r
�%~2+p|!�{�bnr��x���<���y|��<���/]�Z�<�6�j��[��/��{�.cg��ͼ���Kh^����/�'�<gC��t	��j#?+a��Q�o����=ͅ|˸z�禃���L��6�@����>~ +5�ێ�9�c����n���r��y$^�u�K�7��)�].��cY�*�t��}��9Rb�b������'yM~
��3���/��o/�M�r1%���¨�{o?��b#��oO��Q�5�؁�o�m���D��o�?PK
    +Q�Hx�?�6  >9  &  org/bridj/objc/ObjectiveCRuntime.class  >9      6      �Zy|����&�� $��`��E8�&�@�$���f+����b/�jkm��-�jK[�a��.A�b���Okﻵ����������fw������=��y��x�'���#D�D��)h$v4$��767F�7ܨGR��z���x*:���L�.��^�43|э��a����x��+:�'�ژJw�c�:SM�h2���r��5��0fZp6�j���;�%*�3�r�6�xJO�n�cz8�'T��4=o_�iL�P��z�rC�z�v�h46(*�R1(�f0�6(S(_���zj�1���:�C�����[L�\,k�{uS�؈.�*͂�
�4�e ���Io{,�L�ɵc�d{Oxj��%
mMEc���(�/we�5���;�{S�h|G[W�<W6t����W�*��i�E�"#��ф�vL�fZU���>�fl�Zo�N�# Ǽ�"�m\қ�̴�8N�lLW4�*z���L��m>��n��� �鲲6fDv��;'_���HU���HE�x�h2<��xSy4�fw8�%��Pݶ�@�)N�a��aK�dw8���:���"?-��L���hnZ��\?e+��hj�y��Z�R?y�2��iC8��R��Omt�F�(�#���h�5�R�K�����W��&�К�ШC�A	�H���#�l]�~��j�hu
�s\�ф)w�����T�l�!��P�Rm��m�h]SNi�I_8�N����5�V7���mߡ�L6,S�QfM�-���C�t	��Ա7�����KX�3�#rK0�k����(<�7h����{�	B�m���K�t=mg���ӌP]>�Fa�SEr�mZ�+0]\H��K��4DQ�|�ϩ��q��Nx�S\���zi��Ȉ���
�d�	J
:�#�'��`�Z�����
F��4�9�����m�jc�5M�,(�Ƃ�R/���S;�d<h�(h18��K�aq)âD��"�8�A���,!15�&ƣ�//���v^�(j�*��I�BRK�;c���/�E�L��"~�XJ7Q0`+�u�XU�y�_D�<I�uHX�͚O�̝��7�j����x2�G`�u����B��+)�6�d�"s٦��2"F�[w!<�k/*Cj��	=9b��}F�.f �ԟ�)�ގ.OER�mϘ��
�� ��7�6�{MAIUZ�G��U	,
H�T��b�*�Bq�z=�'���:n�[5̬�ЖS=ht�������=�	UȰ��2;Tw}q���L��1��/u��!���M��DqIA� ]�e�vvQR��5��'|uK�}�h��Ī#95IF�*c򍈰,I��UJ8��E�**���8@�S��D���5��}	LB�EVu�(�@m��c��3�]��O#R�Q����F��3~�=��6�+n�A����l��t��$���>��xN�8汗>/}��-V�����}�O���H]h
��`yͤ!e���P{qEٰ���a����!�;�v\�}��+d|�ijn!��2Z1��$�1k�~zZ�|��(2�eʊs,4~L?�B��eĈ���xR��K���B~P�@0$Ԫ�)˨|�_!
<���7KS��v��̩�ۻ�����vn���Ot�G�ҟ���E��f�h�Y�}����t�����5�}S���2�	މ�C���>�=�S~��4)���
=�ƞϹI��ʥ>.��,�k�M\e��}p��a�,��&;��U�(����xڄ���A����R6<��2�6\Qҿ펡�޶��&8�={��:c4>�V׌����!�B��lD^���p,��\���s�B �v��͗�>������x�Fw��?�j�&kt�F���PN�[�i;	#�r���A.t�I�=���%�p��k��/��'n�A2	���#Vΰ�I��hB*V|�oL�G��΍YbmA,�l�������TnE�����PX����]	;���)�{%_���H��rn�հ�l�T^�4��;�Rh8CA�:��{�Įd���Bųh(���u~n��P{W6�I��r�DK�W�hpF3��{��uM*9�|F^�\/!�, ����-V��C�\ô�x�aG�^���	��:�)A���n�5ކ���z�E��b	�p�u	cX:�|}n������v� z��#� $��ك�x@��,�B9T�f`j.�v,��F��s��&�1���7���U�K,�BlP����/k�X*M������������V�{7{Ѡ&�FS;�t��z�wKp�#*��;y�S�1�Y6^^��I;��uv*	��JG�7]��	�����.X������ ��˷!�'��XX�����u!μ�o��� ���6��l��������hV����@Q)^�?r���l������;�.��7#��GFb0��I;y.N���6?��ۭ��mF��zi�P8�qwΛ��نS���+`��9�ϞP�X�~����c�C�����I=�~d�^e���Ka����N|&r�v�� �aQ��ty�#�}�?*;˹'W**���̄&�m=��E��?��G5�½@�q8`{ǆ���x��ps?����V�����Pq]�q>�*~B_F���5(h�^ȧ����T���k��4N���Lɏ���d��};�	��3�O��g���u[*ͅ]�)ЬN}�{zVqP)"�\�	�7法U�F �ש)�S,;��@�˂�{0b�p�O6����Vvp�~jC�^~��������Z�|��</�[��w��l>mgȭ�� ���j?�h�+g>�;���`p@���%V�h�(��y3����?�g����" \��4�;Y%z�>(7:LKϩ��}8������/pI>L�m*�
:�p����^���7UpR-xDD�-����G2��!�H�������Y����Jx�� 6y.�/�k�"9��P��yĲ(��_�$�9˧E(��|s��ko�����i��ΐ���?SF��=�:/������Idsޟ%��Ñ��L�.^����\���M[�ҟ&�Pvy:��d�@�_�����x�R@)CrۻX~� QL���s���~|f��Y��%zU2����K/�0|�2E�*�Nc�V"��.�K���d�L6��9�?\���we$f��9�'�	}��}��MjJ�|��)���/��2�O�|���z��
�s_�{�����Ãw�ND%��YY�uE�z��� 
dkef.��޸ve_�d$
����F]_�|_���
]�������9(��H?ԅ�Ϝ����n�&�ж�q�w��"���m�o��=9y��_�Y�x����NA���R�[w�vg�Ts^$��=N=P����&���P��j_x��FD�qn/�gU��|�NR!�����h"�[O;Zgũ�E�.��4������Q�X	b�`���d�k��3��|a��b�^�5a9���F�iMl�i 7���D�qZv��P�W��h9���E��+�᷅.��&��\]Q�.�?Em�'h�'h�;\�׎����E��'�W��G'\�"�Y���
Њ�7��*0r% Vc����I!�9@����S)i�����i�)�����'襏6�i�׮m:I7*t�b����q�H@NQ��7�i�	�U��O�n��O�^y�n9�%&�˭�,:�ѫ鵠����[1R�B��:z=��D�t;�A��A�X�q�o��@	����o;x�
���z�F(@/�n@��R�@t��\e!k�FښQ�r1�����6��s�[��!��7cd��
��0�?>zk�q�����p��Ngވ���.gބ��i�3[�Oﱭg�"7M�oH���߇���#�U̴6iO���Gq�5�Q�s?��������jO��?MG�6�WV�����Q,ᑖҒ����҃4;�.[ڪ6�T��2>����6nv	یk�@9�'��4���ó��$�d<�!�Ĉ�:l�S8���8� �Fz��y]d���?�ߗQ%����+`���]��.��vI�}��ǝbV���ۺ?%�_%��D���l{f�/��7������np(�@_3)�Bm0ׯ�u�۰�:���C^�o�	�.��,:Y�Ռc��Y��}�������v��e?�Gl�Y	mm�iz��S�RZ]Z�9H�6U�.m-[�2� ��������K����Yn-�Ҟ8���\��&�ך
+��V�
�@am��Ŀ�5��d۠��������`�֎V���mA\L>�ލ�w�|=L|5�r�ܽ��8�b�ɄNn�]b
�<FQ�G��0yJ�*n*}���_r��������b�{��_Q{�I����uN����`�{��HfQ5����^�bN3�
s�;3�2���i���jώ�,7�O�'x�dSXK�F�!�B^:L�a
õwù�����}�������#����m�����n��Yi��O��}�G�_}�T�Y�Ӕ�
+�oh�ZKV(煇�+/��3T���Ӭ R`?�E���S���mB&���⚌U�"q$ۋ��р�M�@�2��#1����y	����R�E�9t3/3�.C�'ܴa�8,���k��YG�x�M� Ƒ.N��CH$��@>	3|���z1�3J���k����WXr&$T�Y9��������x�V4��5L=M��ݕC��@�x�=2%�a�_t����w�Ӑ�W��Y�t&՛�(A�#��f�Y�j=|�3c��k P��=�d�+}pO�/ ��_֯9l^j���;x�D����	�ݍ�[�{�� ��<������@���4o�*oiL�K�Q�F-c���9�PK�&�$��<�;L���p����t��
J�U&�%���V���;X�.��{��>������!"��(�~9��6�/P7���:)���E��%�Js�4�%���a&�S��i��T���iM%Mi~�g0ͷ��In}���M�R��,��4Ul�hM�=Mn֬�.r���9T��o�7��ٙ�)�����*}D�y���_�r�+ʡ�K������û��q�@���9ZyK�����L�ohl
x�������2����4�k������Z�����`�?�������|��Pe|_���z�x0�'�HM�ô�U�J�U���|��?�� ��h�	��G��B�����f�8>����}��~~�?	4�a��σ'Tݼ�����|�̩y�]#�"�,��2.1׾�5�9�
�4��5�:���%Ŗy??n&�Yεٝр�k}t����a�Ө�+��+���h��f����h���Y������8��#.%���ڦ8ߤ�g�2��=M��NV��A���o�O�]��W�]o*և�!j�X�c�m�H��nkf=��i��}e�!���K1�鍏Ql?u6>ƿ�Ok�"�m�*��[RU�3Y��AP���$���^��]u��#Ĭ�Eb�[Wp-M�p�PG�\�i��r#����~D����h�"����/v�����1�o�d�f�fd]���T��n�|�����4��Ei�b�ֲ�D�#/�,'E���(_e��u<�V_�����[�yJx�d�,����S~Vf���6_3��T~3U�[h&����;��[Q�U��6�V�!���~E�(�2�k�]��NO"x����6�JUD��R��EV��:�T �n"P�Ji%'���ߣ��T�6��-�ޤܚ�����g���$�r��ְ�$)�RI+�����8����3���2�i�'��ǕyG�@b�M�,����f/AMU���T�\*7�~?Y���_/Mř�e>��j`�!�zЖ����҅e>�2@��j�\M���PK
    +Q�H��$  |    org/bridj/objc/SEL.class  |      $      ��]OA��i��uE,XP�[d���D����6$zc�t,K�n]�$��(M�^�����������s�y�̙����+�qR�Wɖ<���uK����|B ��_|S��%�v|�%H2�Һ�e	t8ֆ$%�>�U˩d�g;�	��I۱�)�抎$�5t@��_�7��3��&�' ���I�Y��uX ^��n���L�� �ز�u��J�0Z���u������F���gG�8�!�c�����u���[2�\w|{C&0��6e��'+�&��"�m��N���8��N�����٪VG�Tv^��ڳ�o����.`DmgnYN #�UM�E��0�1v���)�@���u�ZV�y�Fx�W4v�U�)�Us=#��l5�V�NY`���M�7qK!o�8�D��{fwud�c�H���V�{d/=��	�/�y�r:fp_�<$���D�T���\˹eqN��U���Нʻ�Vu��l�T�Ee�mG.�7Jl�Г��-t�c�u��mH�s�-�uoU��U�3�C� ��;8�_�z��O�5�8@W��.��,��4Gz�� �zp�9��k���N���ߊ��1�ʌ�"�X���p��K��CO�>�E���,гL�iD��pT9��'��3��CV2:�b�U�˴l�(���;�����ɐc���G+O3n ��p=A��)��z�����C_0�|�R7vp'��I�)�L7����C���쵈Y�
:8����o+��7���v�u6J<�Gx4T=M�3,d�^vfK1b~��lV���Du�PK
    +Q�Hڄ��   C    org/bridj/objc/Selector.class  C      �       �P�JA}�����B*��6.�V
B�p�����c݅�^�_���(q"h,�3�x��c��Ϸw �!ֺ���ѡl*]��*��@��Ƭ�v����l�W�!oX�}H&����/T�����p2�וsb�F���ʸ�	�-�yp�z����wׄ�ӳ?�"E�k��Ɗo���Iފ����Җ�7�.��� ��+�%�/���+��d�+5`��PK
    +Q�H�j8�  �  =  org/bridj/relocated/org/objectweb/asm/AnnotationVisitor.class  �      �      ���N�P���B�i 	tH�'�^�
Z�������J٢bE��F��V ��X�d�C!αR���R/|����L�><���F����z������ܶ#kA��Dgn�Q'G�g�"y���N�(� �dW��s����=���r��#P����CcH���=���Oݪך��V}h�Z�D�4����_�Q41���L��cLFe�HO�֭� �Q����Ư�'�Ә�ׄBr��z����?���[��*��(�"���nm芙�Ŝx�'��0T�o�q�?n�$n�	cY��&V�7ָ�_���/�D�k��"��.�b�w�;i���Y9fxծ�&.!� �P��ۢ}�I�z���y�J�f�,cN�W������M��d�#��Rt"E�b��\ʌ��d�/�t��\�ga-ɦ�s1V,��91~vIb	k����F�'PK
    +Q�H��S&H  Y  <  org/bridj/relocated/org/objectweb/asm/AnnotationWriter.class  Y      H      ���S[Eǿ��˅x�Rh���	ZZJ�Җ �5�����!	MB+�Z���Z�V���Ggtngt���� ��?���s &�����9��=����a@n�'�Q�P2�$#��P0	{x.14	�/F�<�Ԙ�X<�HӱD<���#IB�`����T,� e��
�u�F��S)�pi��/D_?}a�}9�Z&ӑ^���A���h��4�(8����7�k��?����U�Z!���*J`��ă*d���U�ƣGT< �G�*���*֣�G[���{�]#�A�h0����X<ڔ5sBw���)��N��y'H�n%�x���A����J�
'*m��@m��QP%P8>��'��JQ�)V�Nyl�F�@�R������`?��_����EC,��muV��8�F@�ӓ{(�td���ã�G:ͮ��eM��chؘ�e"1	��
�CƏE_�U��1��@颖w8����� C�sQɫ��6t����L��)xB���ᢆ_œ��p=9��39N��X��[#�P26N�!��Y���x
}6@%�2Т�4��
��ޯ`�{��!�}
��w(8�{ԑ��ŘѮ�f���cF��
ƙњ7#Ɍ��Q�
?_��.�~פj|��^!��#Eu������Q��\�e��<I�ը->1&ph����3���t�b�8�-�0���MEt�wr).�Qq��sk��L'�W*tk�E��SX�������[�o��P�E�.��W)&��79��Ul4X��Q]���*>4��GTh�5�@�-k,���33	��Zq�ڂ��6{�'3_1~I�ԛGPK�ꢐ6��YY�-���_[���V�י�z}�z�Q���Rz�����Yt�vWɦ;x�垅�U>�2W�,*\i[\vy۾�۱�е������o���Y�r͠,�R�*�s�5P���ub�tq��~B��V��:h�!�m�r��ܠᰆ#3��B��I�-7-�i�e�HӐ�ͺR?+Ud��B�L����p"[�	�\�B'5���DB�6�B!S(�a`�KI�ɠ���P;�KT��^�K�s�����Ku��$1}��(g3� �Yj+S*�e�B��~���)Hm5��&��2����J��j�Iٿ�r�(����gRj�Q�Q�%Jm5J�I�hYB��(�e��j�v�R�!��%�y�r��j�V��WCz	e�~�4\��K&�g��M��w/����J �#�{�t����T��\\ ���Mp�*���S���f��<�#,}<'���7�W�����i�5�n��%s�;r37`�t,ذ�f����A��p�ؖy��nW��7'~Wq��k=�/i�_�1���&�I�K�����j��*���a��=}�ϲo�k�gjM�i��c�G�fW�$e�4��ET8$��4\sH�����Q���J�q�]�	pȍ+�p��W��x|�������nh�? _K�k�,<<�\�G�EGss��.���u6j�|�Y?�T�uV�p+p_#�R��h,��+y[��9�Q�!ȍ�C�bWt�(.�Q�K��r��2{O�wu�7��PK
    +Q�H�}
�  I  5  org/bridj/relocated/org/objectweb/asm/Attribute.class  I            �TKSA�&v�!�QW��/��!	�A�
�*R���!�6�����.�*	�X9x��x{�(�*�=l�t�MOwO��� � 4�hfմ��l���/�떑i��c�*iU/m�3�e��ۖ��|�{]�녬����Ve�`��pb]"�B6�����,-t��%y*W�Y���Y��
��xq=p�Ӌ�n8�cp�J˅w�b��@�a�ʕŌq�O��a-�i#_b
�R猰�B�9MC�0|��/��K�W�c�qMK%����@����x����B�-G�7��X��,c���Q7M��^ܪ0�OW��'q�*M�6�xЏ�e3'J�o)�I�d�S���q�b+�/�T¡V}8��D��EBC�Pwk"��n��l��zD�����Hk�XM_���`��_�O���P��x��&����#1�ͶCm=���������E�b�S@/cZ��	�
"�
�3M�/�zF�'�DP���1�0'8��ыB=렁H�3�֐T���)^^��*�$=�=t�#5tn`ipⲍ�$�H:�����Y�Դ9�'οl�m���m��Q�ñ��{7b\��\5"U�^E@���{
�C@-aD(lN�o��=�c�"O��hsqP���MG�z�v�')��KS���!:?0�bdq��g��1|Ԇ��雤�q�ȇ�(2E\�d�O�H����w��B��kkE�1y�臟�PNٔ�T7I-,n|���O8b.bW�u<U\�ZG"��b�l�� �����A�d�PK
    +Q�H>O��o  �  6  org/bridj/relocated/org/objectweb/asm/ByteVector.class  �      o      ��Ko�@�����`Z04ԡ�g�P"D郂�RUph��z��Fi�� c@E�9 n�7@�\A�%T!N�K�IZfm�n��@ٻ3;��of'���? ���35�����W�v�R[���b��j�+��ai>kݻ��\uJ�d�l�A[�XيU-go�q2��b��M�d��<�ty���1D�C�*b��!`�
R�f���Y��}���p���5�B��%�p��8��1���n�Y���@�|���k�2G��J�+�*\��p==VpƱ��呮$�v)b���egɭ{^� �q����d�W��WU�1�r�A���m[��s�]�n+��=�tG�C�����$nn��럑|W�7M��01L�Wk�%��
Խ����/:{z��-F�,YI�`4�6�B5��u�3z>��<���0.��a�ۢ4$��s��8i~��QC(���c�)|���a���i|�^��K�~_`�^i<��Rb( ������G��71H-�1p&�BKm��vc�ҔǍ�pG69`�&-�6�I���#�+�g_�9�sNy�r�,�q���Nw�gt��=������6����h���ȉ�.�����P���@7/m/G?���2�h|���#��N0Z�qS4�mo+t4'��]�����I�$��]Ҟ���H�B�����Vt�x�]	�5/>V�Y�t)!o�q+ڄT�#u�57�$��> 7��.Sv4iVL
��KV$;@�}�m������{��R��H�}���v��'=���}���t��Ӌ��fUiR�"kn�o?��H��4Jg�[�,O36l����B"cp������nT(��>��8�����,�'�_3Rk��&�Ժr��'��|�+&��� PK
    +Q�H�N��   K  7  org/bridj/relocated/org/objectweb/asm/ClassReader.class  K      �       �<xTՕ�y�d�s�d� �0�$�� 	 %��:C2@0Lb2Q�m;V����-b�:��-�dB�v[����j������nw�m����s�{3�8h����޼w�=��s�=���v��g �FY�`Ao��ڝ��]{k�#=���X���`�;�F:c7Fvֆ�ծ�	l���"�N`�{�7�k{��ݵ�l��W�l�vՆ��X��@T� �n^�e-A9�fS���v�r����Զ:�B;(;V�C�Z�Aю��������z��b��#ć��hwl9{厕�2p⽥e�VJ`���*e��*�i��n왆��G>�{z�c�ʖy�̀r"��`fz𖞞��pOS���}�h�yg�/��u�lT@��%:н;��آ�\�$��4�B\5F�rbN�֠���V�bp���|Z���Ě:;#bJ�$!b����"�+�eS���@c0��eǪ,X,� IY/���E�%W����5K4X.qИr�%���
�@x弬�eT�N���w#�zZG���Zb�}NX-u-y��a-�`e�[���x���\��D�Ǚj�*�q=��A60�OS����o��A^w4��;6��W��lk4h���[�F����\e긵7�["_��v�A��� WH�k��1���wpgO�	�5�$��J��\�A'ty`'�j�j7���`je����{I��L�V�E4�'u�\4���>t�&u4	r+�{�Q�~p���ڌ\�I� �S=jDh���*+'b7-�� ��&��^��|�n��104�n#��Q0s� ���՜nG������?|��"/e�;=�A�NͩzRZ��#�Q��]�����lvipi�z���x��yeool ��[����p��c��\?��u|Z���]�Oj���z��,AϤ��!���a4�=�=�z��ȏ�A��ۭ.\���b.�QZ�@�o� !E�GR�Zr$ɾ���%��F�����HV��ؐ�7�1�,;��y;V�h�!�>K!m
=}nܬSъA�x���]���Nx`����ԈZ�*����I��P�ιH�l �poɱ��)8M�=�j:��\�4�5�+�4x�p"i&�I[{e��e:%�h0�"��������..�8jp�y�+�/��3����z�].�)��x���<iz'|-��=a��|�L�[�<�P��T����x���;6��8�_�y]goz�?�ٶd	{���߇�v���?�
�[�*��)�V'�y�d����nr���ډ6�P�;c�o~�`�%�7ш�K��W�����SŚ~���%��1"hq���n����8d�p�P���Y86؏T�C+�4�uX��MQ��09&��=�:������6�ŁhlO$�������EX��fud��������Q��A�9BK�,c������"K����2QF�ᝑ��������$��Ǽ)Ԩ<x���n�&�d�ݰ����0_ZU��:E�bv��0�9q�"����`�R>qp3q�A�6����j{鄸d���o��7m?����l��YN��VH�1h�\���YQD�2���J���[��`�D�F�|HS�N�]f�"��T�_��)��2�#Ƹ��B8������b�5ݑ��^�v"K�2A���k4��"YgO؋2�l���eE�jt��5G�4�Ǥ�@ܓ�T��X5�<U��X-nn��:�+<�s��AE7��qÈ֟�n\g����1/��P�m�T�gs�	*]����b����t�Z��-�-��Kخh�ǖ�Y[����I�7({#k��ѱ
n,��}l5k�a���B{�j����]�5.�Z�խ�6��]��KP���θd\$3��A}廉^�l��mb��~E�,����6
g�K_|�l�l���`U$d�HbYLv�Aw����	��$����s����^��$��D�iU�����;(�dpM�ߨȐ����B7��d��_.���`U8ֹg%2A�C� ���9k��Ǣ��^r7dг5��M[����b���Ѝv1�\%c1�YX���Z�����};#�&�F:�����m��;�[�3;oƐn�\���1d��[ѽ���Ф�u3��?U�/��{P�� k���o��Dp��������lnijm�޼����Z�q_��@tR�[��;ه���a�8u�	�7��s�4�Qvn��ݸ�ki�ܼ�y��>.���tM놦��OB�G��mk5���	d�zÖ���� :��9 ��v�t�%?�>E�
���O������G����2)mCX�cЙ,����ߣ�R�_��0ˮ5���#�'���u�����&ib"(�x��Z�Q�}��P�q[(��[��I8J�G�W��=#r�I���;�){NJ�/�.O"r���1�mF&#�$���;�N�O1�rE{{��+��D��;�O�gH�g-��7I���З��֮N)T��9�t��#��v�B���-��u�ve��}�ɾo��ML�u�hWO�ɾm�Xy�^Y} ��mʸgb���X�{��Ѳ1
�R��l� �|��+�|���,����"7�3\��"����:&�0��wL�\*�~��LR��r����{E���駊*�	�"5;ٯx�ř�ꎀ�{��%N�5��_����o��3�Y�D�.����d��0ؐm���6�w�?IO���㴳?Rq�_��~:�w����R�Vc��ٟq+�����	G��ʏM���c��ُr��λ�_��yӖfMa�(cޠ���NE�Q�Ũ�ã��uH+�1m�;is��	s����(E�l�9:�OS��e���)-�V��7.}o(�])P
q��䯝�)ѻ9�Q8M��J��+���bY�Q�*:����5�L�0�ܶ��US�K��eX���9�'�7;�zq{/uLM�:���+�j�Dw����u��>�Y�E�|Y����G�*�Vs*�Rk��_���1J�J���ƣ�)�i�v*�˗���i�4e�\�%�Gf��=�D�9�ye��*
��� �fз�Ķ+�M���v���v.Ї�\H��Ž�Ľ� a\ܧ��<HY�-��+4���Vuf.������J��(n���?
>�L�{I��]xrNAE�(�y��/�BI���@�g��է�f��{��2���N��c���5���;>&_��)�&�������sܺ,��3q\�+�n�w��q�iH�3d���ۏBw�hN�t8��.��/l�s��!�,�Ts9)�)B\����3Q��6�R P�!��;mOB�quY
u���I7�I��4�>�_jQ7Z�M�Ҥ�B��r"�:B�R$^V�+�Vv*%iPŵ���a�gJ5��Ku�i��q����|mh��lC[������z���}OAsPU��o��U����p��t�p�B�y
�;�}�]�)֗=����4�w�� ^���	�mףi8���Wh�;�BO�[Ǒ��	��o�x���!	W&X����$�%ac�ͶZ'ak:�(M�(��#J���{uB�*��8	���-`/�8�.��=�"S)�?0
=;���P(�x���*'�MOzn�bA݋L<�"l�:�� �_��8���hh<��(	7' s�B(�u��>E�U����]w	�9�{�F�2�8n\����ۻ���m(��]U��q��#p_�o����7f�9������5T�zQN�ES��B"��a��
�&�4��SU��à�4�6"�;.$.�����o���v5*)�W�'tg�o�y�i"!�c3U�è!\;�A⇓0l�Xlh���\;�*�A��4����x��P�W�W9ȫ��<��j����s
?}0	��y�^\�|=/��i����\�w���\��#�O�����]�ǂ9z�X8����������L0�6H�tvx��vJ@��&��p|�8����C�'��M�:\g�?#�8�U�om���3���O��$|U���C�)���"'އ�� �<�Q��Qx�i4��v��-�|�3>���Ȝ�#P��a(��v��n��Nu��@�^:N$|Y��q5�1��{%�g���@Б�q�)��B>��|���q�=�u��ąۃ���i�P�S
rm�[����>VO����`>a��"���)x�,	�Y�#�@*�0*�J����f�����'��/���ɾ<��u�<��2���i2��5j����^iØ>�y6#?�v�/��y�EMϋ(�]{ܭĽh[��ԃ8k5�d
|�t���u�[E�mh8��k
�
��L�)�k.^L��Cj�Cj�b�^�9����ʂ:^Ƃ�cy��)m���^&|�H�#�%	����͞\�a�'���ߚ�Ui��Tj���q����૑�t�i7�_�`Z�f�'��;�#/�W
�)���O�V�z�O�,��	+��c�$���Ɣ������:vgn�('ak�'"O�TLϘf3�y1�C�^��6�i����(�XnL������j@/\,9t��F�Bp�>�,���u�S��X@�_K\��WW�1�a6�ѹ���%������>�,�T�%��$���g!�J����eI�Uɒ�-�{0�%���C�T5ӊ���U��U�5p�e�IV<ʦ���]aX�t�Y�a�d
N��P�*ݕd�4�ą_��!���|ig��vCU���|a0x:��\Ѵ:�c;��0�I�H�M�组@����E'%�>��pЈ�B�|�a3|��b�Ԉ[�շM�G�(b�5��|	�D�ݺ3���,6ڝ�F�dط۴�{t��(M�-L��&�&r[&����JX��s_J�>��$�Nӧ���d��V^<�Z���RN�R~�1�E��2�ⴹTJs)ǁ_�?N�2m�����^�I{��>-��؛�.����;�gj1m�3m�,\U��aH��2Wzm-U��nG�1U������\�o�=�O����{S�pՏfY���V�hqyo-��<���}Y�#e��k���-ʀ�L�QČȬn�����oc|�i������g'(��9p6z�m�l� g�b�S۱KĴWS֤�N�`�B�8˶�ϲ�!�K�x�5��sN�'�*��p"bk��g3��ρh�;deʹ	X��	��S	���g���S���F��0������!�����on��ayk��!��W$���ͺ��sFY�6}�Y��s��YM>���23z�S��&�/M�������L>?���La3QMD4�B|���"�M@��E�E�r����7��^o:�39������[I��f���~�o����b��r+Ր^�d{�a��݌�y]X8�\[X �'Yȓ	����)[�W���v�ym�\��`^X��ͯ�uW\c	fC�����eJ�l	�Mޖ��q�Iҩ!S>(��\m��d\C�?I�����]Ta��X�����P��<�QT?0ى�z��9JU[5�B��#�K��9����ib2��||\½�/�:�[+��~��ٮIW!������j��%Y_J��,�je��]�T��Qm3jlF�͘o3،:���f,�������Uc�Ȅ�r�����"�oƛ��`C�Z
�E+��Q>������z_Zw0�,s�8�b�m#,ƗZ�?�6X�|����Ɩi�	VR����ɑU��;�":,qF�M�|U���"�w� �>��CpT��IU���!�'��"v�į���÷K�Ɇ��Ӟm]��ם`�3,��\����6�d��5���16�f��_�k���|�S�>�n�y��o3�܃��C0��ݮ��*G7x0dO���'0�ʖy�'S��F�>�cJH��ɃMV�?+�ځ�~�6��w�L���翤��/�{�>8����ą�T�l�S�Ob�=�z[�$9���A�����-H����Y�p
A2��rP����o�-�2D��N�����Q�k����׆�]ð^�B��,��bմ�������aL*���eD,�SG �T�yh�$�G�Fx�bE�*�_���0�C0�>M��)z���0���#�g�y��9�:�{�/X4�z���.�'��	��S�����?��%�b�&^�d��J�z���"^�m/�7�.O�f^_ ��L��2��b� �W���5Nc�JhXh֐V�5
Q�~J�����O��,��1�vc>��.`!_�Ea�.�Q��(�E\ƭVM~��M�V-�a(��iA3���U�X`"�1B��1�J�;���"c�OL�]��2bfQ\>}qvt\�}�E�i���1�'��Mg�z�����mOg��- J^sѯ���N����7/���O��y|n��*�'�.��N���h�I�9J��[p)����뿢Wx^o�)����DJ���D(τ
��Ă�6U)�%�(%R[����]�mf�=a�ˬ�i�Z�Fu�L�f*��d_�By��Y�bt5�|5#��ҿ�4��Re�	��x�Tc-���r��>}9>U����Ey���3��/yF_�dgʶwQ�=����i���q��
*ˉb�ޘR�#4�K�"��p������B�im��+	��x�}E�N�ZR��B�>�Z͠77�_w`���Ow QT�i���7ɣ�����>��1�J ��jZ��0	W���I��x3��"�/�+�7E����a�R�*'6�������f1�g���5���Z�����J�-����s&Ar��������=�R���I�
����%�w���S:
I�ɗ!f��U2Յ�z�s�0l����Z����o��1��ߓ�L�!x��y�l��jֱ#[�]TJhk��.��1�a�s�f�N]ı^�ZX�%.|��2g�f���Yt�x�e)�r\�ן�����z��z=o��G����P_~����yz��6}��ą��6ĺ�xDS��u�×��8��Ϭ�睷[|��$7�"n�^�3��݄1����9����c`�7��:�.�33�9'ٿ��.:�����a\4;w���N�A��&�n��]h/sz�C�x�ix�T��0���������_jU��w�q��G�ói�)�6p�פWJ�vd���V��������KWqC� ^z�����2���U�Go�� �� ��w��9]=�BB�#^=^t�߈W�Y��+�Wy�+t�_�T�S�G5��G�O�V�^�� f�g���v�?1���z�l_�b�o�����;�?n��y籲�ߪ��ӣ
�x�߸J	�M=�^��9ы�@�=��/�U�.����T��g�TlV�Q����7��,����øwT�51���H�R,ȏSaFԣx�S�R='�b�	����(S�x��i���Cdx����J���qF@����]��B�@�T	g?�w��G��]�����,�ӫ/����N.�>:nI6ǙM|?�2ʭ;Ĝ/$��T��G�t�x�<��:9Jq�>qpYnD�;cp�x�m3��"m@R{ГA�Oz�1���!�'��"���'�`Q��(sLJ8��9A-�RGy��1��EyR:��)ʙz��1O���X�?!�\�x#;�]�8o��'aצ1�y1Z�#��2�13�~C�S�}Ek�W�f��i��2�p�����>Rh��f��V�=�L���v|��*��p�
������p�
!��C5Ah>����3�_�)	(ƶ�'�,��`>)�J�a�>�|�Z(�;���SlWǨ2��ǭ�&����DΪ<����8" �8��>�bNr��$���{��Վ��2���¨C(�S���I�w�����xH��J��E���N�/����蛋:��})�)&}N:YHsSHsL}\FH����(5��,�Pn��5iJ/Js�EԚ��$Z4�hj����[ â��q"l�|)��Cn��}d�m�7�KE�{�2�����%���0ɖC�$[�D�y`���Xj��.�R:w��qR���A�)B�$$>�I��^��7���_*-�/T�-��z��*�����"Vn�(���Z�R��𺅻����[~o5w����ݒ��tt�?}
��;�ཆK����ʧ�]�3	]^�~�Xq�{�ب�8$I/�OAMG��;F�*�s��)=���������O����g����J#].B��%��Ŏ�f�6��FC/^���!�b��O)���m�J��S�I60�*�R�D��Qev��l��q��w���4'�^�`��]��}�V�a~;t���7S&�����o�S���y���ꨲ��l�PK
    +Q�Hb�'~  �  8  org/bridj/relocated/org/objectweb/asm/ClassVisitor.class  �      ~      �U]O�`~ޭ�`+�P�Ɨ�tcPETp��M�L� �B�����ٚ���a"%��K/�Q�s޶�.�v����s������? laO`�����g�Nt��]ӷz:߹����:�9��������ؾ�� fN�3S�α~ �9���G[@���N���[�g�c��ͨ	�j�8D�#�(䑂JҴ�<��������fVE�TȜ����0ڣ}�v�[In�]����2n
d�C���Z�ZRf��3T����Է<���^"��y�ļ�1��q}ӷ]��p��m=a+FDq?T��6�#0�C�ШhIyc)�.�1�z,�p�aY��Y���h0�@^���~O�6�`��ݗV�B�ȣnb����(����.)�2���F6��0�H�l���R�K����\
�i��ݞ���A���ʼ����
�-@Ђ��{�N%�	�Uq����
�J��d��K�4��k4/P���sp��sd�P���jm��T2�l��؃v,�X$b��=T6� �JkA�H>�3B�B�f��KSa�#����Z��sq�i�#p����gBpA�h1-Mh�\�:fȖCd1�0�h�h�a5���Q5��jSV#���jf���uz�����y6��b�PK
    +Q�H��߹S  76  7  org/bridj/relocated/org/objectweb/asm/ClassWriter.class  76      S      �;	xT����'/0$0$�"Kx�!0$�����!	$3q2A��Ƶ�]k\A��ֶA�+�Xm���v�u��U���j�^�s����3��������{�{ι�{_���# 0O�"�GZ�6Eښ�E���@4�\İ�-���e�ME������@W׺H[4�",� ����-&<�Z�����V]RS���&�草ëה�T�1T�� ����5We�sM0���M���5Qk&�ӤP�#��� D�mL�v0�fj-��Z��Q�B�<j�Rc-m�֎��jK`[��=j)��F�B-��A-D-L�������"Ժ�E�u#,IS��P(D��!io汍�e�,针�t���A��Nm�˩�Q+Oߔ�m����*�L�&m'�WQ[I���
j���m���2s�n�	� *��R'��Qa,X� I}F��c��T0���U9��Up�8�G���w�P!rs����@��0^
w�V2m7L��:&�х*L��u*x�h�
K�,mT�D�>���`g��$�s2�!�t��3�jؑ�&'l�f����[��f��Q����?����x2����jޢ�9��h/B!�R��UA��ө�i-���򈤴��V/Qa�\w�
��*L��ϫ0C�����0�GW"d��օ�#M����z#�$�/���(sG�N%}�QR�����kU�-}�z��B��"���JK���ϑ��@ʫt���L_d���V��*HZ��eL�<v�����I����(��I�u���}E��h�+p7k�����b��E�o4�!sy3���0y��T��g5��P(a��T�&�����+����|L����m�5B��ux4�C�Ph��KF��BE� ��0O��cN�B�C�+F� ����>�s¥��I��:>
��۫�'�0 ߎGQY" \5Z��J�'	��YR'W56xa�P�)��� ����Q
wB�U!�jV4̇�,	��k.���t��m���M�N�U6�.%T!��m��i�pxZ{ ��n�c�ȵ��N�UX �ļ$J/?���De��m�W�#�]���OD�g*,�b��s�+� ��Feo~�8�̯U�/O����T�����hW4�(]vx�Q��
D�#A;��"�, �IMv�/���2����j{4�"���w��BM��.R�$g�wM��Fe�3���8ݹ���ώP�5mk��Ӆ-ׂ$�8D��=��x;�ڃ�|Ck>F�3���m)��I����=��X����m��t�ʙ�Ӌt��z�r�?U�2c���e�^ig*M&��&5�|��
QG��J:ഞ9QǢ��m�MhS���I*FBǨ�3Zi�I�8F���� ]TU���	���1�4h�����D���s�C7N`jUx���=�F������`�Ģ����ڻ�*�F� ��TJ��Wb�:�g:�:�
�V�g:q�MLT�"�&�8��T}
D`�Pq.jN,�B:�I!��D��8��%�"B{0���ƛ�G�^��p���#�U��D��N�f&0�U\�g9q1��.�3�E)�b�]�
�ZlH�AG;��V�t�/w�r���ȘW󪦸��Ub�G��f1N�T�v�҉~��Tf̯����O&^p��f��c��Y�M��o:6���[K�n~����ٕ���l�U��"m�t�(�=YB7�E��9ޡ`	�
��Q���|�R1 WmRa�\Eiܛ���B�l��s�l�V�=O��~K�v~#�kG[vel�N�˥3�bD{{�%�^i�����*��&�Ȳ�{�f>��N���m�p����etv����Ԥ�$���^q�p��7�;�J
nѰ�S�*6�6���(�h�QP���P7ũs�<V˵X�O�%����78�̗�M�8[��,�M��ï���\��"�Q�nEf��徃CE��c�.�+��5�J�H�����1&{�M�k���ߨ�M�*ޏ����p�$��ˠ�(R���������L򫒤����#ܞ�<�Ħח����@WkE������[�Q���o�H����x�]����MWщ�EW|+q��'���<Q�/��p�%��ħ�E��-HK'�QFz�G��ϑtd���[��;B���&�����E���A�����s���f�"���v�_b�?�����#��VK{��?e�
	x�?����'�H�]�����Q�&^)������ɶ��u�5�=�f��7yǿ�zADf��NH�H�������q�:��|���
�ů��ȚkG���t	u����k��"��S��M���?�?���J.�<ᎎp���s��nI��IQW�	?�}��+~�ǿ��$�����%��e� ��8^|6���6�n�c�����3
��O�"��VE19T��a�`g{�.�PPQ�j�U��Y;-��p1��4�S�)إ،�T�X Չ���d۶���.~Šz�:��Z�$4��(c#��꾭K��IzUɥ[��۱_ֽM��*Iu49IVɢ�U&SMD����{��2�ΐr;9'ieٯ������ղ��+V��T�_U�����uAF���+N��\}��8W���.�.+����+V�<a�
�r:|k-��G+Te�2�]d�U��Euů�fN�0�&� P@��V@E����F���oL���lя���+z�\*�s W���&�~��O2z��É�AF�S�¿ĉy+L���t��a���L��2�g9�	J�F?�^
��>��3���0��7��Bџi�X�E��?ъ�D���1�_/��RXJ,��kH�
��k9�`�f�A�v*7��1�ktv���1���C�vj�\���\@kVҚ51X��'���-ϼ�l�>0�bp��gI������e�Đ)�$�������P�!�ƠE���f�����S�Cˋ�V-?�����ti�t{̃��i��c�I���L}ࠑXv��:���X�.;5��Χ�1�e*��m��x��E�۶�0W�ذo��HW�nC$���O/U�
�� �������G��h��ǳ��4�&B�;�Үn��q�;�.k=�	���>�T�{L����6hf��2 ���{��1�^���aRK��A���C�{����B��e2ل�dL!-=�o�Eĥ�&|�X�ͳ4�i��c0&�K���qsc�Bi��*�@o�M��@�ܖ ��<��?�a߱��}6hy^��졭?��ax�X9����t��$�Q�x ��c|��l���.�</��[�N�/&��qW���0�!�{��g\������R�R���L:�G�<�ЏK}���0P�7t�T̖�E��c��3汛����c9�9
GJ,}C���A��c�<��?�덍�ZΛ�#V�����k9o��$���A�0� �1yS���g�:r~�3�j9����\@��4ܚ��N���䵼zY�����e?��#cvo��^�(f?1f�'���~j���ܬ�:�����;��IQt�[c)��_)�e� ������C��Xr��y�ė�w��&EG�\��r-o�Ulk;�ve�N��%�+�9�$�י�n��#t��1�'zD������1���hO�Ň�t��oL�Xx�#�/��2������8	w�����(��YIP��׌=J���oIl�����c���=�,9T��L��b/|G.t;��{�зdGn6�׽'�ن��$�y�AZ�^./}8�}��}sSz�@�p$�AC?%��`B?�xT��`B?䠓��D@���P�{��Os��s�����c��za�aP6P�j,q�M<6b9��=Z2�Cj��/`2$?�ɸ���8\R�,N�q�Gq��Ӗj�:��O�Y8K��	`���M �I�<�����!�|�Svbr��X���U�L�1p�.ױ�\����K�_ǚ�\�g��^J�]3����^XL��j�:6[��c����ul�o������D�Q[za
���h�C�Fm+�ja#��1��0n�0�����P��.�8�=��Hί*F�w��A�	�;��?j�m6��!�s��&[�5"�x#k��Ja^�fo��v�:��8��7p�+���$I�n�0}6j]
��.[�A��`3p�d��{S��O��7��?b��I"�=��S���H�/��Z�4�\A�=��N������ڐ����@x���������=�pL��I�ձ�&O����Yb���d�X��>�I��5M��ȥ����Q�Y���C�.�R�q��!&AC��>�Ql�b�G�Jm+��p�o��c>B������!��1�J�n�ǩ�c��$���6����\��,�(V#
ٚ#�J�<Y��ޓuu��=�ͣ'ܶ��ɒ���7yt�X5g���Nf�p[�ٍ�W�O^�XO63�S���Uڀ5���F��,�6f��~�:�O�D�B�3�'�TO�/��U��6^�6�5�(��r�*�(�m �?ـ�ـY��'K�*�.�d�Bi����eȀ���I���p7!��c>4�CT�� ?�4f*�Ysܝ��6�2?K�?B���E-$����ns/�]Y}@ᯘ���n�	�Y=V��mIK2+�aX2k\�}�?�������m��l��s,����'?+�<N��6�%�Yi��z��?K���)����0r���+�Ն�+x�T�_�;&�����į%�C�$k�`�#��Z�x�A|����d��"^Z��#}
�Л2.�O�홥���������ӆo�0��ƚ:���y��A-�&� �R� |�۞���vG(r�prXHN�B�a��N;9�����5#��kK�'L��΃��0��rO��5���{���;c�D���9���9(�6mp�"�CǶ����cx\Z��pB|��\.~F������a�V����g�'�c�'���޺$O��`7���6a�ir��yW�_횶������iyIۋ[h��[pߥ@E�|1��RϏ%t�Ŀ��7Ro�4�`t��B��hm�sY���nM�!]����\�t�a�=�d���#>-}�Sb��Ǫ+c��,�*9�`)�ˍY���<r�Y<�4W� `�e�c�湊�C?9�f�\��0�s�hK�ϙ�����k�ti$O�	��,r}e*�$Г5}Co{�0�貏���ny|�x#.�!Ari���ܸl
Y�Ĝon�b�^(iز��� �<V��R}'%r+gR��J)޶ �Or��y�%־��{,C}CG��L�6���P+��;Xʏ25��)�u���א8���c9@�Q	��
o�T��I�ʌ��E���9w���}e�2s�ii�v�!���	��U�|�������Ǖ���PK
    +Q�H$f�   $  0  org/bridj/relocated/org/objectweb/asm/Edge.class  $      �       �NK
�P�؟֪�.��� �q!ܹ��QZj��\	.<��Ӟ��d�a&��}����N��3���U"�E�U*7Is7J��Etj<!��M�B��8u�$��P�U���X*Sl8��f�78�n�2kvk�8"�acD���6���+`1�h�C��|����)s�8��Gg�PK
    +Q�H��j}  �  8  org/bridj/relocated/org/objectweb/asm/FieldVisitor.class  �      }      ��MO�@�߁"_EP����jlb<�`L�ф������b+Y��)+�-L=��������}��y������{�#?h[�@8+p���-]�R��Vǽ�/n˲{�֕p�NS��$�P��}���^ۺ	�$ℸ�$T'�������k��S�	yFЌz�I81���6u��� �[3&�b�:XH�Β�$RjU$������Җ���Fcf�V�k��sv3���c���5�⤘d�ֳtyZƼ��3��l*�2!*^z��-�3�m����'��J�9�4�c�S��{��"�� I�Lc�^�d#���q�ys��Yb�<�4�^�0������'r*�WFX� ������*[����2�e;���~��C2��;?PK
    +Q�H���    7  org/bridj/relocated/org/objectweb/asm/FieldWriter.class        �      �V�SU��$$!] M�>��UCV��b��G��"���Zِ�n6 ~��t�|c���҇:C��g���X���$�t&If�sϹ����w����� 0�}�����Șzv+aj�ji��
�-m���2	��O��Z.�d�f �M����n��+ 2�����bщ9N�k�ZYZ�uZ�6��8mK��Qw��ڢ:4�²L=S�4��O�nM
|k!%e~K�Q9��H,�Scc�I�m���@� ��)i	t�H�B��=�*���3�7��`�K�Ao;��#�.8�����+͸t��|��W������g�u	�{C `h�w�̍	t��_�E� �!B!Khw�%�.!�ÍbU`*vJy��XZ����
��*o�.��ؒ���m	��F�k��P�[��S�\ic�Q��Í���YZ��|���ƜQ�a
4/�풵�Y0-��4��;����-v6'p����{��rW��ۼ�{9�A�:��M���M�������N㫯ݞF�P/����@�I� �x&��,S�m@����{z�;fF�R+��JZ�����<{&о�gX������
z�B7�mS����}�P��I�5��J���5�LN�w���p>��}!��T��S���[��{3���1�B����in���"��@P�t5ÒPr|�ݛ��W��a��#Ͱ����l!�a��Bz#����զ�.���o�M%��۴˥4kD�������j<r�/ʇ��g�x�������R\.�r���X\���2��r�gs�Ѷctж��&��c�i���!��1��'p�n����h�	���0�0?�e�T���(�,��a���� �Q���(����[��JRQ�c7�"z(}�ot�t4]�
'��b��i�\�������"���i88AN&(A��O��� mbg��?� ��Q��#�RYH9�_5Xs��8[���ɪl��{�=�l�e�a[VAnu�Ѥ�Z��Mմ�ct�2�#���T���D�Z������r�*?E�.��T�\�X���}j
�C�y'�Z�xE��W��1;ow��q��˥ja��gZ��:)�sP'��V�4z��qO�P���[�uÙ�ݥ2W��o]�s�?1�nLJ *׺T�H�99�J��L�JJ�����[w�PK
    +Q�HܡS�  �  1  org/bridj/relocated/org/objectweb/asm/Frame.class  �      �      �[pS�q��z!�}�&]%I��/�`��N��6� Icْm�-����Ih�-i���PK��	P�M��Ҵ��L�3�Gf:ӏN2�f������WF�@#��ݳgwϞ=���K��M@)�I,�U���v���=��`"*#^�}g�#�'�^��-��{��$���,�	F�ʚ��d	����H�KP��ڌn��{֠NB!�ЉЅ@��"��F��D�ra��s�%P
�=0�.��M�g%�Z��X�E�3�n&��-��*��s�nɘU���D�����xpoG�o�F��3_Ә��H..���p�a�������*��D��yx�PB��H)�ѧH�����`��x$����ޚ�G�]k(h_��F��
7��[D}�� &
(����a��|�wt��	3x5��*7���%pD���`s��A#�:2$�ǆz=�hW���	�_$�ױ���ۗ�&Z�+���p�o��>rm�u���h�ك�o�a���.�̣��>Y��Ȫ�Kb\�'���a�n�`IW8Q��G���PK81��F���=� ��"���<�\39��1��q��M�.�����t�S_b
H#4i	��d�5�Ո��vz���Deș����4��.U ��~� 9?�=2쟚��l� |Cq��	њaԶȸ�a0���Ն�;⑾D,.��¬�:�iG$a2�H�^G��9\R��x��93>q�Nx�Iu��G��c��eÉ�X�f鄧$��!�>���3P��m�C��:HT>Q?���̒+-�D�7\7��KDbQ�D�������m.���X����/�9�$�:b�}�0?��b\�	/����/��T<E����i�����T%�w����m+W�?cTx�
�9�
?�
?�
?�
?�6/���#�GAS������m7��c���G����\� �4�ɯ�R8-Aq���j��8!�33�<�.%�I8'���1tC��u\60z�)za
�7V����o��oe�0��/��U:�7��N��8�v�Kƥ�z�kh�����7�_]�_-�ѯ��	���?���pku\r��T��SSW_W_�����>��Ef�����
I��	��y��x���Ba(��6��-�>�^E8v���cݬ8����s���\��aV��S��#V�	Xt���QY��
�λR�4��x��'���-�����-�ԏ@'����RO���;�VW��E�g�/�����\��w�z�6��}n��P�/�+��,|��W��Wo�v/)��>4L��D��BjNV����:a@7h�N�D��|�6���v���fd��rRk��e��u�|g`�L��?J�J-�����|�a�ᛀ�>���|l�(�V��Sb���e�J)�ĵ�F��8ܓ[8
��E�P��%�V�ב}���a�u�v�/�{>,�����l�m�����M��[�b�S~]i�C���M��(�֑r�_S��8������d�N�e���f ���Dx�Ҟ��J_?�P����O��m!t7�Jh�%���2�*B��Մtt8�����\}PSGf�A��J\9�?e�QX�N$%��4���AN9�'�F\�^�F�5TBF��!�[���@�H�S�!d�2��d�6a�K���.�E�:�3�g�;�>%4�K��{/f��[;���r��PO�s���&
k#��~܆Ju�N-^W!QW�̺j���Ʉx]���3^��0o#M��k:�DY��"��$�l�0�5
� 3�����!Q��T�"dT=%����<DCjJ).���vD�������ٱ���.m�e�;�żc�`����[��QP})�ѣb_���t��p���)�AC&4$�n�s��������T�2��$�7��YFg�%�c��_�ٗ��#��i�ь��n�F�ۉE����]�@�d�E�t$��8���Q�o�ߐv#����y^H\ċM�r�5W�Z�xP���.�.AZG�)w��}]��@�F��a��M�s��_�j �j�B=B����,»��;l!BB/�n��W��6_O��Ss�,�C�?#��߂Ќ�C}�O�>�x��B�פ	x�A�Ձۻ̈́+�,���V!`�90ގ�Y����w6�s!]��34oO�-o'�W��I���j9�$H��{R�g�:N|�`�-��|�4��<��U�eǆ�6!t#`��Bf.xiz��c+����2�V�i����:��W�~2�����N��y��t�M��'�9N��p@yV��^
���NѲ����9x��Q@5؀��q�݂���ҏ*��N'�s�3�;�����M�%�y��=�*�)q���u�_Y�0-�@Wӏ�����Ӧ�73M�d������C%���*��Ҡ+�oRnL�ڧ�����:��W/ʴ6ӕ!f�"�M���m粨�י��C}h�i&mm�̱���ed��ʚ9�r!a���C���4t�y()]6���+�K�M�SѲؔ><�tN�j�R��m�	8��QB�����^0},)=e�[z��{)[�Rg��̓���3Hؘ����8����G��5��B�}�̕
��`�x3���7y��e>��7�����@؊І����`I����~Ɖ�9'�1�	N�0�[�8n�'^6�/8q�`����܏
>�%����F�y8�mN���3��q8;��}h5؅�[�d71���
KiO�(0ڒD�(1s���y˱m�G�|������D���t���57xk�N;�����:�O�g4���#�5Gi��9��K�\I�Ӝt�t#�+�<m��}�I}���/�n��4/��ar�4;��5Ӆ��Ç�6�enD.ڈ�
��ǣ�->����x����*�g����r��W�J�Qؔ���i��ҟ"g�"�/��!���~1eSJSR<d�=���5O�Cz�`����p��I���X�����]���2"����Gs�Y����r�?�Ľ�s�Ϙϊ}�$/>䔗}0��3DS!�=�VS�����mVR���0k:�@��^!��g�v��]Bj|^bM#��=����F��� >N�E�u��&�0��r�y��8[DE�O�̒ux�eJPX�����Y��TtX6g��0Z!�#tg\�ྏ]� W���"C���ȭ5�a�>7ށODQ�PK
    +Q�H3�%�B  :  2  org/bridj/relocated/org/objectweb/asm/Handle.class  :      B      �RMoQ=p��"�j�����~T-�E�B�jM4M4.|�+�C���-�r��M41��G[�H��{�o~���@k�N�nW��Z��v��]Q�e�Si��{ *6����Sk�Ao�7�ns�noyA���T�)O�nө��ҩ1��5��{�a�(���O��f涆38��)!��@נ""�����Mk���u���{h��[��2L椱Ub<����]#,^��v�!el_F�|�ϊ�B*�5\ĥ.�
�m�^c�S��ɫ�t;>�a�~}gGtU1���	�ޞph�c�~N�|yICYa�!kl�ʳ%�C`ވ��O�ߔ�[����mE^+�w�>6�|$�t�D���l̳0zP���R�#]��u�sVv��U i-��2� �ϐ?��Ȍ4q��l���x�";N~�&©1<7N�az�����}��> ���?x�P�����#9P��{����&�Xx�ً���di��^�*���X<��I}� s���U�Y^�\��Ĺƫ�l�h�uP�V��|~�W��Л��E_]L������I�w��PK
    +Q�H���  �  3  org/bridj/relocated/org/objectweb/asm/Handler.class  �      �      �R�n�P=7�}��@����6qR�cѢn����	����D��Dr�vS�o�CʶH�Z��H|TәK�z1sΝǙ��n~x����0�aҍzA��m=���cð�GGq���D�8��=}���t���H"/ 4�����a�ߡ���M	TZ�e�����1�'���g�R��;�v��wO0_����M-�V��2�3n����36���=g�p�@#�p��E��k�ț���t��eΚ؊�"J��\�qGևac��O�m<X�`a��m�z��sd�U P#V&��_��k�N7��R ��'�Ņ�_B5��x�B�.Q�%\$|g5���	
��1d�����u�c�T�q������̱֗1��L፱�/�H�8��[�����-=���9�2d5Ū!�)��L�i���X��$�s�PK
    +Q�Hj��/3  W  0  org/bridj/relocated/org/objectweb/asm/Item.class  W      3      �RMOQ=�Z� mK)X*��c�Q����qJk)�6B���L�&��1Ѹpg����*q�{�?E�w�+���ɹs߹���� �pE�(�d��J6�d��s���N��+$����tҴV��D1���/Y-3g�3�u[�K@X�!IX ����@p�	�Y\��3ct�H�������7�g��℀K��k��7	��;��Ј:��I��|D�WZ��c�K�hlukh��Q�ի�YFs=����vf��L3L�� fr�F�/����k=�/Nf��R��0�!`�c�T���̥=hIٶ�b��ϔsL�g5��)N��(Mb�&�⩩,���.Z��S�T�^u<�qFq^@���:�����ͦ��Mݦg�~�f�貭���$��ILq?�4nô7=�F��ϣث�Vm3-��&�7+�[~~�!+@,8���_ A���6*_G��c#TB���P�kp����_Ab�f��a�)��9ZB�9VB�����r�����ty��n4p�'���}TW1�����vYyZb�]�4<�İS'��&긊��Ba�o�ַ�3N��5agU�+�뉟rB<�A�E��&���;^/f�^�d�b^�U{�򻋙
��aB�-wqu����/�'��G7b���d�	_�������0ݲ�sGw�uQ�
�hyL�߳���*�%)y���~�ŐC7aC}Vx��᜕�?5��sT��;�/��OוW����ّ�o�q����H��NGkE��c�Ǌ�c��\#�'���V)X��X�^��PK
    +Q�H����l  �
  1  org/bridj/relocated/org/objectweb/asm/Label.class  �
      l      �U�SSW���>�1A�x+�(������*��X� J+�rC.!rir��LkY�p�R�Ҷ�.\�Nut�3����@����{y�Nlf��ޯ�}�ɯ��@n0�[�L<UȦg�3gM���s���5��/�T�(�����S�B��M#�3���PQ�e���i��np����t�tRt����	Μ���3��9X]2�Ɯ�g��p�Y��*m���:�r,���'�Ѷ� �+ 	:�?c�C��E��d*|~x��вq�\���a�B�5e��Y+�����,b	�y���ȌQ��-;�2�|�`��M3)��{�見��|��ɫ5��p�x��z��rϛ���-dm��[�M_�6G��
����ok��-?�6�v9�L�JTt(�.���v2O��M��}ZA�� 9?��#W�3V��}��D��M}D�sgG�5�å�mΩ�A���Q���K��룞|Ks'8�z�W3�}m�4*�j�w�=�¼�SU�X-��%;�8�3����@��;���H�8�v���v�<8�ga����z����� .B��i�%?�MA�C��('��E�86��$y�+;Ǳ�ibl�Y/�z��ז�a�V^ߍ�i��:�!ؠ��)��������M����B-�`�;��.�M�y;k��řSV����#�ߠ���c�͗�?�[��|�08V�vs��C�K�'�
��^6�.��{# m��׺��.�)�;��S�5��S��D�	2�rl�<jT]�>x�xWl	��{������+x�9��?�T���5��	�Yti�]4�<M�%t� ��Y���2ǚ6q���U��qS�Q�]��Nz�V������UR:�5���4P�"{8��}�0�L>\਷�+8��Q��Q=#�qi����C[�C��k<�}EA�&$��,/T�k�`�7!k2� ��'M^�YWBل���R���N�4_x�QC����ݩ�R�p��~��OߣN�4���Kel_#뉔��*�|!��w.����Qr?)M&|��]��!B��͆������>��wHvP��+#��%��y]9�*��r�[� �%ܺ�W��|s���6ѪT��}�݈4�'ɔ�0�mw�{���x�h��氱�]|IO�.zXy��&��\�'�9鎭�j�#\��IJ�"9irmz�l�P����c�u�9��g�G���C�{]Y��V����pFs��kPʫ��ʘC󀎌qٰ��/�{x��c+�Qu��?�`DW���K�`��^�`BWt���e4�JdWE�ᚴ�kB�;y�>'(Nȵ_�ďh�UrJ	�D�@u���@`�G-�>/����	�`�շ�
�ihx�)�7]7����c���2��D�PK
    +Q�H�)yC  1  9  org/bridj/relocated/org/objectweb/asm/MethodVisitor.class  1      C      �V]WU��0
��	��j�i�U�T�B��Z��ŏN�[2���0y�?�菨k��Z>��?��9s��1	��7�w�}�9�|����
�*\�9���]���ue�)��,gy�)n˒w �Ys��]�^�)oX{��}��澙���Vv-���[��ܵD^���/p�p
��@�˶�y�H*?�!p+�?��~D��ĥ���("��Ao?��5Ї3�iT`|�Ml��L�r�%�̬W=�\j�C	G�Z��8�Y�9��+��
G�\�\���=�7�M�5�,!0\��t͚��{��5
�{�����������W�Ow	���u���q�)Ko�v�M�h����	dR��f�լ�5�c���%�����m �(��
�np �C�l��5\׀�U�s����`p��pW*��f�f�w�.����l�jY��nf����F�y��dS5�dΫ�t���}gG.�f�*��+M��Ngzߴ�U���GX�]V�����^�U"�w\��(��=,3�G:1��k�&�S��c�ʅr�x��#+Xe�5�H޲K*��T^|"0���,V����*��)e։n�؝���5P#�+wg���W'��?�����x"pNe%�UkaU,��y�K���ݗ����QQtMR�n���d��Gpӂ|
�����T�sX�?tVp�-�S�ļɪ��6R�l�Z��k��J���s��n����u��3��=�l�V�ڡa��;r��D�ߏ.���O���&@t���o��(�	���%�0` $踛�X�%�ӉIg^`Li��)Z�g�?c�7��c�xBi`���Ȝ�
:��L�G�Lc._$��ɘ��L��x����$��>�b�����Z�1�7��Q��-��/S�8��
��H��#�=>f4>�i3		W5��[#d*a����m�k���4�ZA3>ni(M�Fl{�ۘ��NF|����?T��yִ@�(���Y�F�}�a���IS�5�F>j�u�5�VQH~}������a��O�̬�M����B��7J�}pKM�%D_���uB�G�ɞx��-mQi����6t5�۔ܮ�OPK
    +Q�H0?uw"  �Q  8  org/bridj/relocated/org/objectweb/asm/MethodWriter.class  �Q      "      �[`�ř~g����l��M�.�Q�?�M@��0�k��GE���
��������j����`�V�m�l��X������]��=����j�m��5��3��nB�K���ٙw�y�g&~�g��$υ���[VO^�Ґ�urK�����5��̰�U���[oK��\�a�䅩�5��e-�������3����͘�$Va�͞�X�a�Zt:f֣Ԣ$QR(�*]pkݦ�ɍuM�'/imihZ�W��Ai@�e� �J�وq��[ZS��Y.�Nд!N�����Z���ܔ��	�Y�e+��Q��|RД��iKVmlM���(�(KQ6�lB�e3���(�Pf�<�5��5%�sP��C��c(�Q�B�8�
�(Q	��
�V��b��Q�A�V�9�����F��	g�O��j�P +O�X1�z/D��	���i] `�����l���	
�� ͡y6�M#�C��ao�"(�%CdP��O���>^@W��*UR��L>m�@x5]���&��Zj�E~n]/�jJ�v��+�	r&��扵6�@� c�Mj�'l
��M6�ͭ�ME��ʦ��M�TB�܂��c�!��(�6MU��i�����-�	��On�k�0���r��'����� 5,-:4�,ݲ>e,r��T묖�ץ�Z7�jJ^�j��Ҵ�ak
Dnb"7�m6�UDn�i�jm�YtG��X��t)��S��i'ck��6���`h�PK�(+���W�G�(�)���n��؈�N�0q�n0�Be��ZP��|�E��ș���ß����~����\�h�Xq��9��غdMsD3�k�$��}�]�����(��Ѻ�v�4Z�t����u-u�R�h��O�#�Y�r��mij]�jm���}6���t
����u�E�����C@�M��e��%J���MgQ�g=��g�l��	�sYC���l|��bC��Mc�R_�J�H_>T��E��p���9ɢnh_Æ9��T��Mpt=t(@:l�*gB�a�V���)�`GH���Y�d�� sW��D��=�X^s�E�`L�&��^bG�kӅʱ�l�J����DY�s�A%9��M������ohj���q��d�O�� }���+�s8'?}��"�7j�J��I?�E~�D�e�~dӹ�G��M�)��]�9y$46�V�5.�¦�m�O�g��� ���;Y�G�.�~�����8���5e�x�үm:G�~㲿�iC�M�)�����.)*h��=3�C5r�E������qJmkj����z��dS���1Z�}`�t��S�Bٚ3�9��!�8�g� }��몖�q}]�@���"`�I���!l���Q�9A&l�`�e8lbPTQ2���Y��@���@��+R�IEk�`���I��!����=��7��Ե�jU)�[�E��(w#��T��RgHܐ�U���L�8���n�T۴�ymj�u���5C�g8��:ZA�?-5\F]����5��6�[�X3e�P����"9�Tsx��fQ��({�I6]���"Ak������ 3\!}��bZ.���.f
����l�#��e�	A�+gsh�)��tv��8��{�Ʀi2���6s�M��O�����[��*;s�x5\���>���EW�Mz���u֭jL-����~�'�q�t��������yVKK�A�&��}fQC,�9V\���F��V�|��ix����|�2v�(�57�ݸ�?3�GB��9Zy_f-J�&y����2.L)U�o�2����*k�q�SK��*�u�f���f6��05q����h�g��?ln݂���Q����������(Y�rl�mD:��6#�3�r9�ɼ~�̝�'m��<��}���|#%a��a{ACSj��u�R-6�u9j�M�Q���º�8��嶲tMK�m���s��м��%v�N�W����#jp��&y>�ZP���{ M���S2�8��a�.աI�5���5��u
��0q?����4 `5�,[<(3��X��h�U��s�����Pto��r�;T��R���,\tx����T5<�uU���#����g,�R��5%�UH�tzq��w2��k���,�<D���7�/z����0/Þ��Ө���[���+��m:|_$�^�w�W���#�7�r{���8ħ^�n��TSRPx��x5!���LG�
a����0�9�xLjmV}H"&�:c�!^��g_�I��I�l���K����Acr����ڰ.�L/����,kl}s25���ylc]���8�����s����N@�"���
_������+�/U��_��?����'���2�%�u�k֭נ�%.�/~��g`ʜ��oʈ�YFl����go���^���������\�/~�cV7յnla�Tr���_�����4_�a�AX�-������m(��S� C�4�?�A�&1�����h�����SA~@2��z�6U���d�����}HM��Iv%�+>����ug� g�u��CX�#Xyރ�<pU��������&�r�4bG�Ж� ��	��%���fP�u�^W�=�rKN)����eߨxFbV����q~�rT��>�3�3:�q<g��L��Շ��{�L^�O�8C^�9[���1�w,����S�)h'C����fϹ��X���Xغ�xRIA~�C���~�K�!O�]�-�Y��GH8���uP�%�x�h��%�Ѻ>�B��발���iY��督�cu=N��u}�w��>_�{���PO��ȿe�u��Wj<���d�}�����)�>��e}���T=.N��z��/�u��.�
�t9	�=��rp=��$ZZs�fE�М���͏u��cT�fhau7-Fs	/��2t]4��e�Xe��Ѝ�XȐ���!#Cuѐ/C�!��f�̣{(E��T4�M�gZ�8��I!T���X�t
�z����"������ ˛�"�B�H��������u��.]6tЈ��nZVZ���ꦺôٷ5^	��:�l/�:�*o�F۰�;3�cw`f{Џ��Lߎ��K���O�}�U��a���1i��9&\���.�=D|M��,=��݄y��]��-��10��>�EY�b1*+}@QmD:�	 ud�a�ώ4�Jȣ.�ѐ᮵��굎b-6���Z�F��
ɝ�a#q����Y�C�"["��b0�B�W��+�� <F�Q��}���������*��!ߒ4U��u��.9����cC>w/O���L��"�����wPY��d�9V�#i
�����yW\ߠ�zz��Fq�^��W]��*�yw������>�Τ��oF���MǌtR{�cV�@�t!����}{���зK_aq�7����q��4]�F�����}����&D�����U5���^�׷/n7a
�KJ��>�L�ٟ#f�j��Gjr��!G��OϦ�!�qZ܎!'�ј�E�����i�@�Q�$i$y�PI�����b�Ϟ?ь���PnCy
��?(�`���7�a���-ǂpJ���Uu����e�塎��<+�3��4}�7z{$�E}2�p��q�6�YɼY��4-w���N
J
 {�yz`ް*5��{�33�F����gG�h/��d�~����y��o;�4��c+���s���+�-���)��¼��k���nz7����3-�����axR���}������?'�%��~
��zLV��#+zH��&<«n��,��z����$��%^ꤑ�)w�,�%�y�`�>����H�0��"�ÿ�]��]V���!�l�4��ǲ_�G�1�#@� �ɔdD!�;��������਽䄃g��p�ҽT^��_�&MVDol���5buҥL�^�(�CM�c�A'�ۜ�����t��'�\)ʅй�F1���	� <�����ط�E{u��E71BkI5�e��U����+�.�r6}]�d��}�GF"n8��PA�1�E�{RV�-&�]|���?�~K.^�LB���)^Q���Q���ڈZ�qv�d7�6p�C�F	�LC��	����KTWAW}H$@����t����#{g�:�s��<g�����(��#�K2�r����9Y.�
\(@�cp���Zq����#�W�!�[��s6�S2g�I%!���q���lg����'˷5�Xf[��+���#����/��ߓ�����X)�י8�����E��~��!΃��mwh�Z�EJ��}̨s���
��1z�%�L��p���`zLW��7c��^$@�
��Ǖ�D�>��S�	m���K�;O�N��&�ҕx+���zz/�h�[��Հ<��j+��x�m7�*������[L��S������)��q損ᨠ�o���F�C��94^�f�,�N�t�OI��^Vn�E�W�9��4"?��i~� !�4v�4�ac�)�~�rx+d�ҫI��e:*��\��;���0�*Z���%a�ћ�(�,���P)+qY���=0�7��KI�q��_S�{m�c���l�6�E��w���xʹ��0��c4*v��[~H\�^��2�
8�Y�4S!�$�(�NE̽�Xvi��1K�Yi�eZ�}8�)~�ԗ󤄳�D�,t/��\��"W���_js��!����zD�B���$X�U���Ҋnq�/�\��q�9)�Z�1c����zG���un�e
X��#�Wiy~h�x6�خ�oUT�QT�eC{X���#��.ԩ� G�w ��w�(�)O�����va�Yߵ@,��l��Y��iœ�s�pBx-�e�OZ�{�5�*��:>C);A,���d�2��<ooV卓I�ϣ���D�)7�嚌;A�6�d�����X�%�����*A'E�+�$�V:�����>P�:��Yb<�d������.%�{����J�r�ʠb�ܥ���k���,�bV^կ�݋�O�qe�g$]wǘ�ܑ����r�[���
�RS�\S�P����T(rCYr_��r�b�n$��Ǝ�tVaV��|BܘM���-�*8�"��EG��p	�p��U!_EFԇ|��
�p�����b�p����Xþ��|�"�h���Mr��x�X��5����u�rL&��&Z��V&���B�<�}��^�8�|>����l�>�t�M�0nb���f�Ɗ���N��Y������++87����d������ō�T���y�
dl�G�6&�&��P�V����~��p����Vz�a)4.CwA𫠝�)n�Ш熉��cTP&�#��jK�->���!_N�CF��"M="vB-�.`W�=T�R���-�͈�0� #���9�F��[@ܴ���ݴ�Z�F��,�,y���L޵l�������W&T;����K�U�Y�������l�/�pš���C~I�XI�j�TDw���b����{<�|�,� �@�VB�^�
t���!���P!�3��G|>n;v�L|"
�,���`�}Ձt�s��\��K/��n,�+P�R��Ȣ����y-Sg"��4�C��x�S���Z���3�n�iq
;�	���.m��<~�
��/�:/�
E�v���_�pLoa��bw�[L�?�7C�b�(�99��%��(rWz;�)W��S�*�]�lJӔ�� �f��6�h�x���Rzc��\PN���{q��0p������eu�QMٝ d�z�+#����GJ����a+�v�tΧ��g���2�c�=R�]�%�������xޜj_��k9�K��H�ɷ�cB�L���kcu4y���{3i�yQ0�Sz
��!��|���O
ܘ'�c�^����f�Yb�^����^����^�~l52����\!�2 �.T��g���X_!L�}5�wK4�^���>��<�<g��t��]?X�_W.�Z��2�D���R8��B��םȢ��l��]���l}�X0H�;H�l@J;"?����}�~�ϏQG`1�{��r�u��>�>Tm�k��1�2�Λ��)��v� �#F"Q㽜�_�~���>2�-!/�^RL ��O�@ u<��עX�
8�r}l��iz���/M��~:��T��P����?�
�^҂����L7#�������?�7��Q��G���seDd�+_���v��Yi�"�w4r{���}"?x�	�RO���<���,���,��b(d�W�Ƥr�I�����ēm��N��W�TNB��18j���!��(@8��"�s��Ƥ��q};��n�Z����#U��y'�k��nn˓���5�����>$�	�ļjW����7�8߄�m-�B�%t2K���\�.�G�i#1�N�g�Q��-D&c�-/+jy'�τA�L*[����)�c�l��(�j���(�(�K��3�QN��(_���;wG�o�����i�vG�3�u�=��Vr|�<��A�Q�<ajD�D���A�Y����>��J�הG:�#̿�I��2��6�n��_kCG��&ٷ��������������7uf���[d�`�=E������:��+
��C���M��leR�}}{�Ř��=��e�wA���J@04d��%�rq�<���r�F8,nc%�O;u~�e>�Xn"�hǑ�O�@V��-D�J՜��\ռ��Y��l�������D�
^��~��=�E�4>a}���'���$�����ɗ���!���)��b�m��1��4xtV1���Mσ�g<�˼�%{��z��
��8�x��ymt<蟡c��ѭ2��h����2��?=�r��idY8X�G%�~�;_�Hp궩��jؿ�aܹ����l����l��l�r���n:�^Gr�q�� �3������]�ď���Dv��^������!8��V���CS{�	yCcb'�R��e%ABr˧e�~���Jk�S�������ee�繎7s���� �_1P�V�0���<��"�g��n�#���ܞ;z�oU�������v�Ū��ےo�G�s �w{𨑔/\��xFv0RuL:{[}0����ЕE��<�]�PvDٕ��k ��q�QR���b
?�*�xO)�o�z���(�kag6n��%�,��٦�7��f}��I��,��[|��� ��ָf�|�+�j�V���Uw������ukW�Ցm=�m̶��-0�����ї�����L��'h4INz�$K�3s�(�-9hK�-ݖ���i��&	�9M�Y��=!C�9��0���ao+9l�m��L�iT�,�/�-��=4��|�l2-��U�[Q�k�r�5<�M|�9�be�(�23tk[��'��#��G�q��O��|�ބ�1>oCl��~d'�G��N5ozK���PMo�Mߖ�������ߑ��۲�yw7�J�>��߰�ySWF'r�[9�׉�`����~�;���({���Z�T�V."����W�T'9\��dt5��2g���G�r^Y������}�/���X�?3ujﮗ�&[���ܴ˘]J�u[1iW�I��1���ָ:�C���w��Gu/��ٱ��ֽ٩�{,�7�̍��R��WY$n�R�R�6x� �-��gQi�>kT&�w&e��O��ǎvz΋9��Hp�d�����X�Gh�N�KPnP�rqH��o�m.ϩ"�7�ơ �"1[���X�X%t�1�r��N�ONI�4�zd�/KA��8�)L���~��wE�c:�=%�(�N�1=Prg��S�Żi<�M�	Ԓ�>~6�q?0����`o���4�����3���������Gkd�����tL+����,􃪲�Q'�Ě�����=��ŸHt�$��x_�|Y`���v�vӓ�R�5[n����pN�Q#�l���R�v�7T�8z���lo%�B�GsqȮ<�|�pa�^��B�0�_��t���_�C�֩C�1ՖT$�����&�J~V%�'O����r��������^>���q�S+P{.ϣ!��|z�竎_�_�_듟��?T}�����ˇ�␕}R�ϰ�5L�(_�D����}BH�!�,���E���g�T�n@��ABr�Y��P�?X��cƋ��I�ᕞP���
Y�OdNQ����B/��(�YbT���hD䌀Zk8�e0�uF���m�$��B���CBA
��i�X��D��yf�ga¬FJLA���v�ڸ���͔�>���H~��^y!�o���%������=t *o"�����~��������!��ՃH����¨� �?$>����K5!)�ɜ���nV��)�5���2d��G��]~w��F�N����Ww���xΑٛ|��?e�#}�ժ϶Rhq�į��Ƌ�b_'�����t�	��.��D��$_��]�Ǥ�
Y۽ZB�8�Þ�N�Y�����r�/!Ǵ��t_���ŧT�U�3��-�t�G���ȹF��/�(ꦆ
{<(��q���<���Wa���P������}�DCV��X����B_�ӷ�N4,�+��kE������z�x=|�`�t��̢���Ovǟ�n��."|����E��/��p$�����&��Ү����#�z�]XI��J�=�I5����I��*?��f��J�e`�\���*r�lՇ��������L��9���ǂކ+�1/�mBfzM�m�ŏ�D�oPK
    +Q�H�����	  )  3  org/bridj/relocated/org/objectweb/asm/Opcodes.class  )      �	      e�w`u�����fE�N��0�*�����dfٝ]ڒF�!�z/�{�b�QQPl��y�y������}ofwލ�Ǿ�۷���of~��;�i����FttΫl�\��Z���������\I���֖��e-���V:��:�[�jJi�K*���U:\T�)�XO׎Q�2��bM���r���"m�W�!9Mq���x���x����ʋ�S<Zi=�h4��T[f�2�KOΤ̬��ꦴ^^�q��k�(Y��2����2��S&nںE�
?��$�%��<9QoG)�6�1�E(�u,�c��&�CW��X���'���TM��_���M�v�4lׯ�1B�F��y�����d7�?�^��/�.r�Z�,R&g��?�݄�Z��������:6�C�-��agj������LQ��ͦ��U;�e��J�\4��rtWZ���[�NG�J0���9���\\]�\�N8)�+WZw�N�Ѓ�,Ǯ!���$r5�7Kۓ�]"�*���"����}5�L1�f���N'��PI:iDM*���ƴP�o��p0�8���0�x.���.�U���dҰc�E4�$9H�t�^�;�ȥ/�[��b�w��k霈*:R����Ђb o%q������1ߌmڦ�i�ݗsf#�42�3�N�9����T�#���� ٪ �c�p,B+�
F�Y?Ek	̏x/8旒{��>8�j3�I'�9�t_��ㇳ���� Xy���1��1����M+��A,���:Dc���4�FL�N���q4lA�i�n�t#��	t�:�0I�O��`, �R= n��ꀸ�J�3`:`k�t�N�ͅ��Tұ��i֙d��/����l~q<�&��/�U ;��i:��Cl�1^�9tc�q�7��~�D��L5��T��-T��s�ޏ�Q}m���T���ޏ[�ޏo���������x!��q;��qէ�,�ET�ǷS�wR�/�z�୭���x	���R���e|�	��r>_/^��y�]��9^EE��jz(�X�+m�*����u���������TX���Џ7Q޴���L?����a��-�[i�*��mr��r�v�q�`�<�N�`�v^�n�`�<�^>_�}���s�/�4�h-�giK@̃��+|����7G|�7G���T��ql�sr�c�_Vwq\��^���^�O��ϙ��t��F�;Hx��$���	��O��+��z�(	�(bN5��P����4_ׇ���1\���4Ӎ��(Z�q�d�A�1ڠ�L���qڠ>AT�'���mP����\x�S�$
�sJ��k"����e�z��{�S��B��S�NLv�{�@�-O�����z�W{�ޱx�#��I �S)���u�2�2��	�a׸��i�w�2���ф�B�3%^Eoc�e��Q����5̷&��49ʽ�q�:��Z�e��ޤS������ΰ;�x'0��mA����qZÆ�U��C=I���[2ɯ*f�F����ڮvE�zmz9�=m��h3��@D��E�"�l/:�r^t,���"<M��틻ڻ�mKhW��
������]m��]+AKR���..�{��#½���}�
�p?���%������C�����__)|<T�j���?"�Q�c!_+|<,����?!�Ix���p��Hx�p<Zx<Vx<^����zL�O�	�Y�xrh�t�j8*��8\�^���2�o����k��[�����o24ߩ�)8-��|���Nͷ.4_<����Sȟ3��Y��l�3���?B�hͣ)4���<ZB�Z�y�u�Z��uk��m���������E���b�.xI�\*�^.�^)�
^-�^+�^/��(�	�ڷ��[[B���о�-�o�ڷ��w
�w��
���
���
����>	�>�-||��}����
??,����c���O�O
??-|~F�,���s������_��_�_~�(�
���k���o��~~K�m�����,�9���_�"�%�/�_�*�5���
����o������� �����������������_������������?����������������/�?����+��
%�X	â/R%p�p\.��)�{	���W�}�����/��	��_
_&|9|���U�C᫅��E_��)��k�넇��R胔�� %� �>H�>H�R�R胔�� %� �>H�>H�R�R�����o�o���G�}�Dߣ�>T��Qx*���,����}��`��(}�J¢oQ�[��[�%���E����z�����,��pNx,���~D5â�Psa�o����/T+,�	���A�P�P����%���A��A-��	/�W��W	������	��7o�7	o�E����?A��j2����џy��\P��Ω�g�^
�9�OawRX��a
K9<Ja��)��*N��A� PK
    +Q�H	0Br�  �  0  org/bridj/relocated/org/objectweb/asm/Type.class  �      �      �X\[�?7��i}����tU�
IJ��tZ�B�65@�Q� �Ԑ`��ӉsnsN��jg�:ٔ�Xm`:;���ۜnss������t��`��{���O>�s���s�=��sϽ/O���c PƖ3p�}��D�w�/��{B�p����ݻ�=�=�n_hh�׺w0l�@���EC�>_簀�@mk
�1`�KmSS���� 
���5�D����h�'��-[��[	��@#'�8�%�T�A
��"�� ����� �"[MssM��j�����QC}�֦:Bhd����x����M��)��'�<���{"�=ɌsO2䉤O$b!l�L�~$z�����X$Y��J��@���TR�f��ು
�ڡ�40�:;����r;x�X���z?nH_8I18�$8��-�D$ַ�t~1�g+�@%z����C��D"�w����o�j�l�*8��i%�ü"�jmh?�d!�/�(e4�E�4����^��U%�Y�s>����euᡞDd0O0��7gg�ΦH�pl"���fc�������v�,y��ڞ�D���a��;���6h�s�O�b�p_8a�vLq��Xd�ء�����}���1X4����Z���e�`鞱Pm<�b�� L\+W�E�{�X�"�"��K7�`fv�'I6�4�߉���h�'�$i�$����g�.>��/�`/1�"�>4Cіh<��.�`?�<��a��>"2ߘY�s�j���+)>ʠ�(���F����P21܃:��h�A�h��w_*��W����O0ؚK^���ZYv\U9�ЧȊkq���D��@8����\�t^ǖA�x�SW�;i��x6Ё��a�e�A����p�n���pl'�o)�N'b��Z"����M;��Jv��F�����J���0��P��z�ږ�>2ə+��{�I���z��h�/����;y8"�|(�I��q}4��8ʂy^F�pE���&�4'�1�<~s�Ewc}���h[�(CV8���&��ƺc���Cf�ʆB�#1$Ʊ�T��5d��c}Vx����
�`�d����;wR����������>8B��S���������<+|W	�c���|+�^#���4�_,ɸ����d�c�C�x�В�Ҷ����h�������y�~��/�<b���H�BQz_���?�_��:���()���;;�	�'�d����/�%/J������a�!,/����)�6^!�p<�W��U���^'����9�DJέ���7��0p��Z��6xn�,(m�¿�l��+��)Q����xL�#;���D73|��Eñ�d���tR��Y�J<�����`O�7�o�)P�a,������x�m*݁�������=Q� V�����??~ (�D���@����)�3)u��f-�^�bɶPt8L#�oo�����y��RH�'`Al5`�̀ ��Bċ�ĺ�#v�b��D�Ā�".4`�o�!.6`b|�pOV��Dٟ$��e�J��e�F����A��O	�{$��~���n\y�5�p`�{Ns��n�Q��v��n�zN��>1~��2N�a4�NC�2	u)�R�e��Lد$��C`��(�z�(Xum̺ͣx�M�Yɭ��jd	XL��3	�Дʚ�]��Z.D-m����]`9秐q��ȝ��'�BN9���Ü�C�>N^B�9yy�\�rO�U3���4� M #����������k������
H�J����Xy��T��Q�R�QX*&�M�pp����B��DL`�	��`:C:���CP�Luy�1�-�H�{ N�z�6
��JWW~j�:m�g�q��qt�V�q��c���sL�v�
���Z7	���(ScS�x3��[�����q�iU�	u0G��pj�p`��w�62�&�R�rS,���j��]Lt��b�ކ�)cP�����ҷIO���]�eQ��G��E�{
��QM��\cS�ԬaScPh�F�i�����6���X������q�ml��:�]��Rl7��kd�6?
�{ �g�ەzx��^l�P�S�S�S��	�$6�:�����|����H-A, FJN�I�5U��tg�g1��EjW��K,|`�[qO�w�=rW�徛ݘ��rz<;�F��r�6`�X�����RQF�RRƅ2�2?#�)���:Fo-�z/�=���0�~7�Ɯ�� ��6�m�Ƕ�������[;m�ご#�rL��_M9����_O9��x�-�v����ɘ���@�8~���������I�3�YՑ���L��ei�e�el>k�J���,�!��~��|�f~��8��,��g8��n�,�?fB?��i���rz�t{&��9�{5��!yk�;A�6x��4�ܮT�<�c|\�(̫�+^�/��iěUg���T׃�h�v
���C�p�m�^x��$:�ݲ���A������=�&�Z0g*sK>��N,X(�̎�xC/�}�O�k$�5'"�
ޚ��F�Βw��p�Q㿂�/��oɰ8��9dP���RY@*���=)1��
��t����)վ�j-�?�i��w�˯^MT�A��/_MoC���ׯ��@p��_��^��/��5ݏ`��_ނ`��_Ú^�`��_Ě�A�����"���[E������06�t�ME��h\�fy�Rav���aX��i��^��v��e�H��#řG�#f��9��y�ˌY�9�R>4
DZ-��ȇ��t���gV�Mro�媺H/ÒX�7�Bq��r�q1����}(m��9aۯ�rB�]��R�>�Ko���s��qϣ`��ʸ���)����Or�v������3��m�P]4�Uav9͇a��*ǙN���b2�����-�F�V>*�Nef�5�@U1W]]�:N=��W\��_ɯ�����l����XQD�Y�"���Q�4�t�(l1;A�K�~�!�"��'lF�/p�pb���-����q����K��b�r>@K��|�D���KD��� PK
    +Q�H�ALm�  �  E  org/bridj/relocated/org/objectweb/asm/signature/SignatureReader.class  �      �      �UKoU�n=���L�0h����WMIܴ��RCJJܖ,�ؾu9�h<N�+*�X�&Re�f�Tb���+$�`�9��Lc�
$���}|���s�?��Ï ^�:Ù�[�U�Fm3��f�j{��w��&�z7x%g��r�Fݱ���s��n��5�`���c皶S�-K3f3�/�C���p��B�ixsF�a8]f���e*I(Hj�"��hdjW�|�cXL-���ˍv�k�2��`*t
��Nݻ.3)i��$����;O�T)]�0�I�aPN��\��M�J��i�{�!��T��;Ä@.[óxN�?�p�q+Sq��Ȏ8�o�[vs��6�d������ē8�F�R�i����Sc8�J?>�^FJ�H3\yD�KO�y%1�$�E�ᰬ��Py��*��h4�2�͡��S ����Ұ�)��co����t񦘻F+����S��jg��UA���A?�Ϭ4��!��?��È�[���?+��x �X���Ѽ�ڷ������c�e�mؕ&�����yq�+��[���K��!�}Zf��u?/�8V��ͻ��w<k>��x��'2<k�,<^!&���Qj�B_,j���N���8�~D�	�К���A+�-F���!��:,F6*��i����l�\6�ǔ^��F4�d�C�c:�dE��>���U6�T>f���]�Ѳ��$-k]�����'��m����|L��b�_�`o�+��u����^�T�d�һ����o"����C��
'û���}�¾J��L��G��ِL""y;(8�dH񲯔O+ �.��u�2o3Y���B�K�@�N�3$ݡ��������������t��=ˤ�C��Y��):�d-SpG�zW��g棑<��|W��ID��������F�K�������L�P������q����\��g���c��(y��O��L��,s(�r�+�%Cr��D�Ή���=�*�?Y��!�J�z�{Ă~���No0)�oPK
    +Q�H�O  �  F  org/bridj/relocated/org/objectweb/asm/signature/SignatureVisitor.class  �            ���n�@��$nӆ$M�-��:A�( Rו"UiU���$"G�8�}+X $< ����,�xa�=߽��ϯ�?~x���@����FK0?R�F�ւ���'6�h8�Bo̩���ŪD	��>�W��)[�q]	E����tO\b���5���s����N���s~��7E:�Tv�`���=���0;;"f�_A�24*����v���FN1�~�z�.��S&� �i�-7�J���n���>�� �#��y��'qD�7�p���ټyb�F3&�ړ���G����X�]2��%Is>�Lz�\���1Y���lĲ��Txt೅o[z��֖'��	8)u٫-�єqI�(��qf�L���v�CI��S?ғ�����?�~���A`�����7R�˩�v�5Q��j�R力n)VP�r�;�[߰��Q�E�$�wP�����ԗh��2g�9�N;�awsؽv?�=�ì��'���qvٓl��"��Yʬ�b�<� PK
    +Q�H�M~(  �  E  org/bridj/relocated/org/objectweb/asm/signature/SignatureWriter.class  �      (      �T�NA>�Zj��Q��v��@��~!%hb��C]��6�-ʣ�_A.�&>�e<�;���d:�s���s�9ӟ��� ��X2yE+r���qV5K�beM���>+YYQ�����+���i[���-��@,�5IAo薉,A��ܧT�R��mY\7*�ͽ=���.�z�����k�@�n��"���-!@ �ld1�AO	�S�!)��Q�T:��0�5��^��F�ۇu��rZc�+�~�B}y�,���z�X^FY�^�L���;L`�2��wp�@�]�Z�6�fS�|�d7��&P�>�x����h�Ir'�V��xI���vxH�ۏ ���pB�t9"���^3�k_�����nJc�6��s~�P��^�,L�uZ��V+��C'�����=
7D��v���晗�W�5fX��m�m#N�BЈe:wK �\�q��yXw��Z3�F�>q\I1�x
�ɳ�.�c�����h��2�� � �j��z��з{����
�#7e�rpW��#$t
<��gpgG���`�>$愩�1�$G7�"_@�"}�]� �_�M�F=p����S=��g�ɠ�>Ef��'0!���3*���.jR�Fڨ� NY4wEK�|Q<�QRب��x�{슯ʘa�i���y/����U�����o��wO`���)L��g\\N�FQ��66��;zSr���cH�ѡ�ퟪ���m�$Ü̞��!�X�촟�u�w+�H�z�.|b�[��)9[tKU@��Ɉ1I�o��+�z#�mJ�4��T{8��eG;�U]��7PK
    +Q�HNL1��  �    org/bridj/util/ASMUtils$1.class  �      �      �U�n�T���$M�vY,Y
-Ѝ4��:
��t�nefm�(�$ǾIoq��v�@H��<Ő�:!��P�s�]'�E*?r��}��7��� Vq����z;�A�	�������pq5�p}�s�]߶"��e�op;����VxX�r�0���� �	���:W���p�_hr�2���­^ۖu>�~���|O|˝��>��Ѿ���[��m�]'dج�H��ky�XIcg�NEo��x�X:�n`y����.�C̦���ܦu�f��kE����|�DWP�?�����ê���}l��;Y�3pF��b4�pc<JYn���y=��oe�������k̔`�amV�L_B�f�4����ȃӼa(�Fs�7�"^�-�L��W1'm[d0,�i��`�r]����7i��V@U�\���=�˶yH랚�|(������x�
BVǢd��SZe8�4=p%��fu<'M�[��E��y!�&J�:y�W�|YC���G:�g3Z1�Fwxh�����	M
3�S�����q5�6`gsT_T
xǥ����ty�3L�0���������*�]�g�&rtߧW���QD�$h�w�$�ݳa�]��\h4v��k��<H"���l�-��w<��Cj��#c0F<�5::�]hŢ�j ڧ�}�qw}�	���<ŅZY��Ze�/�"��6��C���P��y�*���gU�3Z�&�����}�V������ى߱p�W^�_�ai@u7NO��QK���:!M�ejdB�B�BW	e�S�Y%iZe=�,��/��*�'�Z�l@�Rr���Bo�ZKș��ަ�M��|I{V�fOR��8�2h�Sh9a��v ��i��wH݀�C+MU��Ee�R�6F�=�U�?,���r�[�
J��R���*(�
J��n���![��W�"���U�30i�)^���
TWS,�PK
    +Q�H�;ame  C    org/bridj/util/ASMUtils.class  C      e      �W	w��^�Z�-pAI�m9�I�vl'KY�88���hlO*�ԙQ�J�ҽi�ޒhI��ܦн�����f�؎��S�c��w���~ߛ���5 ������5��YF�L����`6}���h9��U�՜Nɝ�5'��-<�$Y ������~�4�_�}\AM��;3�M������lY?�ۚ@">�h��OhNr���%��c�4%o]�.�6�ih]�t�d��n��^¸]�ٰ�ZF�p���k�)�!�Vl��Ӻ�5�傞Q���o�]��S
lb|o�U�B^*��V��9B�ƨi3�5�0J�T���{�=���C�%��G�\7��N�D��[ê�K�a)׎���$�J���DJ��5�h{vI˒Mv%g�T�6����n�v����o��G��'�\�
��ۊ���,uVA��~���.�%S7�{FcY�T{ ��C
>�[#X�!���AbG�O������g�傪r}|�A����a���ԗ�Q���3�Sz^�BZ BM��s��w,�uY+8������u�@�������DԜ�Z��t�Ȁ��O��b'�����0Nq�H�Q�6\k]\֕�W���S-k;[zE#�R�M����@����)���q�RI��~Q�|>[q۠PHŗ�K/�4���I�WrG�9=�T���aN��k��0]�W��l>+_Һ3Sb>O�+�(;���죙��^�Q�;�O�A۳��rD�N����r���,s�VʴMv^<���)|Z2|��yI,<�޵�C���O/��A��I��$~q��V��
����Nw���W�Uσ��45:�w-�����)y��j�;,�	ڳ�d	�k�N�l%�I䓆3��5��d�ɨ����A3��H�6b�<�|0^��7����A}�0�L�Su��1J�ԑC�5��%3��ޔ0~P�8�I�n?��R��ώz���'\�O�W������/�Aʊx	/�x���,��ˌXil�A?[���uս%��E9�&#.�����	���M��04���(�}rH���k��y�ܤ2B�L����������jt.���4���]W��i���~���l�o���hK�
l�i�2Dvej�8�K����k����ڸtk9w��X5��	�'Է��r���</�p��4����+�c�ct��g*Ŝn�v�/g�Y#D�w,֔5�MթX$���z�$����������͌��Z&#�R���C���L�6u�x;c���^�	��?�-�Upt̡�2����U�M��p����Ny��E>�0��Z/`��}^g:����`��Rg���esz['�pW�W��+HTq_�_��*Wr�5&�^�0i�C����j9]��%*ɌJ�Ϋ8.@�9�H�eB �um�߷/�h�-]m�ݽ�Dt�0���y�ـ���'$�uw�[۰���Q�$>��t���$T:���9ht�؁<t��y�R����>�i�P�����0,�e������1\��ߍ(������������G� �����D �Z�����H)���-�����ᏚђUT�t�DK�A�l�s��R�3|�\ŗ~��9�|}1�wy t�nq��	��_4������͂��#t#�8�/�GсQ���^^w��|�h�.6Ѹ&J��?Lw\��Zf;�F� �e��_��Z���K�9���Gh"�j,t��罡y\��s�Eo8����[�1,Xť��� 껞P�g
N�~�q��/8�&9�t��O>�����|�3%�q�O�{��O?��TF'�S�@� ��_�w��p��❮�cD<.?"�7QƉ�Ql�;,�
�Vk����n���ݧ ��5BZȵ:�?PK
    +Q�H(8ұ  �  $  org/bridj/util/AnnotationUtils.class  �      �      �W�OSW~N{{��**����b���2AQPdt��^�Ғ۲��9���m����d��b2�,N�`���ߗ,�G�som�%�ql4���s~��{y~綿��� �qE�.mOF&l+q-2�����T*�5�V:u�3���k��F$i�&#g&�����旎�+ee���M����P�F@�^�2����]`뤙�O]5m+kL$�����gz�F&�^�`�W�t����M�Sf*�>^t���Q�7�xB`�*v�V�3c��7�G�l�q��}��n��K�S;�q��	��V��5lX9f�����;!�H��f�iL T��"E&j*_��P+Pee
TC������5?�M��$�+:,S-u��Z����8��&�è�n��G��(N�����2Y#g���n3:�:�e�a���4�X_��1MܪƦ�؇�����L��e�]1l�yP�f���<-9a�����%x��H:��&f~w66��@ެ@'��7JL�������Q�@���
\��j������Hͩ	��p�������a[�I>�Y�S�����̴i���!�;gY%^$�K�G���IpOLh�{5��{/of�'���6��Fr�ԲGܾ��R���`n�z�1
0��vؚL����:�c����$�J�r�;\�Q�uҴ���2-O��^�u$p���W����+�փ�Q�8=c��>+ib;�h�o��z��1~�p}��X�='��=�.
���:+-��{�xJ_ �WB�Js�16�q�u췹�؄�9� ��5؂����g�������;�'�ɶ~6者̳��1���Q�j���a��<����.-YiX|8�.èǎ�q<��������]�����"	KG����a�cy�Q��>��$�x���/���ޖ��5��!�Zf�S�̢*��　�@���>���3o���&�A��փ7�c^��p��*X�V��fH����9nv:�W��(��8B�n��\{�}8��d8�v>�0'�d�����>HYGe.������P���`ng�Qyج��Nh�Ef�6,�^�������)��2oQѢt�8�sC��Y��j0�Z�b�b��잋���\$q�߆�Hğ���Z��SBʓ��U�j�w;BJPm�izHs�Ι�=Ed��Z��>1f��H�E�!e�ŝ
��S���k�Oqj���[@D6w�f1����/�{�31U�bZH[D�������$�������kB�<QhɛLQ-M
F�+�F���wȑI%�"��:�m����c��<g*>��(gR���,0����y��G��Ĺ@+�)�,��;��!��&/ ���<'�7A�$
��d]�5����1I�-�8�i"�gi=���q�7��-|��>�׸�op��|����reO�ә��PK
    +Q�H�S�y�  �  '  org/bridj/util/BytecodeAnalyzer$1.class  �      �      �T]OA=�o�
�
��lKa�o�!Q�Ic������tw(C��dwZ�7_��M$~$��QƻӪ��<���s�{�ܻ��Ǘo Vq�a��f×���V�1*ay�x�r���s�I0��ia��uX��T��D�!;���;�a��$M�����%ԞgWe��틀�q�2�w�fU��m��!���m��`��"�V�0�`�Wϐ�p'�Ő<@P蔮>��[�a�xA��ҕj�a>?Hr<�P3`��"30���:�͇�Χ���ړ$�\�ԮQÝ�B]^�����������ǳ��b^c_X�h�<h���=]���?L��u(���l�+ö_fHɠ�u�i�\xf`3i\�,�>XEs#K��<��m�o�L���B�k�c��,���L�\�ʘ-�a(�5pi��Jz.������ ��9 %��%o8�i�0�V�+�ۭ��{H��}K<�ڽ�Z�ϯFe��c`�!Fk$�	'���#D���,��u�ޣ���0^,![����u�Z
$7&0I�Mz��:�K=�7�,L}�շ�)~�x�+r�(Y�j=V���K��(F����f_�걇�"J�K�5��e���2Ɋik��Cq]ψ�Ր�r���-��m�c��q��1�":KJ��H�PK
    +Q�H�~Bp    '  org/bridj/util/BytecodeAnalyzer$2.class              �S�nA=�ma����ZkQ�]�xW�D�6!�zQ���;��ˮ�0x�+i�1z��P�o�M�`$^���3g��3;�|�`w�c���J�e�?�hы�(���P���9Ov0|�'�H+Y�ڴ�ހ�9��'y�R_�C)���E���k��~ȣ�������d�C�$�B��֖��ݜ&\,b����g�ú��2}�!�PFR�1�z3�.JKȠ��w�rXe��Im������&��w^�?�0�<�D�t�wt%¸ǵ|��V�Ft}�}9m�S>[��KT(���� /\\��".��4ZTD7�P�M�:�X�}�v�L|V����>u��Q�a�+ɻ�xf&�嶌��h�*e
��H�ġ��Q/�
�D蓘�w[Q$��iD��tu9z �R17I(C��e0�!�Shl}�J�3�}��f�4���ӺI#o�>�p1u�:Ok��+�/���s���d��fjb�nX��q�/a�P֢:��E�p6l��(���{[����n�P5-� [��OPK
    +Q�HV��3  '  '  org/bridj/util/BytecodeAnalyzer$3.class  '            �S]oA=�ma��o���@ѵ���65i����;�C�]3;`0��?�Dc����2�V�`$>���3wν��Ώ�߾��M��@����n�j�9�ZtW<�7~#T���Xv0x��mJ(I��|ȭ>q��%J���Џ�>	�#>!��j+:�x��9�ZI���'���0l�*�M��u�6O�X��=��5�^E	�P�?���/}��J����5$P`HV��<��PbH�Im��OY�����難��B̼X�j3����.��u".��EW���g�;��*��٬�s�"w����=1"��sp1����$�C���Ke(.VE���Nѝ)"�J���ɷH����\I����hbXoI_�b&sUW<�f���zAH:�M�}_(�����S�VX��)��<��p��=���L}�36�_p꣉��lS�Ӵ�h�3����
�NӚ��F�+.'��}���M6c�m⊑�aWM��	%�Jtױb�fL�[d��F{;��`�n�P1n�"6��_PK
    +Q�H|.*��  �  2  org/bridj/util/BytecodeAnalyzer$EmptyVisitor.class  �      �      �T�OA��^[(�'�(W@�"�(�
�>`br�nʒ���m1�b����h4��������{ۻP���tv����ٽ�>�@������i69sͅNk~��{����K[/�N����A��$#��_�9��"�;���_RǴ�-sѵ�0��8�zj�޶	�CAr��2�0��9�T̀@@7�R��P,`��	LU�R�,��p	��UM����טMyv0T� �E@ce,!��n&��V˱7{X��!z��5��(�1#�R!�O�69d��K��7�y��͙�s<�s�TIw���A�EX�N�7"��~3FZ�V���y�`��G�nly^||��y|��R�pˌ�u��c���ȪT>���%sr��Ａ
�u۞P���7�z�SI�4�N�vIEK���}��V�َK�
���0��4��H!z3�L�)&��!��&�.�+�'�[�2���q�s~�����4�b�>8��m���݅�õSЯ r~����Q@%o NK@�|��Io�BFzC���;�^Vz��R	��|��"\R�qd:IGXB*HL���}D{���C�Wz��R�i���v�(�G8Iy�O��j1�W�Z��=��p=�D���A%#y��&_�PRk8��3������F��8L(��8��U<E�*n݅�vMzC�A�\��&�&�K�����p��������L��;��)yQ�O\�����eB���]�PK
    +Q�Hwyq�  �  %  org/bridj/util/BytecodeAnalyzer.class  �      �      �W{W~O��l�M		,�[�I6l�P�H��6e	Hh0���i��,����kU��ެ�R�h��Z/��$6���<����_P�sf���I���d�����~���9�����^�M`��Nǧ\+u1��,;>8�I'e�{�I�� �/���m���'�.�IOC�@[��i&[r�љ�7;ne-�!~�@�xF`�J }Vav��u�0���(P�J[�a��h�x�Ѭ#�!%Lb�~��i�5<�y��.8�1k:mx9�����D!�C����w�3
-ae="��ˉ��8�D��x��ְI`=�GҞ��ۨ1c
�
�f�<�JO�GЁ�:j�E����mx�;���� ��2�]��.�%�6ܭc+��G��WYVF=�6�q�I�e,%G�p]cV.���)���꽗:�M��&�ⴖ���܋��dq�6Uq+�[�״��ᙩ��sT[]1��Fv�_tʔ�4��\�e���z֐������e�@]trЯ��:�p�����\�t}v�k�����ò�K4a���r��Bo+�Η��γbH� ,Tn!��>�(�u4�!�I����5�0P���6�G$�c�p�$�� M�Gq�{�\ޥ��ܷ�@���+3�L��e�)�r&����.�1����(�,�~����S�:�L�ܬy�Y.5�JSU9SRG|�S�"8�{>�C���K(h����4sƌ`J�6���H�s{th�bE�x\V�4�gI�N�Y'��U۫�W��⏞J0ػ��vز�Q�vr�T��~V����l	>3�z�jP�1��l����r����NUn�r��z:�9B�Q
�������ʔ^�ڊqk�<ŋ	,�nG�
쾈/���,�/����0����k%"�������7(�K�����L�IS�FE�kx�>����1��.)�|i�39�� ��:�ËK��n��h~V)�K��ܵ�2<���m�/	��@'r^B�+:���l��@�u%d�
�D�}���nr�ky���ɈR��u��#>K�N���cy"���p�<'A�*�[��\�s��U�V�%S|�������#m�69��IH1"����Vs�i���_b-	J�=n��1e���
����hnf�t�=ߒܻ���J�	Vr\M�O��9�d�r6��%F�;>�Tv�ڀ�~�/��r_H�8������)��zMUI�MW�7�����a]�k�gw��W����y���A�y���h�F��'�8@��h���
`�m�k�ߎ�~�'�{po�S�f�G^C�(�E��3@�3鯱�{�� rO���=���#CQ�`������3k��w$W�{�"�&���y��ს��h��|bG�c]G�;F�gz�4c�n�搈�pjU8{}�|8�A8rt'�\�z��}+�8E���Ϗ���3	��9�ʵ;���'�8_F�=R��%��>�k���OI����:�>�֎�����.u�t�u�z0~�#���D�<&����>j��0�r$��>UXr$y��,�_�1ս�g]Oi5I�O�+�h�D)<�i<�����y�C����K�����r�G�y^&�Y�|�ϰ�Zs�ΚC�yOs|Vİp�VU��Y�|d�B�	ЮqN�ȑE\bO��r����sǻcsxj���ع{"�h�*�Ƥ�U�lO�_��]>=�9?t�F�If��ٸ�ķ�l��N{�ϟ��U�"��e��c.�w��@E�{�-�{�*�rUyY����&���'��Aw2��E\#�W�o���h��B7��mcI�q�?���*4��L�/
�}��ś��r��̯�6̯�_�7�j����ɽ[�[�VH���iy�6��fnbDQ�μ�QTWԇ�}s��$�M���zȫ�xi^6e!G�8/��J��tun��[��7+���_Ԩ�}�j��]��Y���ɿ�PK
    +Q�HӐc�   0  !  org/bridj/util/ClassDefiner.class  0      �       �N�n�@���$�����RQ�R��:��:��E���(�|T��(U��������������\�Yg���.Ų���J�Q��B��(���ǾP��$}�7��մ�Ɠ��2q�M>�-�bm�^�H�G�����!D�T}:m���&:7�U���*��o�[q�6�TmBnC����ȳ � =�x���F�_PK
    +Q�H��G^  �  $  org/bridj/util/ConcurrentCache.class  �      ^      �VmSW~.	$���T��b���U!`�P_�Xߪ���M�l@����������8S��7��~�����������{�yy�s�=�����Q�/o/����[I��L��-�d��r�5}Y� 2����+ښ�65k)}#�"ugda�X�H`�VYA�["�RZ���eF+��f9��B�u!�
4���U� ��i�o�I��LS":������#�#c4��ifI��Z�(��G�Q�{�,S��W��[E�.�N�8�ӵ�ɜ�}
4:��Ʀa��o��X`f≅(�p0�f�7�!�������M8�^�S��Ag�(�|��:���vQ�J�tu,��5U�5�k�tYp��B�T��{��&���F�6�ߘ�]�G��`8%pdG�ND��e]�Ţ�5�[�{Q��P���,{�(�}0~O��#�W
�B�.Y��*}�����۰���3'<��ꀁ�|L�B�rrQ+�NL��VLW�ca\b�i���r���x�KO]@&�2����a�L3�k!�|V[��ami�	&U6��N�"���bZ ��d~�ίk�5Ri��FpC�I>�ަQ�?m�\�"{�҉�?�8���(N����3��u}����B~.�;���Ŝ|L�L�.�a�ے�m|6f����C6��f"_�@�v�8�"D�żz�B5���|[��L-^��0.l��.aY97T��D�<��b��[7�fG�W����a����d���r����w�"�e,��Ph�3�,�)����sR% ��.h��<�k��>/l^�6,9[Z�J�*�i���ѫ�k�n�isJ��,F����m�e|��_=o~�??s����	C��NY��]4��c�]3�8��5�yj��9���~\Q#�;@�]���%O顉kW�z���{��{����K�~q<緻�İ���˺����~�}�}���A����U�|�?��*�����,&E�-&���c���K$��1r)���hS�`_���k��}�Q�������-�/Q�2>�����W����� ���s��o�o�6�T�z�O�:�0����"-��e��.��(��A�ì�����Ҫ,�)�5�d/�]sw7f���W���R���mD��5ƵG]�*g)�*)<blUR^U���jU��(&�&o;&�X��m���uT�Nː�I�ű$w���h����`O�Z{�3/�<8����,�;qO(�>�Y�N5àw�
���`q���Y����Y�,{�&-ke��t�V7��&�o1�m$Hl w|T9��UT'��$��2��ھR�pC3�}�q}����w6��^����񿼶��GU��Ѳ��{wm�nl�~�ZZ�PK
    +Q�H��,(  �
  -  org/bridj/util/DefaultParameterizedType.class  �
      (      �U]oU~��,�]�m���`���m
�@��¶|��N�i;e;[�Y5&b%���z�&�pÅ&�%����A���s�L����b�s�{���}����OO �Ť@s��̎���t�����1k�,�Ӧk�X����Y��o�ZQ�M��;f6o:��S��֘EX`g��Zy��e�#[+o���1�h�%�;Y���@���ZR�S��pӱ\y�\Y,�7}�u]�c{=�T%�J��a��©������M:�X_�:b����ϫм)���s���La�x�%.�q�l�y�s�k;ļ&�~F���E�j^o�Ώ[n/�фMT\��Q�h�^W:���8vb1gg-g\�5�Vp�nM4#%�J��2������@tŰG ��C;�=1�1n��d�����+Zd7�J��F;�?�t!a�"ad��NZ��rcҐJW�E�@d,_p�����чcq��5�.N��jK�b`qʞ]�ؔyc��0n�y�1��2윎8)'cH��>�4eL��(~S��u��Qˠz�}c]g�w��t����"��iI�K��e(W)R��1o����Y?�D�0f�M�6G��yI6�l�*Ό�f>'~�PtǬ~;oa;}h`�#!���	�B�UWk���U�1��J�1񢑙G��:���2���a���e����I�B�Ր�IaX��"B������[;����
<��m�k���E4��5��o1�C���R>��k�8�;�P`�wjK}�1�..b{���K����v/�H���HF��#\�O�3��+���FŹ����$�-K'�}#s!���2��j��G��+xUE�y�0A~'��T�H;���FtS�0�8�Z�f/g���{C���Gq6kv���A�=�����E#��å(j�� s����}�S�&=Bo��\%w�Ls�O�[2��WA"%�I9d��l`""�Z9�F�mҁ��u�W�H9��<�e��\��.�g���A�<��
w+H{���6�CZ�������P����p��~�l#Jg�����N��q'{�o�N�'ϯ�n5w��^#�yJ8�hm�3p�������BA�p��%b��/�j��3˛�	?4���F�tW��R�>������Mv%��w��-��}�?�.|�[>Y�c!�e�
�%���)���jrR�MŔ�����uRum}��wh��Ij��}�9Jj�����4Y�g��~�-��a0������J*���zj��ɩ�ߛ���H��O(�)���|��s�>_P�KV�+b�5���z�b��ܥ�	O�oPK
    +Q�HZƾ	C  �  0  org/bridj/util/JNIUtils$NativeMethodsCache.class  �      C      �T[WU�N�S ����Vm1	б�DKlmjմ���!��a�5s�U�'>�諮���������_Q�3�\�t-Ι������o���_p��¨��Ez��o�����/���OԶ2�p?.�j]93��2��;{�j�����UkXx	��1��Ah7ֵ@�f�b��R%y�-������R�F�D:��5�|7��m6�f��g���Ν�Uudt8��dw=x�q1��@�K����$����9�=L��@
�̭����4_�ѡ�W�j�2�K��W���L��P�)��<^uq.�Pǭc��Ὰ���*r�:���[�JO%�C�~I�lO�K:6$r	o���7ɿ�����6*�&d6���Ŷ��x{W�ae�rN]�e��$���2V&����A�������\�~�l�W�9:X�T�͌���I��A�A�а7ps�q�P�X��f%�%�L]�˥��c|��!��9ey��̐�w��a�=�}qH�CS,��M�n߲��8�g��pO���NY���e��}��)y�F�&:�I���&VecWFZ�5�C{��ׁ*7�T�ָ��d�+/F�o`w߭�ͨ��j���@EIIU��Nq�������&1B��iʟR�=��_!����0��3��K���s��BV`{�_�;\���X/�~�����ʩ��#x��?����w��>f��5���y��1>��@"���T(����|��i�����E{i��4O񶴷�f�,��>N�U����k'��w��%E���	J�2��պ���.�wbicu��%}ĳ�H��8�����8�PK
    +Q�Haa?�n
  �    org/bridj/util/JNIUtils.class  �      n
      �Wi`T��n2�y3<H�`� na�5
�	!P��@%�̼$f�gAp��ڪU�jWܨVŢU�v�ծR�b�X�ז���w��L2��c�w��|���{߳�<�$�E�L��Nj��/eŶ7e3V�����b>�>����N�)n�M���ь�SO�4�i��$&��42�Ns��tb�V#:h�P&�8�A��`y����7�-
G�v�"�ʤ,{����Ѵ,�E]�n4�;��c�E�YJ��I%�x^sc��v	�US��T�r쮤����8����me����߬��� (��Zi��d��j���׊��@�J��ʀ�4�mX�+j&3���Y:��Q�jnuA�}�e$p�X�.7�~��1g
f#�H�!V��g�t2K��1}�������9�-;c�l#�7��N#��y�n�N-M5���0ҙN�^��I�b;���:)s���
J����L���@fP1�M�B,
�	�
�^��B��6�ߵ�_`F�mr��'םO��A#��Y�Ե�o�ь9�����1�̇$��J��,��u�+�2�7`Q����H�!K`ǎ:1s��ɬ����c]� 8+3rA�[_{G
m��X�ӕ����г]�4L����Q�J�,C�k���i)E*m��xS�h.�w'���K�r���T��ͭ)�U.��L�ے�(J+�U7.���#�Og��jBj�E�o�ڗ���%�zu4`��iH~�M�.*��H����QS*��U�ǀT&��gWe�xL�n{ ;d�+3�IӦ�E��$��$[�p��ӕ�����.GJ��%��4d��|+��q���v�
쒡��13e��	_k��F���0�.M��� ¶�	�;Y;��pT�3���	7�w��v8��K"���8{��ٝȃ�f]�l������MLB�S�z\�s���[e_H$�!��!��o}q�����0߅wp��:�ӧ���T�x�<��ߎ�ig
&���nH��2cHDٙ�7}�ȁ�N�5��V�������.ƜO��{$i�ƽl{t5}�M�F��)�c�3�8���noq3&r��_��<(K���H��J��I��Ɏ������Fv}&�Lmڝ�4a�l���G� �c:�ǝ��xD�dy��:$Qvw�"����S���=���I�G�"�������8��s%�D�,�<�T�c^&����"Ӭ�%�P�l������)�y^�<M �z6���E���1<�a���Q�G�_��+x� �5<W���A'�k�����R���|��U�3�ۏ��U^(���q����E?��T�h�a�c��e���c?~�4Vk�Y��q� ������V�/�<�ܪ�7�6;I�;?~��7k�#�>:Q��X	s̡�g:���.^2f,5Ҧ���� �o�sO���\��F�j�c [Z�Dұ�	$at�GR�n��:^ձG�R�kD�h����h<���zݦ��B#=(���, |���G[�*������E�F��_U���p�.��0�T�$�hT64Q^�3ym��AܫCW�qϹ�{��]����O�꺘�Nob,�����1��Ӫ�o�É��Fʒ]w���B�mvf},fw$0�~P��ɦ��ZK��m�m�T��i�eA{���A@���U7�o%��j��r��P�g�z�!�'
5O��b�	>��#�<(��9���A��*@�)���oJ:Z��<�)PKΜs5���[�O��Q3��0|=�|fO�Qԕ�������2�W��_�D%�ULr��H�y��sU����&�8y��s�T��xiͲH����X,����Ol/*"���rX6��;�}���W_,ytH�5��
����`-�荔J�j��G7R7a_B�[x]�ʔ^H�n>V�L����C�0���A�#}I�b�s�.S9�U��Qo�
��Nײx���;�sز��'�m�"����T%,VCC�[≔VQ���h��j�6<�E!o�R�yP�s�����|K�Ii�r�fo��#3�-�S����,�h�h��!\���Be9\۬��chƺ����ۤ5�%��+�Rz��|9��e��.�����KCe]����5b���&��{$i�ݤ)�+Q��(��O�M��|<��s̋��(��fl��m>�A☆��JrЯ6��������H�y�N�;h1��<;as�r�M�b������a7�ǕxW��5闍.��%�(Er؛�x4Z��t|��K�%�u�q?>���4�JBv�Af������>�M���oxry�O�g��5Ty�m�և�C8��ǻo��}����/��>������(��~6�.Q�60O`�>gb>���� j�)�i����;�͵,���	=���MUÍ��M�w3?�ob��`ne�ܦb��E4�󲟨���Cx�!��t��W��5)}SJߒ�w��=)�@J?��O�����K�WR���~+�?H�O��rO�G���{0�o�MZr��I���J95$J�����]�?f׶1W��k����d�,򰆼�G6����j�f��ً�r�ъ��������j���#0�9x )d�Cޑ.�W�pհ���a�T�@NL;����}͉�âꐨ�3s�z�)��ǲ�CX��i�C(��a��n���~����ۼא<�r#��6OK^q�:Kdw-!1�PK
    +Q�HMw§�  ;    org/bridj/util/Pair.class  ;      �      �V�sU?��Jh�G�-���iVh)�����VZ���di��I�$�:*����3������KtFʨ3Otƿ�g�w�ݤ�RGe:ݽ{����9������F��|Ϝme{*e+�3mXv�4���rfb�X6zrF~�gjn�̔��.��FQ�d��T4lc.g�O��ꟽ�7�����$4�F��H�l�8j���ɧQ��� ���� �4
��n�j�}(H�4�$�w,�T�(Ҙ�F^ĥQ�df
�,�����[���Ʒ,��$ҸO�u�M�M�6�v��0yh�N��i�F��U�(�e�4ju�C�7ˣ2��x�-�03*�P�A��d�1�KUx8#�n�4�w� 1�S;u4!��O1
���FAJ�tPbSip����=�5��+Ԁ�����O�+�*fʶ���/����^6T�rY��r��6�Ӎ���`�&ק+�h�Ѽ2է�Y`k��nnj˛�|s�:BteK�hT�����|�\��H��)���G�������[�e7�,���B��F?��5��e����y�6K�x0�V�\�)\�.��%@voj�"�����S�����-�-�Y��`��s�d�{�J��\ND
oA�4�T,�0�0��6Ͻc���5�7���dn��B�ȥ�b���y�I�R�P윰���Ҝi+I8.���O�%�o�=X�
$��u���O`4B+�7�*v��ؑ>�ϛ���Y�HyP$�W���i4��j�ﮚ�$�;�� �}��x�L>�=�·�/�zH�!�g�T�z�H��y>�a-nB�T��� �����3�P��t��r"�V<9���������K�
eq��ݲ�0Q\tC�Ť�tL�D�~�W&Br\E�����f����)e6����2{]�ёjڤ�iF@5cq�.��ժ���3�_�����[�۵�?nt����7���� *��TO�Q�1'S�sg�P�o5�	���顁�7䏭�ԥ�uj�B?����<�]@v	��Ix�@4��#H9�D?N�p�T���"b��$N^�QR��d����?��O�Yv�6<��Fσ�#��xCmǑ�%`�ps���eU����������y��N_{Dg"�k�
Wb��##���8��X=���7p�*���nn�L��g7	�j&a�&��{j?1;������u�vt��:*���cN�-'��+�"jc9���Y��T���Ꮭ���*����~����\�u
zP�����y�*�
��պ�{U�^�jt�N��<5��)U\F&�[3�.�%K�6s�� �d�����v����3t�r�;��|L�I��c�
)���o����hJ�"���t��)�Ў���fc*����?�>��T]Y�d�M�i���;����=������Q��[>�L}D��1��	��)ݤ�`�s�5hNcZѲ�7����D�o5~Y���4��K<3��ץ���a���A�WYY�R[9��~��Y5)Kv
�;�b�����$���w��������@�oPK
    +Q�H��$D�  �  *  org/bridj/util/ProcessUtils$Kernel32.class  �      �      �P]KA=71��h�֨�� ڇ.���R��Jp��h�g�A'��03�g����?�?�xwmf�sϜ;g�yx��mB3��abU�f^��¦]��c�<��H��s "L��@�Z���{җ]�L���§\BX���
c�X%V��CBe t&	c�Cg��q���4^�����6�m�%K���EBk��Q�x��ߩ�o���_���(��0z���_	�ݽN�X�b���a'~�� s��G��<c(i�
�{Ei�g��iW莰J$Z^��+#ϳ�D�!Sm����o*?�Z�Hi���4~d��Nv�S,>1&�"尉�<�J�8k�B�ĵ���~��מI,��u��h��8V�ʨ��B]ak`�Q	�����4w�����7Ǎ�HT1�PK
    +Q�H.Z��9  �  &  org/bridj/util/ProcessUtils$LibC.class  �      9      �N�JA}�I2�4�K�^�xP������{Ϥ�&=���<	� ?J�=iC���U��������aj�Ad�ldN%��Ici��� T��:�A"�<��2v><B�7�$����A�u�'�0�g��J$�$PL��C�G�PΥ	Ց�ʝ�ãi-�5P�:�ݣ����?�,\�K��fő	�����i,��0JD���?B;TZ^e�H��N�.�L,/U^�&ZK3N������vj)��*&_h�:�T�-�(����8�7����X9~E��o������բ3�:z���C�`W����i��&jp��:��-j_PK
    +Q�H���v  a  !  org/bridj/util/ProcessUtils.class  a      v      �Vk[G~'D6,kŠ�X[S�H��VC�BQ�T�k7��&���F��k��^{��{���� �i�~����h{f�$@"��y2;�9��{�y�����o ؁6["M#5�;F&:$�$��4�0��	����f::���IGA���~�҅a�
�Z�F�GA-�_�ZVr>ʅ�3�v*�c,��P�e�����&�:�A�j~�EI�q�f�_!k��1͝���t�������!X���EKd�c�3�Q�LY���yZC6�X��k�1�4�+h&����Ⴁ=/�ד�m;�_s<o:F��4܍-*6��y����hT�"D<P9�LۤIACS���������"M��Tb(\��4�zf�˰#3-�*{B���
�*Z%㚻jX�CF�+h'���s��� :��fx�� 6������p���+7n�4i$՝*�.���B\-<�"�=��w�L����+��$3 *�V��I�# ^"��(��\�j��t�;w���#`$y�\��$�X�u�u����r�ͣ:v�����r�������A�ZO���Wl��8^�!�_G2�IR�{�I)�Μ�0��I��B�:�g��3�i��j�"/M5���<;Uy�Ou��
�y\��eGC
�'M2,g�+EC��ϐ71᷍+�+�F�Sv�.]�X��c�"g��Ta��M��2)5Yc�R�����Rax�>��v]5bHUY�0]~K.eʻ����ڊ�&�eX���5y1�ay�A��߲ܿ� 7����Yt�����Ë+]0�����I�s�T�*��
�R_�j�Bv�^Sq�k؎T��&�+]�Y]�x�jX%�r���wd�w	��)Cб�
a	��:)iK�����}��*�5�|՘��>���00�|���q�X).e%�̈.=��'�@�7L>��&��,MKݦr�u�F�ԝ��yW�J�T�O���Z:<���*	u�ʋ$��b�L�7	���C���䫟���]�d�\�6�5��ć/hԊF4`-=���T���c�C�^�n�h�Ŧi����wt��
*����h��9�(#ЋZ����G�~�G������U�5=�ֱ���#2&��Y�����K��]<�+�1x���gp���9��a4Y���8o�V���}��5�1���h���>d�����>?��w$2��w�����'.�L�j\�v�I*d�����1�+�F���si���x���&^��_�uk��ْ�%���Kҵ���:��9��8�a\�q'q#��S��=�o��*^���X��S��Ǎ��?�7�E��g�V7G#T䇣����A�J�Ct���>�g�&W���]�;K���<}�]����y0�����l~pc|�	�"����PK
    +Q�H��?I  T	     org/bridj/util/StringUtils.class  T	      I      �U�RG=�F3���H ?b'�X	�(A�rldll��#��4�PB�F��l�a�l0���MU���&�?�.��hxPL߾}�{������)p�j���-���j��r�X����Ś!е�o멲^YK�,o+ujO�Iu̬����'60�
- >��n���ϔ��ͭr�d�bK��q֦Yv�J rZw���jX>�S�V��-�RH�.���C�d�KWb��څ�]D�W�6��c.`��ET�^��˓ݲ�ږ�\6*��$�&/�������[z�j	��8�Tu���02Ҫi�h"nŖ
��Nm[���n�D� �0�>l���)���p�쩸'������
�D~�=�m'i�|��E �#-�9��ɺa��e�ⰿ��G[	w<�P��=g�6�%9zw������k�)wv?#��EL:z"���v�C�0J˹�	^�u�6m�T���b�0َ�x�A����!t�Q����H^�F�e٣�TV���D��,J�Y����1�v���ecӨ�iui���l6�=�nm.�W��[}[�������
h5["�70q	E�߬P�����u˔G��#�Y0+�tcsٰM����֡��h�U�zâ<76�9Kp�w����A����:P�6�c�,���A��Q!��ί�]���ꍿ��W
mX�7�T"�v�+�0 ?�:���ȿE���Rr�Uޥ���V��_�U���vm>On������z~V���߉=\yu��9|�\�5���>�u�!�,ċ0����*s���]X}�Id>���-�b��+跱&x����R�������(uw��+�;3��[���H�:E�F���2�{�q�C�6���>��G�8@�y��R�t;�CT�c�����q-�����ȑ��JZ�����ި��� %��Ԩ�;�݃�����B�����B2��ana�����%(��S��BQ��.M��!�L�X���^L�[��M�����6�
JGI�E������K�6��o�$<����>a�S<�������)[����!c��-�����Ԣ���QsN�5��m��?PK
    +Q�H`�ݪ�  G    org/bridj/util/Tuple.class  G      �      }TMoU=o<cO&�4qk��Hm�qR�i�B�m҆8��*���xdOd���
�ؠ�	`�Ħ�,�T\	D�VbÒ5��p�xj�t1ｹ��sϹ�������dpS�X�QNni?�n�����A�	AL��w�tծ������V�s8'�Ԓ��v�����e�`֭��U�hr���@ 9�cB�a@Ũ� B#P0F�V�m22?���dN����^����z��0iP��g��("��\vZ��H�D'�_��1�b��u��0]��S�>瓶]mJ�!�
&^��봀R��e�<��}���`���JΧ�6%�h27�N�]�ڦ6�U�n5�Z�mK>/�k%�ヶ��[-9��[|�ci�����E�q����VH$�_L�C�lobYF0����4rEFr8�W��z)DX7���<ݠ��@�c8�	��{vu�n�v��ܖ����[sn�?.:�bl�ۍ=gí:8��P�ɰ�rJy�y�1�5Ƿ�+��L+���M��h�G0x'� �6��p=M�3�:�aN��9s�Ì�u�Xva��,a-�Hy�#>�7�Ӹ���������0m%:H,�1�)��1����e��"���g���v���|ӄW���*d?����}R
S��H�P��u�3DY�I6n
X��^�'?��_���.���H�
�kh���/Pnz��L}+m��jD���Q�
m��c�S��LcZ,���JU��}U�̴HEg�hX�	$y
�˒�O���+u���&�0�,����:�K�R�*=�,F�¶\��Uz\c�ֈv�17�c�7o�m��-������>n�?$�
��)Y1_�~�����z�r��Y��Er�9�4�ݟ�鮽���H���a^����]�7OܥoP�>���Z}�>�W~�~��������/<����J|��O����Ԅ��F�y����]o>�H��up}7��F�@�M&���$E=�ϜO��:��M~��G�ޡ<�(2��Ip8�w��2�S�w�ˡ�PK
    +Q�HJ�,
  �    org/bridj/util/Utils.class  �      ,
      �W���Nv�M���0D"`�N1)�MB8hjH���f�lf��Y0*�*��¶��m=��X��K ���W�}�������3����&����>��|��}���� hƇ��pӀ��oJ�z�i� $	��ՃjST5�����"v >	�ðZ�$���nwH�ՇwQ��?J%��=.aQw!�m�5{���qm��4ⶕ�ئ�C��Q�֬�����fKX^�=놥E�GS�D[�KB�G�0OBn�"Q�ҍ�Ψ�w��ʝͶ �Q!c>B��X�*r=O)
b��D�KM�7�hfa}x_;Kp��S-A�HX�0O˲J��Jە�U��b�b�'ʄ�=�f�f�FZ*�sZ��7���B�n6mJi��^�ovs��\B ��QEF4�f�2��*�qVK�i��W�D'��i�f31M[���5��0M�5մ�e��&���V��I�ٶ;GT+Em��NP��t23"�Pf�����S��L��&m]��Y��;��� :�M�,u,b��$(����Ͷ[elƵ̷%`����bG=�1XR�x�6D���x�>lh���6l�Q	Յ:M@�)v�,����>��߱%����7��X���`WvBF39���2�� ��7	�ώi_�-��k����xq�3.7%���`yl�mlV�I����&:{(�[ė#�u���7b��T���-��0kmK�h���@)0�p�t[dӐa�ѹ E�A����*�Uw��37.Â���(��L}Lh��ȁ>�s:�*Ê��6��8�ۅ7��棲`�$��_(A�J��"QcDW�{���_�vkB��DĴ������s)T�*#�a����̓@DA��N�#�%���I�y�vmP�0�ADm��tVlm����a�E{eM�,���<G� �vEx����])a�E������#./�����Do��[�4i�X�:2d
�T�9Z.�ꝜȞ��"�����}��z>���A#Ŵr�9!��V<B�93�R�8!��3����(	�{�ڡ.��!P_W�IW8)A���2�����V�Q�G�FT�+�K���w��0y'����C�!Q>+�ˈ'b1N?mp{L�T[7�-�E����TV8n;mJЊ� �e��S5Ӯ�G�F�e�֊�֖�v��iƠ�U��)Fy&�^V^ˑL��GJ�HH�X<Fr�4eؙV�eL��8�$�M!��Jh�X �i��TЛ`:#�m��6�no�m���\�:����-U�Ɖ������Z����v��	-���l�X�:+��3š��	�h�/tu�7/����S(��b�U���MP��X捓�u���X�U��ijb<�5�p}��S�[7�m��r�;��٨�#�e�����5?���?M����ĽU�5VD۪G5\ƪ�!~�C�V��7�����.VN��E~��|�MȘ����+qv�QF�\O����+I,H�^��Ҟƙ�j8�y�����O���9IF��\q�P�K�.�{�cֱ˱�.�������3.W-��3!G��^E��ɿ����
ϱw��(���5��h<��jw�:�&�lv��I���w�&���r��\��5b��.[�h�u�r]'}'srw ���]��1�����7��F�	�x�\ëg;�E'����/�c/z�bt�`h��6ª����Z�y�e��>���T6���p]�dړZr��ou	G;��nZw����>Vx���7���ړ��yV����.bRN��J���3����&UJ�#4��=����lU^B��TB7L@�b�V(����b�)��	�s��	�)��R��-I+-ޜ�Z���]��<�T+o�$�d�+�W&1<Ip�9*��?���$4c���y�s/�8������厉��i���랆��p
��1�;��3;���a���܍�R�b��s��\�;-�s��o��;�w'9�m���H��ENa���MSC��	�N*�1��x^����w*&���*:�q�V�^V�>�| ]�W('����>4�b�h���hff�v7��W%pjt���W�k�aIc����xI����K'��a�'Է���c)��u|��e���37�sw�_~z�c��S��v�\u��%��� �y�����{��\��<J�Y�-"���D3yŒ�R�I7�r�i�x$?-�����{�O�Yg�7��xQ�^�t0'���i$%t7�Z��4���q���M����$^?��fdx����g��ʒ���3%.i!����:<Źs�S�iN�	6�	���u=�F|�t,|��y�{E��*�+~:���)�,�1�2\q���$,_�ڟ���;領��L;gJeO��c5�(5"�G|���3&�8=d,�/�:����gK�7aJ	�_;g�lcL�~��3�`��3�g��o�n��M�[�
������m }T��09Gu���<u�{�oVff���Sf:��˔�-����Ɨ����c�~������F�bT�OD����g���<�W:�1��91�<4�/ޤm�_����י�������&u�Emo�|��q�w����/�n�� PK
    +Q�H����  E  	  w/a.class  E      �      �T[OQ�V�]׭��A�ڻx�Zi�[mL��a�1�.�����S�4ib�c�ljb�֤?��u�����93�|s�s����G ���k���H��h����n�����7�Ʀ�_�Pb6%�7�8��N+�*mjBclᾄ)��\4�2��C�hV��6Y�s�f�C�W���eb�d�����s�Vu]UdmQV�
�l��lX��-��S),6u���rj�y��䍬N֮SkRU�����>j:���U�Pf�[�R֌2ӂQ�jm�MSŬ���kUE��Ԟ�����h ob2��<:xxxxyt���ǣ�C{xe�|�x2��Zٵ����=_K��+|��މ��=���K]�T��������(�̝��U ��'�s�L���R�H�hO����v\��G�'%��IB 7%t1�DL�Cܸ��m��ô{"�ы	!<F\DF�a�Ƙ�db��G"�x��4�i}�]��y�nu��د���5�7o��4�'�݇�]:Dd� O�|	sz�v%� ��I�@����&�]�h�"�D��E��T	���pڪsY��d�Ӛ�x?A�t�b�"�����g�R�L�%��)B�L�V&�U}]�csr��x�/��֔/���������K+�6+0�U�v0���ƲuPV��#�.+p�3��_�w�������5�'�%�ڻ���hA+z���*��S`p?�/�a��
l����<9nPK
    +Q�H�6ot  �  
  w/aa.class  �            E�[W��� ez/R�, �*����ĴXX����{�cH"1��ʹ�'��|���s�νswg��.�H��k�~[�rЖö���o�[l9j�1[-����-I�����Y��� �s<�E��\�X�Hҋ�G �C�a�~�2�E�!��u2�##�(r�ͭȕH CƑ	$�L"S�4Bf,����p`n�786���,FN!sȼ%��)�X$41�����4A��Ck�AށK,!�Ȋ%	+�@�ո�	W���]�\ͺZpqu��J�<��{�Ǐ�#kY�Ǔ�'���`:m�i����r�|y�ށ͏	N��}������4ɒ�4q�l"��%�|��($��b��(%ʈr���$���D5QC�u���F\Fl'v��h$��f��h%ڈvb��� :�=�>���&z�!b�!<��&��Ndp/��W�K��r=q ƈqb���1M��b���9b�X Nb��K�2�B�!V�5�F�&�f��V�6�v��N�.�n��^�>�~��A�!�a���T�JK����T�V'� �$��+�;?��������h`.����x@'1O���E�%����(��|q\�G�v�u�ڧnT7���-�Vu��]�K�[ݡ�T�Q�Sw���=�!��zD��v���u�:O��.P�����u��L]��PW���[���u��N�9�x��d�F˂-8q�y��\��E�d�ḳ��Sqoz��N܆��!����?aC�X��b�\;�׺|���N�i�<�������Ir��먶�?��s�d'�\�j�c��%j��h�Gݢs7P�r�Dl�+��ͱ�9r<���(���~���Y�Eub�b�E�lS�C�17�%��bf��������駱���Z��?�j��_P��$SE-6{}��l�Y�R3�J�y�<Vp�P*�e/�T��J���2J�y��I6{x�֬�J���u�)o�4���nx|f�-�F�6뽍�d��Ai6�xe�y�Ŭ�>J�� �͔Q���tm�_�/��PK
    +Q�HF���   S  
  w/ab.class  S      �       M��n�0��MB��O[
�}���#�LLl��(
�}�N�:� <T�s3��wt?[����7 K�	���N��*���CR�'��#9���0�&.Mu��i��k����坢�h��FK��4� � �.H/��xr>�^r�.���)���p�����^�>�e���[>������˟�m˟��Ǭ�sƕQS�_�D�h�?PK
    +Q�HO����  �  
  w/ac.class  �      �      u�]OA�ϴ�KK�R�O@�~�k�6%$����&h��jڮu�2�l��W^����G�[56t�8�l�ygg���?�~��+�l�v���5֤{
�Mi�K��>R���2�Pay�ϴi;��t�a/��*�N*q2����4�ҿEk�@ǜ���~�9-Gs�����e�E�)��XVlN,'�����
bE����KV<\���P��c>����z🭐�N1m�`¨��|��}�C�:Uq��IK�Ys����nMj����F�n]k�sJ�@��/b�|vl?�q���a���(�|Gc+':1#Ӎ���ƩNMl�
�f`u:N8m�B�?������"�"����S�1�F]i��ȹ�#�W��3�]����,��(�>n0\���(��-�"�͂ی%׌Ʋl2�.�%�o"��D��/t���ȕ��%��wd�Z��o�s���g�K�k�e��K�@�PK
    +Q�H��Ö�  �  
  w/ad.class  �      �      }R]kQ=7�M[MM�5���|�k|M)Ԃ	(�ҧ�������ҟ�SA����l�]�]��33��ݙ����� zx�Pl�G
k��w���&�Ą���DD�g�S��T_h�m�OÉS��$�ǉ	���K�w�(_�ٜuJ_}�b����������Z��tM�E�ܮ�N�
��M���.L�
�����?N}�k�Y����U�7���҅�#�Z�u"~�H�m_��K��'�j{y����m{����VMt�t9�8��Nb{�u��*�֙/�Ȝ��,<�6v���OMd��'!�mr�U4P��|Y�����Z���W2�=�[�'��^��#{�Lm��x,����3�d�U�%�F�Y"���W��c3/���ʔ�\~/S�!H����Vw���[z�%����ǆn�[���Wx��,:��?PK
    +Q�H>�gWz  �  
  w/ae.class  �      z      mR�JQ]�k�M��~�����sDE�/>u�#vƣ�g�$�}T��X5k�={�=�����8AY ^�4R5��9uB-�Mt�����H:}���u�絍@��N+P��sg�a�|7�#�r.��H/N3� l���!aC2�ɓH#��t����7���N�~U���yȧ������S.�{L��?WsNSg�K�3J��S��JT����I�=�2<v��E�Jc1��XFɆ]n���p���Cmԃ�P��{�Z�F��@�Nu�4��C	+R�$�-pȷi�:1S�)՘'���#��&򤩨�)�U����kl��ef_��l҄�¢=u���a�;Qc�9���E�v��1r�zEq���f�|PK
    +Q�H��l�b  �  
  w/af.class  �      b      mQ]KA=㪛�e���ǋ�ϊ A`,	��4�&#�,��F?�'!�Џ�Q�p��s���3��� ��d0��C�-�P�#p0&L
3����Ծ�ܱb��`j�1��}�c�C��]���Z�	�V_�Ć���C�Y���Tn�b(��r)�n����p�	��������{Ԙ��I�mK�P�#��_"m3naÉw���y$�t8Ȣ�#�ɪ+B�U�C�ģ;s1�ܮ���J�rΐ鋩�*\�c��I�I2�Q�Q.�=�)��MJ�8b�����B?�#A��o�6,]�nP����d;QE�Y_��%zZMW��ha�r��0ް���J��t|PK
    +Q�HB��   �  
  w/ag.class  �      �       M��R�@F���"(ȟ��tj��wh�����1&F}.*f,| ��Tw3�̞���ٿ��_ /x��OKA���y5Ȝ8�"k�!)y#y'9)��}�d��,Y��t]	���e>�JT��W��*TE����<�E$�5ny�l����lW~T���n��b��b�p�`��f�Lwء�Kvd�ˮ�������}fz�n��b�L����5��y�9������8�#PK
    +Q�He���    
  w/ah.class        �      }R]KA=�g�w�}g�=,=B�!��4�f#6�X��z������Z(��pν{�{g�����;�c��|U q��2%Q&$Q'D�p�;�ٶ|�NG�sUo�#����S�U�����0?������.����(��������c��~��$RIL$1%��;\{J�/
,�D��Ω�����r;MƳ��T��9{6n�D]�]��7`��mю2��U~�.��5<���m��ID ,��=K�����Wnzڨ�����qO���4��]��[����|;X�2 �������� &˘���%fha�Y�$ָ���al�%z߂9�[�q����*�4�#U�~WI�TY�� pH�\��=�Ⱦɦ�	�ΰa�6U8��a����f�i�PK
    +Q�H����w  �    w/ai$a.class  �      w      mQMK�@}kMbk�֏��o��C蹥P�P{�K�7�l��,O��g�G���R�f�d���ُϗ7 u�3䪵.�ݔJ��d=�Ґ?p/�j�]��N3�a4�z���k%w��`=� ӏ����ϑ�c�߻ˁ�`�A�aџ4���"j0,��r��v�QF�T�����Q2T��}#���Lӟ��d�E�E<��1��M-�p��]Pʭgp��~��H��-b
̸��n����i��3�D�	x��a�*QZދ��e/m�B�5ݗj�k9P\'��.���1=�K~��f	�Ȝ3��@���VI	��	�X4�-�9�Sc�&Z9� ���O�Ú�
�)�$9EX8:νb�[c�Xi��h�tf�p�0).�D��_PK
    +Q�H"	R?    
  w/ai.class        ?      mP�JA��k�5Q�_ x���! !�����l2�	�,�������(�g�(�Cu�P���������K�|�3e(��z���N�K��^��»�b��8Yxa"�Ko��l����G�`(<{\��I�<OS`sPr�8�8�24���w+E4�����J��KsK�E�U;ۈ���V�ߢ��G�C�!f�Q{pM8��F񜎫���(�i*R��C��|S��07JŚk+�*�P\g�������sz�Pn�c[q��X0�հP�q�b��҇C�d��\���o�]���\��MҞ�r�V*��PK
    +Q�H�w�  �  
  w/aj.class  �            mPMK�@��4�M��j�����sKA�PP,��i�.eC�@����SA����FD��]�����|}0�%������Die��1#"�b�a"�&��b�2� �6a��u.L�����D�KB�9��氅<�<x���W+�o�L�c���!�S����6S��x��U̎Jf'�yy��5MT@��}�Ԗ3���y��C��z�K�UQ"��N�0*�[B}�6Z�<����`�P�	|kp?f��ssˈF�� �3�.N�;أ�b���[K�Q�����{�3����PK
    +Q�Hy�m?  5  
  w/ak.class  5      ?      mQ�J1=��P[kG��]��떂Ba@�Ѝ�L'��1�L�.WA?��oFD��8�$9��ޛ||�����jw�šTR�ؘ�	>aFj��n��ܽ�b��(��~,��;�q2�?Fa��D0�]�hQb�r�,[6J6*����H*-�C��)Wʽ�"��ѕKZ8�<3D'�x��w���3b�=/{���r�ȁ:(����#��:
h��}��|S��~(���4�2RK��D��I,p�=J�Lz�3�UH�	�1�$�,c���Ʀ�Cb��i�~S0��UOW@�������v�v�j����Yo��q�sn~��PK
    +Q�H=p*  �  
  w/al.class  �      *      mQMK�@}�4��_���y�֏C�9� � �x�$K�7�n���T����و(��{3˛�}�����`�k8Z2tfRI=g`�b�^���ϹJ��(�f��2��R&���e��^��g���!f����q�e���R��y��!�e�x�?��TZ��q8j����iC�l6{�Գ���C{�h��"��N*��Xʕ�rq�T����Z1t2U\W��%���,N��>���)�[�p)����MBm�� �_g�=���żr-��ѽ-��xb�aw���s�8� PK
    +Q�H���  �  
  w/am.class  �            mPMK�@�״��P[��z�֏C蹥 �P(z�i��%�@�i����?�%���"9�{�̛�y����`�k��,	թ���4gF@h��Nx�Б�����IyA�µ�0i�2?De'�L�{Ol6�-���uQ#t�_��ڻW2'l��C<&J�Nl�A����ώf�#�8�dƚ&J [�u�ܖ����E�)�Fm�RmU�[�#�J��P[�H��78a�ʼ0�o�9��*ED#�X.�j�'�2<��b�/�[Kw٣Ľ>9oh����叟_PK
    +Q�H �$�D  Z  
  w/an.class  Z      D      m�KK1�O:m�>�Vm��j]���n)� 
��n\e:����f��rU���ěQ$�sN�/7ɝ������K�ݙ1�RI=b`c'��9) 	�#Ce����Zx��R�5C=���`�Mu���ȭy�P]���ʡ�`��s�e��\]�\l3�&��q��)�`@״���H*-�yw�&����[�{{�Ք�3�(��c���uPg��Di�$fr%�P\)i�e�V��\(��X��:�yP%���*Q��c�P�l`�"o
��[6�GQ��}�a*�&�j���t78{1cK���:���,v{�68���2c�1�PK
    +Q�H���w%  �  
  w/ao.class  �      %      mPMK1}�ڮ�նj���[?��-�BA�Ћ�lJ�5�m��.OA�?J�DD�=�7����||��⒡���*#��3�	Ab������+~'ra:&[�8S˄�l�/�Pވ4�;�\�} G�Q"���О�Z�[%�eDs��{���Y�������g�vXP;L�-Gc�# stTCmG���,i���\[�$�j��T^km����5Cu�VZ�<��B��ܾ����^{[��ħ�"�N�R$�;[䂤�πr��w\/�ܡ�ZPz����5��8� PK
    +Q�HW���  �  
  w/ap.class  �            }S�n�@�Mܘ�-����[�B!��;$� RP$��ҧMbt]�uQ?��JH�|�t�ZX:g����<ޟ��� �Mz%(]*we�J+�%H��7��@�>� -��FR��ݡ�3X���=@��|�n��CoǄQ��3����	�9��g:_<��F��$�RLi&�i�)���R �;RLH���[h�8��Kg\ʹtY�r���w���k�r֪��k��<LX��Q�'�Ro��C�׶�+����� �5�����I����db�fҁ�v�xpl�3��(�jY�GϘ�8͠��,4=6R��d\���6j�僧���ց�F�$hvG�4Q����k�rT�0xX�<XZ��X��N�OM�g-����u�9K߀��t	z��e�Ӗ�@/Z�
�d��g-}�r���s���K-��p���26>�+��V�!'��|tY>�-E��������:B7�D�*��.Z�>��t���6�15`[�3\��=�_-.?���\I�V���t��^L<���D�PK
    +Q�H��s�   �   
  w/aq.class  �       �       MM;�P��v�@m�������_�y���sY�Xx e�G�nf��������ł`����5��{,(!i��Y��˶�4�yd|��Y�l��I �\���T��WW�J��jy�X��#LH���ݑD{#=��2tҡ���C�PK
    +Q�H$s�  �  
  w/ar.class  �      �      }R]KQ=7��~&6���V͇��sD�B!%�R!/>�$���x�ş� ��%=����҅sf��afv���p�@-�l��S(kܡ���M�1$|�g�!F
K#}�������?�N�F�׏�p䝸h2p����OX'w��(� ��2BY��P^�����=:E,�TĊ�j��͏�X�Gm�r�T[�E��N9�j���[/�t�~�˵�ۇ������ � "��h۲�zZ��|����ְ�M�,��{��@	��u�W}����^8m]oz՟�̹�3�?����v�"��X�&���`��*�,�}�+�1.$�2�b"�Л�c���&���*�,�f�9~����	��Q�S�A��WJ�R��KKH����:�r/�i^%�z>P51�Yq�=ʖc���q��M�B%�MH��I2��F3{�w�؝j��j�_PK
    +Q�H�.��V  �  
  w/as.class  �      V      m�KK�@��4mӗڪ��w}��"t�RA(n\M���	����\��(�ND��9'�w&w&��� �8g���;�l_H�lH�$�4!MI���3��N���\�3o�ja�;n$�3g��x�~@f�������[�)�1m)m�������6�F�Ɗ�5���we.�s%�`ڣ��M(�򢞞�e������v����<Ko@=%����Pǡ�#�2�Ҍ��X*��݉�p�B�Pq%B9gȏ�/��#�P�u�q0��[�r��:D�"c��	�S�&�A�3�M��	T)
&P�(���>�D'�*�]h{�Ƌ���4��)�B�c�a{���3�K� �PK
    +Q�H|�f-b  �  
  w/at.class  �      b      mQ]KA=�n��e�٧��ϊ`A`,	��4����,�����I����;ka��{/��{�̝���w u\2�˕�FSH�Z�C��0 �c>���ˑ}�b��`d����
f�Cs>�y�g��8�6L��6q�S2�i"i"͐s��|!�4�\J�|���dH���]������5Z�����*QD����P[��6kN�Zhl��AL��r8���t�i]�ǙT��뉩p'^[J_q%|9eHv�Hr5<�c�ʀ��6�(���2�(b���4�BBA��o�6,��Ȍ겣���D�nFu�ӗ�_5]$hڢ1�j-���%�V����/PK
    +Q�H7��1    
  w/au.class        1      m�MK�@��i��~���j�o�8��S
"��b�O�f)[��M�]�
�� �8Erx����Lfv?>_�qIp��9�<RZ�1�&,�
XVHh��Fx��K�.XɅ!��d��
W��$�����FD�$�=�:�X#kk��5Bk��Eh��*�>7�����F&��������r�9���4n�5u@�ZU4ql���Cާ�j���\�U�k�c#����P���&M$�p�e@\ɫ�����U��Ρ�v9���7��y3�5�P�o�y�W��#��m�Q�X��74�8�ι�O�_PK
    +Q�H�l8;a  �  
  w/av.class  �      a      mQ�J�@=���^�jmj�_^zy}n)A�}�Ӧ	aK�@���Y>� ?J�M��&pf�9gg6g?>_��pŐ��G!��2�>��2�|����}�L��b��з�P�S{��h�~�̂�"�!�d�E��@���C*��g��4�5�g(���!��ʿ�\J���9�#��K���)����}j�4�KR+A��>ԓ��������9Hv���G`:�P±'d�u��cՇH*���\83�'e����3d�\E����1 :I�2� y�B���L�Ei#�ئd�L�����XP��[�Kc�[�?�`8'�n\���/��j�JдEʹF3���%�V�զ#�PK
    +Q�H'��4�  "  
  w/aw.class  "      �      }R�JA�ɩ�6�#�9��爠�YP���$YÄ8���g�$�~�X�Qfq��{�k�f{�����!�bM u��2��J\���Ixĝ�t[>J�#u˹������A˩��vnL�m��B�Qv�ܗ�9�� ��Ĭ�[��&�D�K��i��1�Ƥ@��U��6^P��J��� �O�s�u�̧\��`w�ݑ��[�Oƫ�W��We�œXj.�[�s-FnݿC��Q�e7z��-����f;�e�Z��q��MN}麫���j�A�;މ־�F��A`�F��4��C+����	���_'&���K!1\��Kc��e{��	��	3X��-�#��2K7�������m?7�~�N"gN�L�a�^���([�"l9G�}�T��a��>���|PK
    +Q�H��.$  �  
  w/ax.class  �      $      mP�J�@=�4�M��j�k宏E�:� �P(�q5i�0%N �T�UA���;Q4�s��9�1�/o �8g���Cc"��S6#pB��Y��S��&Z��f�<�\�+��b��	{��B0�}�dQs��48����˕�H�F�dTx�_��L*-��,7�"�ÿە�q�v2
����i�f�]�У;����9�+��b!�2JťR��Zfj�М�Dq]��#L'��r2ҫEy��3�K�F�?�*='Du�
��[x��K�K0�G�k����zE{��/�Y9��PK
    +Q�Hc�~}  �  
  w/ay.class  �      }      mR�J1����ֻV�[�m}X|�*������v-)5k���|� ?J�l��fafΞ9�!'��|}p��@�Tnd�J+s, N�!�&�"�D@���|�~O���-#P��ߌT��ߘ��2?F�Q��\�z�� ɦ�$,%,%-�,�-e�~)y���ݯB�M	,��J���(�G�\�6��w��G'9���u�����Q�e���#�=t�V��)�m��G�R1�el[�����6��t��F������D��H�B� 0~�:Z�~��.<p�H�K��Q׉��)�1C�x5��Yʘ˘����yJ�e,PrX�����,2�.(`��qZ��g�L�T^��?ko�.�a���$߰�aͰ��PK
    +Q�H<؝�   �   
  w/az.class  �       �       ;�o�>C~F/�0F6�̼�; �\?�
L%e�30�3�02�i����'e�d��g敤Y�tIb��Ѳ��0010�v.6N�4�9?%���383=/���(�A��(@�`����	10!���v�` yv ��3!H^{;D�l
 PK
    +Q�H�U)�  F    w/b$a.class  F      �      �RMo�@�m��u\�&��.���&�QQD��*U���*��֖����\RA%�̏B�6��v��x��{�����W ��uQp1+P�Q���8I�Ԩ�@!l
�>�td��ʼ�A]���w"���H�a����=!��I�4���2ӂ��+��}��(���=V���Fz�t�*XH��#���S�W���S;}�9(7�ρ���w0�`��'�]�fǵ��G/���(�����h�C��l�?���q�^�a�s������>nXX�M���1�;>\��PÆ��xX��}�e�bK�؍���n�3#�9��1s��U��k���Hf�ʰ�5���e��!�TP�G2�ȴ�ԙ�͝�wT?�U��������́���M[�b��\�vt���s4*3�4�*�0A��o�O���k����Xb�%
�O�B�GD�q�c���PK
    +Q�H �r̖   �   	  w/b.class  �       �       ;�o�>C^F�DF�ĲD��ļt}׊�Ԃ���<F��RVjr	#s�~#+�TIdg`bg`fg`ag`ed���A(.)��K���A7�ZS���ni1#�g^^j�sNbqqj1#;0�42 �17���ـ���q�I PK
    +Q�H�`_2�   �   
  w/ba.class  �       �       ;�o�>C~F/�0F6�̼�; �\?)Be�30�3�02�i����'e�d��g敤Y�tIb��Ѳ��0010�v.6N�4�9?%���383=/���(�A��(@�`����	10!���v�` yv ��3!H^{;D�l
 PK
    +Q�H��٣   �   
  w/bb.class  �       �       ;�o�>C~F/�0F6�̼�; �\?)	Be�30�3�02�i����'e�d��g敤Y�tIb��Ѳ��0010�v.6N�4�9?%���383=/���(�A��(@�`����	10!���v�` yv ��3!H^{;D�l
 PK
    +Q�H�{���   �   
  w/bc.class  �       �       ;�o�>C~F/�0F6�̼�; �\?)Be�30�3�02�i����'e�d��g敤Y�tIb��Ѳ��0010�v.6N�4�9?%���383=/���(�A��(@�`����	10!���v�` yv ��3!H^{;D�l
 PK
    +Q�H\��գ   �   
  w/bd.class  �       �       ;�o�>C~F/�0F6�̼�; �\?)Be�30�3�02�i����'e�d��g敤Y�tIb��Ѳ��0010�v.6N�4�9?%���383=/���(�A��(@�`����	10!���v�` yv ��3!H^{;D�l
 PK
    +Q�H�P���   �   
  w/be.class  �       �       ;�o�>C~F/�0F6�̼�; �\?)Be�30�3�02�i����'e�d��g敤Y�tIb��Ѳ��0010�v.6N�4�9?h8gpfz^bIiQ*�"+P
�������b`B6-����*@��@�gB���v�<� PK
    +Q�H^�)g�   �   
  w/bf.class  �       �       ;�o�>C~F/�0F6�̼�; �\?)Be�30�3�02�i����'e�d��g敤Y�tIb��Ѳ��0010�v.6N�4�9?%���383=/���(�A��(@�`����	10!���v�` yv ��3!H^{;D�l
 PK
    +Q�HkG�
'  �  
  w/bg.class  �      '      uPMK�@}�4��նj���[?�甂%�X��ӦY��t��.OA�?J���������f������V�7c����z��n�1�|����Ŀ�b��,O�(��꼘�/�^�յ%�1�Á���	��\)f*	�֯�Hc�{��]&�y`v�m#��˖��-��A���`L�*`���Ñ1:k��t��}��|3��Q*.��4�2SK��T&��"��>�`&�J� !eMʛ�[��\�%g�G�Z�*����xO�%�&ڣ9�n`�����g�Y��!�PK
    +Q�Hҋ�ͣ   �   
  w/bh.class  �       �       ;�o�>C~F/�0F6�̼�; �\?)Be�30�3�02�i����'e�d��g敤Y�tIb��Ѳ��0010�v.6N�4�9?%���383=/���(�A��(@�`����	10!���v�` yv ��3!H^{;D�l
 PK
    +Q�HS���   �   
  w/bi.class  �       �       ;�o�>C~F/�0F6�̼�; �\?)Be�30�3�02�i����'e�d��g敤Y�tIb��Ѳ��0010�v.6N�4�9?%���383=/���(�A��(@�`����	10!���v�` yv ��3!H^{;D�l
 PK
    +Q�HА�   �   
  w/bj.class  �       �       ;�o�>C~F/�0F6�̼�; �\?)Be�30�3�02�i����'e�d��g敤Y�tIb��Ѳ��0010�v.6N�4�9?%���383=/���(�A��(@�`����	10!���v�` yv ��3!H^{;D�l
 PK
    +Q�H�ɬ   �   
  w/bk.class  �       �       ;�o�>C~F/�0F6�̼�;F���t���̔,��ʂԔ��̼��"��r��lvfv�*�:�k�9�X$l��r<L� ������DpMu�OIed��L�K,)-JePd`J� P=32�yB�@����%���{#XH��!�L@�����������  PK
    +Q�Hr�o�   �   
  w/bl.class  �       �       ;�o�>C~F/�0F6�̼�; �\?)B�30�3�02�i����'e�d��g敤Y�tIb��Ѳ��0010�v.VN�4�9?%���383=/���(�A��(@�`����	10!���v�` yv ��3!H^{;D�l
 PK
    +Q�HxG4��    
  w/bm.class        �      ���WW��c	EA�kID����Q(��v���!�$��E��z�hmk��.ںKmk�s<�TOw2ȭ�r��f���}�͛%��׍�D���pP���jo��]�򛆣�X$բ(��:Q[�� ��ю؆؎�@`� �nD�����.�^Dbb'�_QA�wɤ>b�e 1��Ԑ�ܡH���v#� �"tEY��c�f�}��z4�SF�t�H�y
iU��@rL?dB�Hx40���P`0i$ꑄa/��E�#�g	EN����Z�~D1��xT��Q=6���)4@Dc�"��(���l�E%s-}�H,œTf��H�90=Ϋ�:��TD��0a���D|�GOE&9ל��6z�:xI�I���T 4f��qO%")c ~��bq8�(�����f�0ry#��d���f2J�e�Ō%�rF��X��2|?��Q˨c�3kk��M�fFcc3c��d�1�2���}����~� c0��GT��jvP��69��®��ר�,���ׂ���q��PQ�5�l%�}Q<\���Ѳ�N����6�^�6�6��sVwM��ȷ����;��e��M��+�n�ږ�m���ӏc��j��ס����N���y��x�/GWݑل�"є2����/ڂ�.�����]_5���v˱iӨ�^��˸�^ר��4ʥl����|tJ#�֨��ը��ר���>�h)}�W�s'���N:I_��E�袗�+�L_3�e|�Bޗ�o�\�8��F0�w��ǒ)=�ڥG'�ZG,f$�Q=��/��?2�S	t���М�tD���_`Y���k���	���W	����F�|����u���7��_������7
�$��f��[�?
��[���ۄ÷�;��N���=�G������G�y�G����£p��1�Kx^ <ׄ������'�E�b�)x��	����§�����	��/~�D���r�O�+�?	��|��#�*�G�w~��g�˅?_!�9���W
~����w8>+��L����6Z~FK�2
�"_IN��]���3t��s�īk�X��Xc���L��M�f&l}��:c%V"1�b$�*�ed����n�O��:�
��?C3C�.\�f���c��E�8�~�r�v5�g��[�+K���Ѕj�H��]��3��_����ǳ�g�U������]��M������JQ\S�-���kt��9s��V�Z��ż�e���޲ٱk�Pp�����f]6;Am�ج;�_g{G�2����f�[���豞��Hl�8C����+����C"�ʭ7
r�~��~�>5�O[��2ǿE��T��:Oa�L�-�D��O/�G.��]�kʹ|��t�B��ȁ�{����
�p<���7��PK
    +Q�H�o��  �  
  w/bn.class  �            uOMK�@}c���Vm�jE� m/�sJQr*� zߘ���	$��'��?�%N�A/Y�켷o�~}|���P����İ�S���Q��@��Kҕ�&z�a��	���b���ך�I�p^E]/�k�	�ZŹ`}���q�p�hN�U�}�e%��,���|�i��S�'��N�ьpQIO�SQ��j�����HB�g�:b�e:#r����&3a�����5f���i��2Q�
q+��E8�[�� g�������F��wq,�ѮԶ�j�ɰ%�����PK
    +Q�H����.    
  w/bo.class        .      uPMK1�g[��Vm�j=����K�ܥ({*� 
�6,�1�ݴş�I���G�o׃���{��7a����	�=B�?��Cm����G�IBǥ��S=_����3��JkE��JY��%�o�����(Bm%͒{u-b�`;@�N8�lZ.6���,	���{��W��`�ǲ�p��+)���3��tT�N�B%L�y7�j���ܜ�7�֪422�TF�=,9ˋ��L�F�Y���1W���J�L��+�V/�b���qQ�#���	�]���-��"XrZ��8��b�׎�>*<3����.���PK
    +Q�H	�7�/    
  w/bp.class        /      uPMK�@�g?bk��~�D�C�e��P��
=���Ǎ]��u#�6ş�I���G�/�t����̛e�����5���`8'�}m���[�IB7N"&z�9��'B��֊ ���Nǖp�����W��L���Z�/j�<��t��p���uf�?�����:��J�a	Fx([��K�Ia��Ą����O�J3U�����&��;��5�V%��i�RB�~�Y��\�:4�����<s����t�$��"k�mv�E8�[�����;�r��/b�%'���c�m�rm+����M�-�w��PK
    +Q�H0�P�#  �  
  w/bq.class  �      #      uP�J�@��&������zm��R����B���ո�ɶ���$x�|(qzh���~fg�����%z�Z0#�GJ+;&xS�D"M	$�̓8S�cP��xx"t�@�u���*�	'U��Ծ���.E��쬂�Ń����� O��!ᴒ��̒��dH�S�������pUi�	�댣�8lb��G�7�L�5o��Y��<�9�w����L�*N��Ɗb\�S5��.��?��3��[q�q�}���
p���{+x�_�.K�Jq��[,��ؔ�A��}�Ml�{��PK
    +Q�H񒶻n  �  
  w/br.class  �      n      �S]S�@=K[����O��~ �H-
�ؙ������v'K�	[�������P�Qߘ�G9��0�E��{oN�=���������i�(8�H2�{^ђ��&|�[-����C(���Cw�q�c��
��+%���(kW00�V�"�%�B2l[{��xƚ�r]���a�h�rm#�Ja���{��-��/�2צ6[��S.��ؕB��|���Ҷ��QyE=Ŋ��Q�v�������]�٫RY^Q������z��L4��J�ҋM��_	h�}���9�q���������e*t��a2��X8�73���0�'X�/��6v�Dr9���`*]h�}�>��T��U���|�m𢭭 #��׀�1өV�8��A\�EXG7":���ER�E�t\RfiC���p�	�pW�e��ps�ⶆ���XP枆q�Rf^�f� �x%:=��Z���ǮQ����{
��)���ώ}D$|���!�����:fh�32c_`��:��XZJi���)2�c�k��������<� �D�7���/L#J��T L�N7�i%��OО+?�F�0O2�4��I*��<�,>I���1s��i$s��I��PK
    +Q�HTy�/�   �   
  w/bs.class  �       �       MM��@��v���\�����!G���eeb��Q�=*v3��ݝ�����Ǌ�n�%!84�1G��Q1jB�ʻ��Wq�ZU�����Ȓ"1��"�X�V�_!)z=�M)���	��s���[;����X��ʱ�93��c���'��PK
    +Q�H�@֨�   �   
  w/bt.class  �       �       MM��0<�/(-�l��D숥[��T�U��.&$>��B8�j�N>�g���o�)	�1�=��PͨY��Jv�\�I�ue	�Cj��ȑ�E�$�	�U�皐��Zel��[�/S;�
>3!wvLY#�Gzƕp�93��C�O�PK
    +Q�H:�,*  �  
  w/bu.class  �      *      }O�J�@=���^��KE��V�R---�}�A��4�����n�w�$���Q�D��,3�3����׷� u��h���TR�n�B�Z��ٲ�"�MGt\Ӷ��
�鞵	���8�XA"�[k<�[�xfy7�N�KE�?��4"�,� 5�A�B��B��������5��N�i�7�%�3Ro��.c�t������?\Z�}o��*r�2*��:n�V�W��r��B��Q*־��ZJ�r�|�&�P��P��g����ȟ<a�1É���������
��؋JL��G(s�l�g��wPK
    +Q�H8�4�h    
  w/bv.class        h      �RKO�@��)� �f�4Mm �@H��Є���}��Y,����'� ����8�"i�v�����f&�_o� �A�@�T��̲I �b�ymz�ct���ҫk=�ڠ�J�j��Q�+�5ݨhu�8��]6����L��j>�'.��@|A�B��:\D1&ȍ�-��Dv�?
�su�\ϧN�7��6D�5�N0�YnSVp�����C���h�����0�m�d��Д�̲��Y�b;D2��������%��,���!��_]����{�{lj؜�ù���H=0�S�w-8�]t�#D����+� ◯p�"q�_!������ iW҄T@��cH���3�IȬ��K�b�PK
    +Q�H����  d  
  w/bw.class  d      �      �SkoA��Շ�V[��Z�
��
T����K�l���H�:��T:[������(�[+r9sνwv9����; ���d��D�e�_��W���m����qԫV�|\3��ɋ�����Ua�n)T��NƱ\�V��:����o��蟛��K�\��{�Q� 5���&�;I�u�����,A�`%	�|	�%�,�:a-�lwf;��fW�j��?��m�6*[���&Rya�ފQp��S���_�Z�-���LL�S���k��QkU���IW]��]�|�����	��_����}��<����^����*���e���1#kv ��Kս�L��H*q�u�P��%e��hb�{'|��(�`��
GҐ�� K`^�x6�ȳ1~y.���Y���+1~�j���i����'��(ץ�P�BQg�/��h0��}8�t�i��aojx<o�MO������	7Q��[(du�V�1��tް�y@GCH�PK
    +Q�H�6�  H  
  w/bx.class  H      �      ���N�@�g9
�YA<`L� ��E�`$$4�pa4�΋�A\[RZ���2��𡌳IM��δ��g'�o�/� ��=�l�M�XR+��IQR�Ʊ���ϥ3��J�r��ʙZ.+"UƙS#@(.�N <�=�$z��G/F�A"B@���(�E!F ղ쎬���ʔs��lǥ��ߊ>Ⱥ՗��*��te1��i�I@���.Q�GyG��S�ꂮy|���7���
��o�nb�g�����us;C��>���GM�I�aG[�t����m6dZ�T9��0�	�nX�SǵM؇%,O�p�w�V�/���3l?	��5�A 2�@
v1�#$�h������y��i �?����	��i`��֪�B�PK
    +Q�H�G�r   �   
  w/by.class  �       r       ;�o�>C.Ff�0F6�̼�;F���t���̔,�����\}�м���<F�r��Jvfv&F.Vv��s~J*�"��@�&9�<A0���Uk;�F� PK
    +Q�H�*���  �  
  w/bz.class  �      �      ��Ko�@�g��I@)}�EH�V֮�U��D��j��׉�nIו�4����? $� ~b�-��m����̷�������; ��@z��!�z��*[oZ�(6��0�fѰ�e0f1gߩ�J�&����">@�nתv�e5�XU<3�R�)�b�T��N� �8|[aԧ~$z��{~N��u��;�%��>2c�Lc\����2j�e!����3\J�Q<�:�����;r���oM�'�������q�.�m���i��~� ����F��t�2��ާH9��KmO�D����57�S~���>�?�R3A�����	䯞��z�Ʒ��S忟5��b���{�΂�g^ת����E�!la�9a�.8��8:b(�A`I�<�X8}��Q�+x���7DY��9�';��~�g���`C�H�6R�/p]BhG΅�ؘ O��%�o �i`9��>6���(�*U��!d`�j��PK
    +Q�H�UY��  �  	  w/c.class  �      �      m�=O�@��'�-o�
J�6���C��qP&7w�b �#��I�@H��'?���I}z�_���<w����ݓ~|��8@�!�6.T��l6���j���Őt["���x0�OX�f�f�f���o��U{t�w��o�����\X�0����GyZO)�H�a�V%�� 26�C�>�I`)+��H�*�
!	�EGB9�&K�h'�ӱ嶴,؏����C�p�PFq��p��9tcB8_7�k/I��&��H��� M�;R`��E�L\
��̈\@�4!�~���vI�R,[J��J�}���O��>����%�������	�T�������[bAI���e�L��C�����ħ§bOŅ-R��b��{���K����{��">�PK
    +Q�H�;�3  �  
  w/ca.class  �      3      mOMKA~^MͲ+�TXf�H
Epw=,�!����.2���:���:���hV��v��y��������3B���Z�v�ֵL�e�mò\Ӱ��0͞��[�ӿk�!���.�x�F����x�d�h��'9��F
k&ag��<�?C	�J�s��ǥdC���mB�������\���|��TA�΀��Gx�w�_sr9e��
��{'�&Z�M�+ȃ�PƑ��Dݰ��H%�P��(zRF�+��<S�U�DjKW���]կ���o8~My��8вӭ�'z�kQz�v���*)�B�PK
    +Q�H��3�r   �   
  w/cb.class  �       r       ;�o�>C.Ff�0F6�̼�;F���t���̔,�����\}�м���<F�r��$vfv&F.Vv��s~J*�"��@�&9�<A0���Uk;�F� PK
    +Q�HP�=.  ?  
  w/cc.class  ?      .      uQ�N1���A�!!ttG+�L	Q�D�@��q.����_�]TH| �X_(\ly����֟_� ��<�2�qL(���C��H�M�I��3."4s<�gm֚PY�$�X�a�%�����j;����Z�Uj3�m�ug��Q:p]�����R|U�2,J�F#�N�T����%��3��"�:'bn�ٷPF��]��|n̔�ԽϴU�h��j�D�Z+�2zI�?�XK��.��2�* �����or��N_O��.��M�����}>� ����`�h��'�9q�cy�Y��PK
    +Q�H4S+WP  �  
  w/cd.class  �      P      uQKO�@�� O�
�'��,��!1xi��h��e��Y,��l�wy2���GgJD�2�~әo�}|~� @�X��c�A�v(8��5��g�g���������TҴ0���C��B�x4�}=�ΣzQz��'"�<ԟ�k�d `kV2�1(����xW�&A�/3�� S��;-���&�f;	̊��VR���l㢮��+���-�����P>w0��H�iX��&���:����G�ȡוc��k��Fj5f�{��&
=8�-l#K#�C�v�3��ޠ�J<�g�=,��[�T��h������`�(��Ocbw.��\���Cʎ!�PK
    +Q�H�4��-  ?  
  w/ce.class  ?      -      uQ�N�0�m����Rn�B/�ت���7�"�ԮR��.NH� >
��PImy����֟_� ��'x�eP��P��GJ+;&�$��,�LE3."4s<�m֚P[�4�Y�a�%�����z;��ݯ��ZLTfs�	]�uo��q6t]����R|]�2*K�F�c�N�\��Y�
Y9�+)R�p"ᖜ}UTZ��	���D<��C�����T�4���Xi��KB�Q%Z�<�q�=��U9�.G�|���p��x�/�tgn�8F��6��ihD� �?�.��ˣ͂�PK
    +Q�H�k�\�  �  
  w/cf.class  �      �      ��QO�P��es�
��PQu�4��ۀl!���,�@ܛ�]��-�:���Ʉ>��pNKƬe�&�۞�=�s����� 9��V3�6��b��+��74�<,h�|��Uu��t}G7z����LW������Q�W��V�)4B~�Q4"<���a��z]ny�s��n���Y}W�P1H]���a�r�k�F2E� I��H�I�i�I����]i�oK��^�A���i�u�<,��k�P�Yʍ��]�|�+��ڊK�îŰ�֐[?����*t��#�~��m�ehz4��ԙ��'T�׾	O�d��4����+~���������A�f���9�����@���i˾�z����_��� s*�J�ρuX�mte�Q�����+�����?)��?��|�Ɇ���Y��1f��8 VG��(����&
<�;��(0X����(����1��Q��I�����I,޾Z�]+��)Ȇ7�PK
    +Q�H���   -  
  w/cg.class  -      �       m��J�@��4M��ZA�\�0d�Q�d�@�+���4ԑ6)m���Jp��P�m��{��s9������c��j�p�i�ű˥+c�8R�8�C.D,�L���u�K]���^�����W>�7*��wE�D�D���h�.�ov>ݝg-CoP-��x�'/v�X�y5����p�p�O֧���}t�LV��=��Zϋ�^��Hʲ�G���αG�f���#�N�0�?p��tIO�@���B;��PK
    +Q�HC��-�  Z  
  w/ch.class  Z      �      ���N�@���殸���f�,J &!i���RqNM)��<^�x��P�3E6u���9����߿�yy}z�llm�n���3�A�@�*�v�R�bI)�IMQ�=U+�m_%�s��C�K�d�T($��^����t�Ó��U�2��	�nX����[j�w�� fوl=�d��-����Xv��l^��LZ��f��X�b\_Sú��ʩ~��z�C�]ej�K:��pL;'̮���\�F�L4��d]z����E_�[Z��f�?�}��K�������NJ��O����I�G���!-�Bz�aVq��VG1v��2���kMS�r��-�"�w��9mۄ��c��"]���)�+����kR'"0���gX�u\���a�>�����]K^`�0,~+^ �@�+���� �{�q7��0�5�v3r�!�unoPK
    +Q�H.�[;  �  
  w/ci.class  �      ;      }P[KQ��5/]�J�=h��E�
>D��G]�c�Y�*�������h֠,$g��.3̼���2H�+�2��]9m۩wm��8�U�uږ-Dת^V�Bԯ�2M�ʴ0��D�>�j4��������z��sD�ԂU�FBX2Y�`p��1KD�W��d���|�ub*��V+4^�X�[�h�렱�KH��x2^�E�YO�O��[�$�P�m��#Z��.B�&^_�� �n��Fi�1��+��BN�H������=�J�����>�<�C�6	�H��S.�h�~օ�R���h+�f��PK
    +Q�H"���9  �  
  w/cj.class  �      9      mP�jA��y?L��TX&!�uQ��(,x�����:+�h�g��!��
�1v��������?>��!Y�x[1���^��9�Us�U�ݺ�p��թ���}���m�LK*��LP���}����i��`�Hd��E��4�Gr:�B)>��^���י,�|.��=�S)�XO�Tڏ�1�d�m�b#x Ԍw^��l�t�b�j����y��f�S���y��\�#����w�
��2T+��PΔ����5��͜�y��n�Č8]}�ٛ�m��Jf[8�q�B�TY�m�t�3
dd��td��?PK
    +Q�H���B  $  
  w/ck.class  $      B      u�[KA���̼t/�ނ\a�(¦-,�I���,�댬���z
z�����Fvac�9��������+ T �/jC�ݶ��� \�f�\�z�֨�u�j�7�kC7n�]Ӭ4��r��9l�ɔ�6Vsf=ʙTk��Xq7�v�l<��g>��D����0�����m�V��V��\�t���m��Y��]�l4-j��A�O�W��\:̢�Cl'� �Ӭ,� Ӑ��EWMh%��@�bn�R�\ېR��J.R�H��������a�B猪�M�(=��S�#Y�!9*b�S����k��8������~�ZB�PK
    +Q�HD)�L]  �  
  w/cl.class  �      ]      �QMO�@��|ȇ���L<��)�@H�\�x0�h�j�%e+�˓��?�8�DlL�d�d�y�;���� u8%��U;�!��j�C�K=�}�y�j�M��jԴ���k�f��̚a���aXV� qp�T�?�G>�<���\�n߳GƗ�@���{,���`w�@$�$(�)�JA�@����aLR_���ɬ��d
ju���	��|Q�H�w^Ft���^�顝a���Oo��8�2�G8�Op:�ۀ	:s�tAG��g�GP��wt��.�A��J�.�<�1���(?K��wB'r�P�c�Y��Nې�j�ȅ���F"���N(8\	����5��Z@�PK
    +Q�H	P6  �	  
  w/cm.class  �	            ��mSQ��#(����K�Y!J�H�J&��e��e/���b�hN�/�46Ӈ~@?��~�Φ��ᾁ���9g��9��_��8mrxG�'��@l20��!0	�#�Q0��-D��������kƌ �B)}�&���A�=�A[�6��v �	���3J*�mn)���FnG����z���(�AT��U��t �y�l���%>B���	�*6��������V��f�c�gk`kdkbkfkakekckg�`�d�b�f�a����������E\tQP{�r�K9M7��iA�'����$��QP�R^�x��+iŏsT-u_U���Q⸐Av�L��qI��#�1m���?;|A:K~���5כ�W�g�fD�~B6ö<���LOY�C#��B�o�����U�w���O���	������ߗ|3�.ݟ/����z���j(�@N��o��b��E7�Q��f�YE�9���_��&N4�rA7��tR��R�tD�s�jh9'�{E��QȧiE�|��	���'|
>�|�h�s!x
��$�eR��C(��i�Ye�je`�-W �d�*@�\h�/@�� 4ɀ�YF���X��h�U�Ze�:@�( �2p�S��d  �- =2���M�^�e>��˱d��U���I󭩴|bL!pIV90(a�.�[޳����50cn�J����]��xuᯃ��7��^�ѫ��V+?6��J�nl>'7+f�G��d��N�v��Ը����u1^��y��9~PK
    +Q�H��,\  �  
  w/cn.class  �      \      �QKO�@��)� �f�5͢Ph!��&�F�4�bْ�B��O&��(�l��1l�3��������	 7P$-]A�(Wջ��W���J���)���S4��ukU����M.��"@�3ǵ����	�ft�L��$����f�&�ؒ�D[�D�HI�!P��:0!耻����_d�m�ɗ֠{��tr���ٟ��65�`!���a6ە��5�ٿ�;/���[!����~�,� ��,�{w�1>{����>�C�l�x�㎘H=rK0�wM8�]��"]0���L0ǯ���M���p*���9��=�IRA�6�t ���MBfM�/Ks�� PK
    +Q�H��v�P  =  
  w/co.class  =      P      ��]KA�ϸ���wiV7Aj,�n���&,xޏ���:k���
�����3J`"5�9g�}�9����� TႀV,	$Z\p�&p���6�������~sg4�NǬ�]�RG��3M� c�����y�����_�@�+@%�RL%-	�$�	�A��Q��	eB�!eļ�og<�b�ZV�\qź��N�,Y
�V�����������pi�E:�%z�j��╊�BH� ���6>��	�}g�g|�9��d�bF ��]�d:p	�xL�8�gw���78}U>��p�ȹ�>���B
ݶ �@|8Y�$�갃@r8^v��H�J���PK
    +Q�H�$��  N  
  w/cp.class  N      �      ���N�@�gA@�ꅉ�i
!Җ�&D�F�h�BْR >�W&^� >�q�*")�fg����f�o�/� ��C�T�A�8�jYE+�%EՊRA������*ժ��U���ڹF Xf�9��hHZvGnڬݕ[��ܲ����{ܚp�15G��	�~,"|"�C�2�x�ǆr.7�패Y��L�PR��vk1�v)�8�T�锇����r.׻tLe��<:F��U����o�^��^��n<N�"=�6��˗��"G�_G�#ư�$+���V�6�=q7��6dMӨrn9�a߳���6�Vq�x@��I��pW��<C�I��1�����EhGH��lM��y �@`��Q�as
l�1��S�"5�PK
    +Q�H�I�{    
  w/cq.class        {      ��[KA�ϸ^���.�=���1/(º���C���"#:k���z
z����3k��-��0��;���y�x}�+8!�e�MO���^Ε�Y��(e9����FV/6
��Q*��"�p�.����cM�`bΨ5��G���$�DST�@41���h���>eB�6w��?k4��3���D'�Y�n.��VՇ\��V�M0ѣ&&z��=����)U~�;�'�?C����ߪ/��o<I�hF�7 A� 	�����N��&B���c�غ�d�;bL z�{�ɉk�)lb�z"@T�C�%1���8xV>�}��j���#�q���G � �.	�C��[V=@�]2ּ�>�:?cc!��Rc�>PK
    +Q�H4��C�    
  w/cr.class        �      ��[KA��xɼt��f+�A��Eؼ������nˈ�ʺ*}���� }��Fl����93;�߹,g>��? �W��l�@ �e57���
m��o�wżR,T���m+�4ԖR��7J���ܩ MG3О	�l4�}`A��j��X	�#����KA$QɎe��o���2!h��Ό��}2��5���D%�qI��aW�d��lڃ�ut��֗@��9�#&L����z@�U���
���ʭ�i�?�t�݉ws2k@"�3�T���RO3����S����n�)�p���93ۀk8�0�l�Y����r̽����	^8\��CҸF:DkC �Yv�B�72��"r����.�d�wU=�GS�PK
    +Q�HM��7�  �  
  w/cs.class  �      �      ���N�@�g�POx�#/@CVQ1AZ�&���/АEܚ�h|,�L��|(�l	�M��f������m���� 2�C@I�j"E.�{F`W?�j�J��Ν�szFO�d��R)�׵�^�*Gèc40�V,�E�6o�i���6�;j܈[a=
���Fi�Q�1�Dd
ɤ�4"SX�Q�	ī_�LZ��e��we��Ф�4��K�״)��b�! �m��h��=r�������B��
���&�����f��+�R�+���Uu��n�o8! �������1X��
�ߙ5��z�,	a���p�]�`n�6af�L*��&>ż;����x�:AkXFd[N�c)@�9�1��8 ����,�U?0�@x�a�L!���4��3x�/��%�OPK
    +Q�H�=ȁq  �  
  w/ct.class  �      q      �Q]KA=�_i�_�}���l����*�BQ�S/�Ȉ��:V����~@?*��&�ý�{Ϲ�����|{P�!C$�o1DsN�a8>3��U,J�U(7땂]��
W�m�e��>7+�K!��10NѦp):�G�y$�d��ɦ"���Ns:Et�&�J`�!s�]��N��R-��W#�Ã���q���sSЍ/��>�ipy����s�5*t�[�OrN���f�tHI��&�a����o�ED�RX���wh��ۑTb��P���-����2$�DWr5
<a����*���km��N^���qƐ��p��i�Ӿ@����E"đ�!dg	KD��f��qg�B�����,au�gS���|PK
    +Q�H�X�R  S  
  w/cu.class  S      R      }�]O�0�O�K>�V�2�4K������.�&ܗ�,%�#���啉� ��B�d�����}�Ӵ�����\HT�C�6\v\[�n�z�N{|����m��kZZìY�u��h��a8c��#�@�:�U��>���v3��(�У���'�	A�<��[�g6�N0���UJ��О.���6�b��6Fh&l��τGm,x�v���A;��'hZ�걛��*���A��
�xk��HH>u�|�G�k
H&y ��/�LF�W��6�$��.����h9HݼC�M��#r��8�2�<Br$ѷN��<�g�@Ӻt�JsH� PK
    +Q�H��^�Z  �  
  w/cv.class  �      Z      �S[oA=SZn�jk+��KkU@�ݕ��@���MxP�$>.���t��K���/��&���MZ�f[+V�n��w�|gfg��~�@�E�!�δ��v�fXHہ����s9KъE]�n*ռa(�Z����s�KX=W3�UK1M�S���+f^3�V���U*�	fh�z��x�XE���:o(ŒNؚer�`�R�!Z�]�����y�Hshthti�ֽ�@��ޞ�=8P�޾j��w,hG�pܧ�ݣ���C���4?�9���	K��z��0$��!Զ;��ΰ̐j���j��Z��U��J�)�S��n�9G�:t�@m�#W��سi{j�K�~T�1%?�+�8WC_���,�)�6M�;��B��ʒdz?S�թ����g�fKZ�M`��aN��2ݎa�H�Q��txL���zt��,O����g�+�z,|w��v�ΰ_���%C����G}lSJ^6�ԑ�����sX�|i*_���T~a�I&Y�f��3��d?R ƈx� Z��T�ڤq�ƭ �}عH�%�
�!�睓�@�,�ٍMF�g<� �#J�oy� ,}���v����	d�ӯ�?���_PK
    +Q�H�a�E    
  w/cw.class        E      uP�N1=�)�B����d2�Lp&2�I��� R��3�]�L\�~���"�6���9��~}|��B��j��Fk� �f���+��s,׶��n��M�j��4�c�M�6M�yC@<��&�0`�gc4�#13��b�	ү�4�e��1Z&�P����"��A��[���� ��i�/��M]�T5J��|/���\�5���"k���D������1��ɣ�c��ci�����[����r.B/d�/r�l½0
|\`W��H��*r�ʬ����;N�Nd�p��T�p�����'W�"2� �1PZ)�6	�5;�Z �PK
    +Q�H=#��6  �  
  w/cx.class  �      6      m�]KQ�ߣ��ч}(]]h�C�Cpw����Y��~X����~@?*�U/�̙�}f�����p�:C�ќ0\�wf�m�L�g���G�64:�fu[�ν��{�.C�A*�C1cȭ���{/�Yl�k�F#}X���� ��4��9J��D�����\r'Xp۶ȩ5���@���M��f��0����P�I�����Nz�D�GԓvUh{VB't��辋�D�r�Nd$��;T*�E,1���D��..Q����lgTU�? w��ӷ�g4GȠFE�8�\&�"o�H@n��J�~��T���PK
    +Q�H��GN�  ?  
  w/cy.class  ?      �      �R]KA=cb�g���F���CT�cJҀ���CQ��$Y�h�������S���Q�gV�[�Ҳ�;s�={�;?~~����Ta�%�ih�mS`�Z��V˧��^m�X9�����i�x��R;���Y��6�!��/��=�u�Jvnoe'��ޥ�6���ߩ����Hv�S4 �c.�\H�0�B.��,f��~wU�Ȗ�P��V��yǬ,b�ρ6��[t]H(4ήԝ�}ez�����f$����c�Ƕ�OI���_��g,�cc��д�����M���AL��q#GA���=
��*c[�ʟ��7~Kt��Xe5E��g��>��m�q�4V�J�<�9�l�ϓO���d����t��3�эs�����~V(Y�~xK+�4E�Ĵ��H��I�.�Q��	���x<��\j��/PK
    +Q�H/
��B    
  w/cz.class        B      uPKO�@�D����x M�" 
�p0�/�4�eKJ���ă?�e�ֈ��afv��Lf��_^�c����K�[m��F����]]���U�ө��W�ZU��6�RI���É�Z|���f3>r�ܸS��Y*��Bؾɰ���(-C�X�8����Y(���|a7~3��F7`���ڑ�3�F�`���!.���D,����A�E�V�.�[�\�Qd
li:�%��>�q�t��<95r.���V��'5gH�JK	�wM�"E�ϯaa0R�	_@��O�h4vA���pD5E�4Ŧ��P��d�
T��� �#�PK
    +Q�H�s�=  �  	  w/d.class  �      =      �TmSU~6��7�Ra)-�J�/$
֗����I��baI��ⲛ�nx��T��ݏ����'�Τ���K���f2錙�Ϟ�g�9������?��,�!ܹ+��o1a8���	�~�'�dx��i��A����0��p��u�� �\�6�Ćm��42�B��8�s�_�J�q��W�c)N����ɜiX�wF@��1�9��%@:���TvF�@�Hư�[�䢖��lI��1)k��c��Ȗ��,1���7�	]����ii�W+�;yrViQ��:�e�$�H]u�VA@{A����;�61EJLy��Y�+����ݤa'��򲞣k�{��Y�乭�^��ڮl���N%;p��kz�;@Q>�����T�0�M�g�]O���:�h42�v��N[e��ѩ.�%ޫ����%S�Q8�L�b��i��.�:�Wݠ�n�l%4'WL�5OK��yݤ���ף���s4,�8BDa	/JxI�i	&%�,ጄz2-�9A|,�<�	~�ǆ2̓!�����C�T����jK~�!<54ЊoUp���j+���J�	�8��-���z�ᘂ�+Hrx�*xW���`�(x�ı̣S����<4�aU�9�#�e\�b��Kpe�G��(ʘǻL���\��u�2�*˔����ơD_�i:[:�m����kfY�=-R%@�q��$}����G���6�o��h�g�O6�s�5�oB�C$�Q��K�o��'�E��>��������S���⃟!�wq(.�n�:��U|�>Rŧ�ᶱnG8v��W���T�ĺ*�T2���'����N�V�U�X�wtid덌`)h���c�T1}ۿ�FO��Eh���5��P��.���M�IEy=�0�د�k��Q��_�D}�@�	t�@
��mߛPb_�Q���U�}ձ e�"w�dc-*wS]�P��$������AG_�/��h������q�U�ɏ��+q5J�����s"q�!�}/��\q�oJdʾ�*!�j�_Рj=y�H�>���fx|?�l@��߱��PK
    +Q�H4hd  H  
  w/da.class  H      d      �PKO�@�ߊ"�L<�IS�v���`[�&�F��
[R�D��'� �q
F�q1�ٝ���������<C���fHօa��i�kVI1xQS��4+W,�j��2/VlN�3ӲOˆ��z�\�x�T�v�RLM�%�ȍ���\�Á��N z7jw4R��Pu�����a��L<��T�qz����J!͐k}�])ն;�1�[�ۚ�+Ǫ}w}^9c��g������Vp�?��_�T������{��"��*��w�������c�xM)���/��+їn8	<b�l�I���=��f�t��ǈg4^�cا"���\!�:Ų�	��ퟂ(��,�4F��$�PK
    +Q�H���O    
  w/db.class        O      m�KK�@�gM߭����^U��h-��U� 
�o�����l���$x������J�?��fgf���� L8!�5��N�ݶ�N�30u���9��Ƶ�ƕa���6�z\p�'@��As	4�ȧӈ�3�,�	���x���L �dA�ȼPw�aPB�l(є�P�C�@m�[�	A'<�	��O{�H�^c!ҋ���i�7��%�>�1�cr�+���T���Cg�?&B�7�1��%D(�䡈	��/�L"Na��������VEO�g/���Uq��X��RF��V��� �6���֪��j�M����mL(���Y�P�7PK
    +Q�HWYOe�   �   
  w/dc.class  �       �       ;�o�>C>Ff�0FS3G3'3]G]CCgW]'cG]#G7'GssF6�̼�;F���t���̔,�����\}O���Ē�FֲĜ�TF�r��dvv6Fq,z<]�y�������S��$�J�J2sS�2�3�rR���KK2��8�JA���$�'f10�jmg��U�$��4'�30 PK
    +Q�H1$�K4  W  
  w/dd.class  W      4      u��J�@��m��<�Ck=�xE�eKA���Bz�%!l�H7�����|(q&����f�of������+,��/t"`�w\�FJ+3�bJRDՅLr����?)�hXK��b�Y��� �bo��p�I����L.�!9���ݧJ�(�3:�㲬e��Bz�Ա��AL���%sF����.��pW6*���p�����C��z�&j��It�uj�Q���U��ɳgإ6��BzBU����]����}A/O�hRާ��h�Q+36�뿱UtW����6:��*�C���[��7PK
    +Q�H�k��  �  
  w/de.class  �      �      ���N1�OD�}�T2��AM�dL�F�LH;:�+/| �xN5�X���?i��?�}}{~�$�	[i�A0n�`~s����ٵ��u��L��GɌ��Csʹ�͌��m2h�R��*`�JX�Q�+O�.��͍Qt��B^I�^2��J��Qr� a$-$� I���$L�F!�����H:H:I����C����F^x~�W�?���ه�ƿY������H:�vR����Wo�
����K~Ǎ
�e#��;��ȯ�7���G�D��/�se�A	;!h��$���n	os�&}q��EU*�%��s_��� r.ʒ�5ρ��}=�����ѕ/?A�|�ofX���Bw��4V̆NP���R��Wr��F ��Q��u�j�m��ѦK��V�� ]bP��$�T���,6�*Y����5G�f4k���M�j\%� ߚ��T��PK
    +Q�Hzoz*  9  
  w/df.class  9      *      �P�JQ][S��Ů���B���eD(#���8�����O�sz
z���h��P�=�a��Z{?��Ϸw �8 dk�.��,��Ӥ����Ҹ�$�J+�"��t���c��6n?mOY~��P��	�� 'T�PH�EW�&�����Ǣ��m�0sW�F�J/���m����T83���&���
j('R�R���x+D��F��u���P	TٲvಁG�6j�uU�߻�:0Ҩ@G��hi���1�|�L�$��V�O@�񊝗�'~�-d��K���^f�g�F���%nh3�"d� PK
    +Q�H;2$d  �  
  w/dg.class  �            mNMK1}�ڮ�j���7��V�� ^��^z���n'e�m�gy<��Qb�R?�2o2��d>>����O(��>���jv�/Cw�-qqI(�+�!�#�Xg�d*��d"�z,�~b=gBi&�<&��E��g�P��{?}�Y�Ufr����U�_ҭVl�,h����ə��D\?�8�XkE�*�ٝ�:����l�8���6�(�SB�^%,M��8�ks(��{��U_d@��;/N';[ֶ�0oc��5�[�niU����/PK
    +Q�H�Tө?  I  
  w/dh.class  I      ?      }�]KA��㪛}�fEtaE�B�a7^D���.��:+�����.�����Za"������9�����@��z�$�%��L�k7�&Ϥ��5��kB����Z��z��T��KH?��7KO7�2�2b�X��#�;A�^�C!�]F����x,��H8�;��u(�a�<���p�s��iv�r*�/�'>�n%u����+�8���E���ceA;�@*���������A$#�	!��<-�8tq�u�f"2UX+���L���{/�'J�>o
�7x���7̴��`�(-E�sv�չ��a��PK
    +Q�H�p\�	  M  
  w/di.class  M      	      ��mOA�g�-E�`QA�ϻ���k��^�}���yY({x�B�X�2��e�YH{^� ���nw~3;;�����/ h��L��h�0X}�e�l��6�>xc4�wF�ڴ�ڰ��V��޶���j��H�Ѻh.���}A,�Q`v#���ٙ醧��I���B2ȝ�� ����$�d�$C�%ɑ�I
$�$E��I�d�@������\J�#"5�濞aI�z�j1ׇPH�GMjM-űwx�Ϲ��20[ߔ�����������i'�)b153v��U�q�rl��1��1����0jw\���p�Ϸ>��{^�,L�`^�صC�o�ʾ�Ru.��z4�J���ݞoK*�B�E �D>,���I�*�!L���u!���~㩨�q��oF#����4��'x�@C��E3��S�;�"P����6ḫ+��z��S��I�>�1�ex�@1�&�9J1�Y�G`�"P��$P�E����5S�HG�8�k�8�Ķ�i���PK
    +Q�H���[U  �  
  w/dj.class  �      U      ��KO�@�g@@�Do&��i�4�А��	1�74�X���\�L<��P�)F|�&^<�������l���� T(#�+U�X��uCQ�F��H�j�KM�D�Šj��ij*BV炇md��?��>���t*��l݈{��Bf���AX���q��A|a29�!���b&�ls?�����Y�ZgԩV��.=.B�o%����G��m�\�ٌ�.#ټc>�t;�BO��m�,����?�G��O-�� ئ��ސ�sЋD�'���wC/d!�D����#���w��${�!.�.e[�@��;q�6 ���أX$�D'k��X_�?�<���Z\
 �PK
    +Q�HS��Or   �   
  w/dk.class  �       r       ;�o�>C.Ff�0F6�̼�;F���t���̔,�����\}�м���<F�r��lvfv&F.Vv��s~J*�"��@�&9�<A0���Uk;�F� PK
    +Q�Ht�T�  �  
  w/dl.class  �      �      }R�n�0>.P�����2�֭]/�RC� �B���H\T�ƽ��K�.�V{�^M�E�5��L�1o�|l����~��� �pL U,�	��~�'p�ݳ
c�*�Y�:e^תWZ�V\�}֩z�#�z.�H�������Fk(�8V�ѶE�Ki�:��S%@8��!�B��A,F�����F7��I~�ѽ$����4�v��Q��A�
)�*dTX��z6	�z�]��v_�ɔ������ޕ�i��������t	�qCP��+���,�d�(q`2��|i45�1̚ 53ՅQu��r9�}L������E^�kh�-HـW��ˋFxm�˩L�M�1���Q��	��+1�<���.�ԷD�����»=�N��
&�p�����4����i��e�3$d�Gx�	����\y�L�F�ڂ��ev��	�e��_Uw�W�	d 7[�~PK
    +Q�H���B  �  
  w/dm.class  �      B      m�]KA�ߣ������M]����.*�����Ey?�"c묬�J?����~@?*�U��8s��9gx����@iB8����F�R0�v�4��^��Z3��k�R�X���N�l�5!�W''\8��]1��t�΄���I:I�̹�[��N��1��!FHw����'\��v���^k�%����9Bz�[͚����H�MR�;�s�l.G���Y��
��+�5S�%���2v����{_zbb��L�m�!��qO8rF�?����Z�BR�����A8V���Dr�8z	tR���NUR���I�TDMl/��5�������	Z3�� PK
    +Q�Hy���   �   
  w/dn.class  �       �       m�AQ��5�`PVb�,Pz�lHil��b�����~�����(yf�9���s���� �A�`�B��i}���X�!5�,�!����:Jw+և�X����y�����O!y.[HZHJ�?�ɸ����BV��^yv�P���F�*\�Rq�*�:��1"��W�`6o���@^��7���xPK
    +Q�HB1W��   �   
  w/do.class  �       �       ;�o�>C>Ff�0F6�̼�;FgC7G]c7]C�c]K7']3cKWcsF���t���̔,�����\}�м���<FֲĜ�TF�r��|vv6FIL-�>��.�<L�\�\@-��)@��A�y%���a�řI9��yy�%�%��y��@� ��L`���X��3po�*���@��Y��PK
    +Q�H��e�   �   
  w/dp.class  �       �       ;�o�>C>Ff�0F3''cC]SC]C�]'c']GgKCCgW3F6�̼�;F���t���̔,�����\}�м���<FֲĜ�TF�r��vv6FIL-�>��.�<��\�\@-��)@��A�y%���a�řI9��yy�%�%��y��@� ���`���X��3po�*���@��Y�� PK
    +Q�H��Jv    
  w/dq.class        v      }R�JA��6I\cL��-�a�9! � /�&�1v�=8�����(�:"�6�j��-ݯ����@U�x�|-�jH%uS@��&:�O�-�%�)0��=�﩮{��-P��ێ��s�t4��/#��������C��aH��JJJr��8�u0/�o}����ATgϿ��J�F��)�ʠ�s=��&F&�d)hFQ�7�����,��j�>�z�9ӈA��b��8����V.�J���Zd�+jO�P2W��<=��`�i@��6�̿)�1w�%i3()N����86c���J�֣H�b�G�����%ʔ��2e���3�	J�r�/>���O�aM���E6�Q��j��c}�|V�> PK
    +Q�H;}��P  M  
  w/dr.class  M      P      mQ]KA=������k�Ioj�ϊ A`,	��4�.2���:k��z������na�܏���93w>>_�tq��o�'ž�B's*��v��ܾs�L1Xa4��Hx{��x�~Ɗ��Px��(O�ЎH3a�(��b�9��PH�G=���*��FΨ�?�^tHiII�?]���|D�9)je`{�����������r�C���r`�Ye��H�&M�:�h`͇X*��O�R��?�2T\�P.Jc1�\ő�K��1h&�l���)��#�(P!�y;L ʾeTu2��s�G�)��I�5�_��v�L�-��Q,w��o�]�$ŤJ�PK
    +Q�H�����  �  
  w/ds.class  �      �      mR�n�@�m.n�@��B�M�-��;$����"5(/<9�6���l���P| ����>�̎���x���@m�R�ZO ۖJ�m�Kt	���'�o	I�Gޱ熞�{�Q0�|���CB�@1��n?���}N~)�6{���d��m?"޳������̱Nx|���Sl���9C)CiCCYC��yC9Cy���X��N��r_� �[�jg�-qp���ǣ�U3�V�^ER� n���l����Lk���v�c�Dk�{
( ]��p7��vw��nu4��tv"�C:�������Zi��<zr,�a�L�H{Z�H וC��I�6�XB	Y�鞘��2������	�A�K�
}>�7�~����?�_�6��.b�`�r�lP���T(K�`��l{���-�BY�W)����-�N)ق�0���Q�kA-�O�,���篸��\�i�-����t�Ro�~�z�G��[ә��PK
    +Q�H����v    
  w/dt.class        v      m�[KA���*���|�C�x��P$t���n6f������J���������x�wv�of盝���W"�ұ�p�t%(V�J� ф�u!���B�����cճ�;}����NP�zv'�n�n�`���0:v#�y�]��M����l�([��b��%ؒ�Z��h^P���!G)�Lz��^ZX��|�WŅ/���w[2����v��UCm��2�Xk`N�B$����Il�h��w�{�r������PvމR�v���PP�-{�ѣ�ï��4�a&�IP��i�6i5�ED�r��	,!&��H�@����`�6�UČ	�!�L`��w*Ae��t�;S�P�o��B���g�oN�~��	�>k����>�PK
    +Q�Hn�`rV  l  
  w/du.class  l      V      mQ[KA=�m�n���]�����s"�B���O��f#6��[�'!�Џ��Y�v��wΜ�|~�} h�!^�R-!�n30N1b�N���S.���h�9��諱=R�}�G��9�Cba�A��aKb�^,$-�,l1�{k�;_H�K��ƔKiw����+�M]�����z�w�⎑n�E^��C��/2�Ԣ�a�-!��m5z�~ѵ��b`&3�ÑIe2���c�>�Z<y1��ב��\_��}1�\�������z��8�Z���i�L3��6u��aH6�r&�3�pBP.�d}����C\�0p���Q���w�.QYqV�%�PK
    +Q�H�o+n�     
  w/dv.class        �       E��Ja���Uw]�R���.4X�_�E	�%��.��MEVd�X�����衢ٌ��93������9s�V�?S�kc��@����0��o&:���"-��H��4K�kEu�ۨD�\'�$�$�*�{\/繢���llǦ&�iA�����t�?��jԟyTixT(�F�c���GK��O���^�b_��������T���='/�P���X?\�����>��PK
    +Q�H1�Ձ!  �	  
  w/dw.class  �	      !      �U]we~����v[�h��6Ͷ,��B�gj
H5ԏn�%ݺݔͦA?.��F�r��hREQo����q&ْ��s�9y��g杙wf��?���!�=�T��@Q�A�P�Q�&	� �JD��</!��%�O���(�2�$] ���ږcy#�þ�9�,����8�<��w/B�����`z����lo�*D����&�'Z����9z�3��X\4��f�?K�y�hؤQr��)sFa�H>kJh�7���m8�8+%l�ǖg�E��;v�ؤm�9�N����xuF�uF�g�LW��q�g��Y�)j�s-''�k-5Z��lmѳ�x�u�+|D�tr��˻���ke��g�E$��G����jTe�p&�%Au�Eۘ5�M,��-<)Ns�8S��j��'���,/?QS��B�G��,D])�*W��i.ǳ�4D��2��񬌈��d�񼌝2v���1H�O�;�MHk8N���ig��88	�ֻN=�����[˓�hjm�x�7E덫�����l�wF��O��Y~�:�I~;�c}G;��쪋�І[z�cN�������T��o�ё�Q�̓�=|�ƣM-����?Q�4l�f[1���4��fP5���%��UC7�4���Hj��Љ1/�UH�ݸ�>��Ѕ���gY1�a�b8ߌ&^gȨx�*ࢊW�eȩ���aA�AL1��`0�*F�Cx�a��b�Wq����b��@�a�z�m=[t<k�<o��L8N�3�����9�WtM�$���PiH����^h�'$7�8>������ٓ�^aa
����d�'�Gd���be|p�r7���W�hM��e��T��_��d:�e��ƾG�Zc��o���<z	7&k��}oW����\L���2n�����T�`�_��7�g�����J�,�
��Vp�������;�������̔q�#T�5�z��������=
�N�9��~"g�0�H�,5�~�PV����n�ԉm����[	�Sz`����-�z�*��i=T�1�<}ׯ@7N�Ά�U�ָ���]=�5B����H|��~�q�7$�������&�w�#�aG�p�q��wSOv��ÃeܦJL����ur����)�N-�W�N/�k�2�������Wu�ԭ��3WKX��r�&~M�c�'���n.�

��%�_b�jc�䥿��;�W](���	^����DƟ��Xd)�3�P:
�3�@:#+�"�3",eAz�bE�h&T�J�"Z5���V�6�F�AlH߇S��PK
    +Q�Hˢȩ�   �   
  w/dx.class  �       �       ;�o�>C~F/�0F6�̼�;F���t���̔,��ʂԔ��̼��"��r��
vfv�*�:�k�9�X$l��r<L� ������DpMu�OIed��L�K,)-JePd`J� P=32�yB�@����%���{#XH��!�L@�����������  PK
    +Q�H�K�b�   �   
  w/dy.class  �       �       ;�o�>C~F/�0F6�̼�; �\?�BU�30�3�02�i����'e�d��g敤Y�tIb��Ѳ��0010�v.VN�4�9?%���383=/���(�A��(@�`����	10!���v�` yv ��3!H^{;D�l
 PK
    +Q�H����   �   
  w/dz.class  �       �       ;�o�>C~F/�0F6�̼�; �\?�BU�30�3�02�i����'e�d��g敤Y�tIb��Ѳ��0010�v.VN�4�9?%���383=/���(�A��(@�`����	10!���v�` yv ��3!H^{;D�l
 PK
    +Q�H�,���   *  	  w/e.class  *      �       ;�o�>C!Ff�0F6�̼�;F�DF��ĲD��ļt}Ϝ���Ĝ��ĒT׊�Ԃ���<F�
������9����,���l��>5�%E�y�� �Ա����T�����"���x�8xX��SR��N)z�(L@37� �l& ͧ}��g7{��v���*����h0�  ��X�@��� PK
    +Q�H�+��   �   
  w/ea.class  �       �       ;�o�>C~F/�0F6�̼�; �\?�L�&�30�3�02�i����'e�d��g敤Y�tIb��Ѳ��0010�v.VN�4�9?%���383=/���(�A��(@�`����	10!���v�` yv ��3!H^{;D�l
 PK
    +Q�H�;2�   �   
  w/eb.class  �       �       ;�o�>C~F/�0F6�̼�; �\?�L�&�30�3�02�i����'e�d��g敤Y�tIb��Ѳ��0010�v.VN�4�9?%���383=/���(�A��(@�`����	10!���v�` yv ��3!H^{;D�l
 PK
    +Q�H�w�   �   
  w/ec.class  �       �       ;�o�>C~F/�0F6�̼�; �\?�L�&�30�3�02�i����'e�d��g敤Y�tIb��Ѳ��0010�v.VN�4�9?%���383=/���(�A��(@�`����	10!���v�` yv ��3!H^{;D�l
 PK
    +Q�H�]�   �   
  w/ed.class  �       �       ;�o�>C~F/�0F6�̼�; �\?�L���30�3�02�i����'e�d��g敤Y�tIb��Ѳ��0010�v.VN�4�9?%���383=/���(�A��(@�`����	10!���v�` yv ��3!H^{;D�l
 PK
    +Q�H��&��   �   
  w/ee.class  �       �       ;�o�>C~F/�0F6�̼�; �\?�L���30�3�02�i����'e�d��g敤Y�tIb��Ѳ��0010�v.VN�4�9?%���383=/���(�A��(@�`����	10!���v�` yv ��3!H^{;D�l
 PK
    +Q�H��7C  A  
  w/ef.class  A      C      mQMK�@}۴��P[����[?�疂B!�X��ӦY˖��tS�gy*��Q�lD��7˛ٙ�}�xy�G��jw�šTR�ؘ�	>aF����+�\��k!f������2X�'3�mV<L�&��{��3�3d��(�(ۨ24����R�a0���G7x��i�ʸ���"��;YƝ�w�4���;�y�[FTSE��A�84tDk]Fm׼M��b*��ŅR��ZFj�P�ȹ�:�Zأ2� ���`8�S��A���IR�2�H�Y�6��Q#��2�f��d�ӈ��q�l~(��	�v�k����Y��Y��+��� ��'PK
    +Q�H���z?  <  
  w/eg.class  <      ?      m�KK�@��4mcj��Z����]�D*�B7�&���H'�w�*��Q❈(��9g�7w��������V�;c(��z��Ƥ['y�9�'	�ڂ��r8w�B�5C3�ǋ��p�:N���<L�&�����`�����m�mTll34&?Gq��)Bߥ:��}$��kZ�f����ӽ�����$�ywD5U����q�cc'4�u��P��Di�3��^(���4�2R+��T��$h�Ae@�?h~���P6I�1v(�Y`���5��,P�(!��AR1���+j����y��n��9�r�o�b���=����>PK
    +Q�H��t�  �  
  w/eh.class  �            }P�J1=�3���V뫸�n�-�BA���<bM30��w�\�~�xR��9I�ͽ�y�x}p���sz6p�J+3c" B""bBw�4��a��?5Y��p!##Py��A�'_�;�K�Rɒc�l���!К|'�I�62�B�t��h�0��+%����%��"4P����}��2����m��z�3�Ta"/�NM`T��թ�����	vxp���#qW���1�)6V06(.ڬ|lF�w�&��/`���W�&��n�ئ�+�!��j�������	PK
    +Q�HkrD�R  x  
  w/ei.class  x      R      mQ[KA=㪛�J3-�[/^�!�@X(|�it�fa���Փ��GE߬D��p�ٝ�]������@7V�5f����z���N��� Js�����y���T3Ԃp�LB�͝����52K�G��~u���1C)C��������"C��+�H�Eأ�ۧ�����?�+��K�{t�u��o2�	͘�$��ݜ-��&��;n�н��3t�Gg��iw�G˨?EJ�1�9�ŭR��Zj��ə�:
8�4 ��1q��
�G���$Z薱G�M2�I�$�D��*]��<j�e3P�+���]���śy�خ�]�&)�|�c}�`��u̺�)�PK
    +Q�H�$O�@    
  w/ej.class        @      ���rTE�� ����񮉚��������EE�x�$K��bJ�K��*��|�װ�Ni��[����tf������ ���4���a�8�'<�`��S�e������E/1X`�������7Xh�KhN�-��Rm�:��.a�LJe�m�\�B��)�d��N��\�.�*�����{���<��xc���]�At��]�\��������]���SV[������ݬ�9c��������`r����AC�:D��S�r�R�^[�S�|
�'�h@Id��2q]��Q(ٗbp$���R�U�Qx�ۀÖx����>�!+�Ů,�3�K<'�c��Nf��(JT����u\x�bWyLE�ԬS9�$��E\�2d��a�<����L.ɜp��P�r"k��Nxdh�Y���IgK�ieKt��{.D*��F�e�6�薽+
�$� D;�	F�c��g�?6SL�kkkk�uk��k��{�G������K[{��C\����u� �&�wX�c�������Wwn��MC;�M��^7h���ƿ_>�59ؽ��9���s�*a��LX!�%�#p�y�*A$A4�,�:�'<�o��E3�~���P=�M�[��	��%l�#�O�D���!�#��YX��g�Op���u� N�<]m��Zsi��!W�<;�!���\R)�TC�!͐vH7d7��y�8#h`?��l0��܅���^�����T]��gؼ�V~�+\�r�݅�w�J���W?Q���T���L�����u��տ��p�o��>�>[}���շ��Uߩ�P�q�����S�w��~����{W��PK
    +Q�H��q<�  9  
  w/ek.class  9      �      mR[kA�&�M�TkK6�zk����f[[��B)��B��i��8q����7���P����3�jC݁s��\������ <-�ʐo��	)�C���C"N��D�Ʃ��?�|�i����,�	�Eo�����{���x�4��܎�گ�Q�+3N����`d�d쫿��9��!Cab�T���� 4c�劘���\3p�aŽ��&R��.C}�ʥ����ʰ�a����¤t�O�w/?r��'��5��������[o��w���1��������8q��1�:�~�͞/���P��
�ivO��
n�A&64{TEi�q@�h�K%>�q&�(ܗ2V\�X�1T��Pr5NB�Q��R@SW���Az�^��	���-b�DE�W7HT�"豈i�e���	�+��i0��]��`F�ؙ��%��O �6	�#Y�t�?P��=��*�SC��������8^fSt����?PK
    +Q�H�?    
  w/el.class        ?      mP�JA=�n��VZ�ի��ϊA� 	��4���l����w� BP�GEw�}����;��������+�ӝ2��7�0�J��)8E�P]�5�B��]�3�Ј��r��&:Nf����<LC���EC`�9p�9(1�ǻ^��w+E8З�?�}$���x�f����Rm?C;썳�F�S��|���"*81P/����M4�͚���IL�J��V*�\�H���P\'���V�ȁ�	��ڧ\�(�iY�"Ri0����`�[�����t�nQen\1�����mo��	k$0�F��ܞ���-Zߚ���1�PK
    +Q�H@�P�e      w/em$a.class        e      mQ]KA=���Ge��}=����!�B��KO�2����'!�Џ��Da�p��s�|~�} h�!^�R���2�{'�c���/��r5�F31�eϟ�#_Nf�@�����K�.Cbe�9y��q��	1��Y���k��I���f(��r��;)�ID�YIOQ���K�YٓU�Kj���]�^����VDm��D���և9��L8� �Ni7=oB+���~��A ���Bi9Cȑ+n��4�4i遜*��@r1�$�0^�W�����#G��v�R(�m��P�.�3��pA�Ax��5�^�����ej#�4��w�q��ٸW�?E���/M%�d�@�PK
    +Q�H21�:�  �  
  w/em.class  �      �      mR[KA=��kb�Z��xmԶ1Q�#B	�@^|�$�t�:����$����3�`��o������ Nq"���δ��\@t�!�1$F�"~c�7�V'�N��4c�r0QC+P	��?��h��l4�W#'�)�����-�s�Pf�
8�2���r���]xX���Ú�����-���V��%�؝��e�>�sjcU�rA�Ҍ���$I�iJ�Y���u�=%d ���CG_���}���Jc��Q�:ƨ��8V�@�zj��U}�A�~Zi5�zzl��F
5��T��*�#��a�zaN�S{s�3�✮rU@�ܤ^b�#V;�(PL3>�,�e�R�QaYƗ��7�uZk�
�7�����]#�]�3��F3���{|��'I��p.�.��G�PK
    +Q�H��C1    
  w/en.class        1      m�MK�@��i��~���j�o�8��S
"��b�O�f)[��M�]�
�� �8Erx����Lfv?>_�qIp��9�<RZ�1�&,�
XVHh��Fx��K�.XɅ!��d��
W��$�����FD�$�=��	����5�Ŏ����5��"��n��B��w���Xi#�N������e�Ü��`�?�?�:
 k�*�8�v��!��yH�QOr��*��ֱF�zM���R�&W8�2����	��U�xȪNP�P���y`�����g���	(���ث����6�(p���[�~�\اa�/PK
    +Q�HmbZ,�  [  
  w/eo.class  [      �      �R�JA��6�-����0xv�H@Q��S'��Ǝ�gy� ?J��(��U�y�ޫI���|}���@z�X�*�̱�����I�-
�����R��E�4�@!�C��f˿6q�a~��lw؛y�(MCX�R�Җ2���rYtC�=�
LU�_FJ� >����a��L� ��O�X>9�g*h7��s����
!��#W�?�m��u`��n�����>�\uo����0R�6�ǖ�m��4jr3�Wm�]PS���N���4*����*��t� �X`���X䰒�!�Pdbv��`�!�-�~a�!�&<�0�0���_0�0��f��t�%�<}�`�n �Q�ד���eɉ/����9Zy��r��)�|��~��v�5]�M�PK
    +Q�H[eضU  p  
  w/ep.class  p      U      mQ[KA=�m�Ri���^�!��X(|�it'��Xg�w�$��Q�7V��o9߷3g����7 �3�+�C�%��m�!\8�O<� <0�G|ʝ1WC�?�`�����9]��c$�|�\b戧8C�P�P�P�P�B�B��C���Wʹ�b�5����&߅PTؕ?���TZM��eܻ����mD���nt�f�fr�����ơ�#
y�{��t*-EONd,.��5��W�tW�a P�6�)�3a������;���IRQF�Ģ�\2
$+Q�I�ec�$�Ҳ�e.�pBVaQњjs?�E.�=��m:5F����(�Q��93���	PK
    +Q�H?����    
  w/eq.class        �      mR]KA�㪛�e_��e�~T��JAE�/=��fc�,mc�����~@?*;�-�,�9{�ޝ;�����锑Q�t%�B
uƈ]m�6�z��}���Qv�_��rٷ���Ux�������-����V��������g��r���x�c`G��i�i24�5%4%5�&-��l�*���{.�u)���_ˡ��R9~C�Y�
�Z�3����f�=P���Q����4��P�&��z4s��ť�L/��ONG��uΥ�WE�Rmї\}�v�0v�
���0��ӡ<|2�x̐_��	�"|*���!��j���c�Y�.�rEk��� ���d>*X�d�Zm@��M�RTP�G�Q�b��=�����oR�:�a;1h�Z3>i{D�I�I0��/PK
    +Q�H��G�    
  w/er.class        �      }R]kA=�m�I��&����V�a�]�`%�AX�4P�6�i����v��.�!���G�g6Ո.�s�;�ν�?~~���[�Jy��<�u��1H����\�������so�����bo)��C�B�R�#`#FȐ�S��Ip8Q����p"G�@-N��0Q����t��6��A4幕'��H&G�a g��q�ƚ�7���^���Z�(��z�)s)�G�j�_܆��w͆j��J���Ne��e�{�ߑ�\oIn��/��{�3�p�������K���eԱg�I�x̝��Cn�~<թ� OԙF��u�����@i��:H���6kԹ����ꦝ�&V���z�|����H�UҵeF�t�%���j��E��Z'r�5C�y���B.�kL̑˭��wfh�s��x�օ?�����|�滍�O?��i����(~PK
    +Q�H�1d/�  \  
  w/es.class  \      �      mR�nA�����18�$�#�� �89�HHA+a���wb�Zf�z� _��p@AH�|���s������������'�.�X��}��6���]�O�Ā	��bD�%41XǇ�Lc3�{��Z�z��� ��X>%�ؘ��|:��R��I����a�N٢x$�$�xp$���J�ʎBGK�*!VB�	�*�͛����Z�I���#�|�(àь���� �H������r37���e��Uyϭ��3�D'�0��zr�;����PF�ƿ/�p�\Ԭ@�]�Uܩ�:��rUϲ��|55V�S�z��zbLfc�33�����v�+�U*;��L�N��b���q���3�S*��6)U�q���3��ϸH9�3.QN�Ƣq�RGiѸ��`�h5j�}���U���W����,�6S]�֬Xkw��:F�d�#�L�� PK
    +Q�H��F�  �  
  w/et.class  �      �      M�GSSa���$@AXK�^%�[p�� �J(��\9��, ��K�՛�sϹ��E����33k�[�ś[�+k�F�bG`A'K�4�bݬ���>��B6�F�(˰�l��aY��*N��|�%�s��"�wY��c+���{�ƙ^7�&�T`%SɌ���#�8�{��*s���Jy��+�eQy��S�+�%��IYV>+_��ʊ��|S�+?���/��G���S��#a+,fA��u>L�0��U�.D��0*�����5n�5X�U�&lŬW:���έx��\�|W;�5�I�����܆�;��;�O�Z�3���,��|�v>��8��{���}��~狸��>�܎�/�F�|��
nr��;w�s
�8�q�s.s��	����ot�����\��o�y����+��֧v㉭?�PK
    +Q�H�k{��   �     w/eu$a.class  �       �       ;�o�>C^Ff�0F�D Nbd�J,K��I�K��O�JM.ad`)�O-ed`Q*��,���l�\�>@�Jk��6�g^^j�sNbqqj1P!';��02010 �Js�if�8� I.�&6N PK
    +Q�Hc��/�   �     w/eu$b.class  �       �       %N�j�P�5jL�F� ^=�P�/9o���(�B-����C?��*Ϋ�����]����`����湠�:��z-���Y�����t��l���Ղ�GbΌ[�.�.\:Z�K�e9��pZP
�� ]=�<���@eei�ӓ�*S�Sp!��T��@�St��#vSj;�����+�����}&�����PK
    +Q�HN�J�  �  
  w/eu.class  �            mQMkQ=/�f^f2�$�X�5��ɘk4 )��U E� ��L�XR�D����+����$l������o�7�`��s��;�/�>� ���Ơ8���s�z-_c�Ԣ�j;h�kD��ꭍ*�Ț���#���o��A��|�C2�v�`�x�����Im��O]Jw�
⡜��q�ߡ�CҜ�o
��@B`F�@R %�f���yK��N���!ն*RԌ�W��H������;�܄	ۄ��	!]|���&���ee�t�uX8c`��!g���`��	,&0���-H�H�'q�ݖ�`ւ��w�~��#G�s�?:m΂�
EK+��.�cy�vG�����k�b/�?�a4��gMG�W	?�6o�R?Y˾���w�r��r� �l�1$�2a��(s���ר��-�m�((=G��	�;.uZ�n������b��Cٔ���wp��.<�lw�~:��?�
���b������Ӆ��oЃ"�\~���!#T�=�Fe�����2O��t'�#�PK
    +Q�H<���  ,    w/ev$1.class  ,      �      uQ�n�P=�qrc�mRBZ�P�#��u���hՅQ*HE���*���j'�_aŎ5R� �X����L������3�;�;��|���G)��# ͽ�a�y�A�D@8$���".E��G�M��������}�wb����]�DdP��~�R�Qq'��8�>�4��Č�!1+1'���K�K��Z���M���:�@�J�̳�<T֬��]�M'�l��S�<�I��g;�~�">�ݷMT:����C�@
�A1��E�]bu��K�0��P�U�k�upS�"j:.���f��<���=��m��n/
��m?~ӣ�7�0�7�n�ꔵ �(�SO@>��f�S��O�<� rV������1־�?�=I8;�IN]+c�6����u��,�OP�]=B�Ėa]�����គ����<��� ��P��^�ޡ��޳�FiR��}ŝ�Ϳ�t�J��i����*=���o2Uz�U<$V��P��h��"xcK���_PK
    +Q�HH�7_  �  
  w/ev.class  �      _      m�XTW�ρ�)��+��bE�"v�
6+XFR`T��,���j/���$�"�`I����t͖l��[���&9�3�|�o�����{���|?��ߞ:CD9T�L/0�a���`I�QVUQ]Q7�)~D�urLI���*�W���u�E�:���pC8�*\�({�ʲȲ����L���饕�����*����ԄWV��ٖ?�����V���VdG�uPZ��Ai�BC��!-'z�*�զ��^j�V^/9/%y�������K���K)^�+��\�d}���_=�,���r�Z�*(�n+�L�a�@�$:���`�8�J����e�uEu5����%XR�/a��:C0�y;�H�&��|�N� hM�H���DjAA��qGFY������Sw�l4 �4���P*	P��Ց�A�zuh�z҈ ��Q	ԙ����/-��^��G��)���:R�_�����G���K��u�{1'4;�����M14C���1jF�	*8AS �̴��:��>:���9N]y�RC"M4�0�8��׸��#��D�OФ�q�'iӂG(mjVl#�-�=5ؓ��9H�<�2SO��z����E�c��w���x�)��4�e5Qat71�4���o#��&�U��3�/�]��7R^�f�n��������^w|�a_(6�8�'�Cq��P�,yc�C>}I���O���� h���V� h$m�d�-&��S��W�x�|G�q'��T����Wv����$(����X�&��'���t ���>��/��r��� L�m�ʃ��!��P��0��p�V�mk�mk�mk��r4��%�b�<ܗ�ù�X`'b�I@�M���B`*�&W+�c87��}�p����)gc�9�Z9W�)�I�R�y�|�v�$)/���K%�������]�@�+��FY*��e�FY.۔9�\hoy��P.�<e�UV�c�+$YY%��K�ye�|�\*i�e2@�\J�5R�����:{��� ��r��S����U��\-�WJO�U�Ky��V^#A嵒^rt�d@kd �VA�d0�^�@d(�Q�A�d8�Y�-2�*��et�L�n�I�MR �,��[��&��v��9�N��y�n	A{d>�Wʠ}R�t�,�n�E���C*�;��Kj�R�z�4@�et����U�Y�+��d=t�l�~&���&����l�~%[�d;tTv@��:&���zP�@�^�I�A'd?t�ptJA��0���="�@g��k�zT����ǥzB�AO�q�)yzZ���&�Y9=''��r
��<�V��~��9��<�A���(�@�˳������^����E�y	zU^���+�yyzM�A��П�5�/��Wyz]ނ�&oCo��MyzKޅޖ���>�| �+C��'���)�|}(�C�/�ȗ�?�+�_�5��|}�<8�$�4��~n�/���Ư���m������c��������Ud��q.p�]�؅8�����n�a=��P�H���y����(��Ȕ�V��ʱC��F�'�[�� V��Q+�m���v������4�qD�qG4�q'D�q*��3��*�+"���;����8�r��s��r��rD��[�8�>��n9β_'�A��E�g�o��!p�s�6��7�P7�-o<��ƃ�k<ĺ�C�k<̺�ík�k]��5i]�Q�5m]�1�5k]�<��[�x�u��[�x�u�'Z�x�u��k<ٺ�S�k\h]��5�f]���5�a]��5�e]�"�[�x�u��X�x�u��E?Z!�Ϸ�q�u�/��/���e�7����,o��q���,o\ny��Z�x��[޸��ƕ�7����U�7^by�j�/���2�/��q��k-o\gy�z�7X�x��WZ�x��W[��J�_ey�-o|�卯���u�7^cy㵖7^gy���7�`y㍖7�dy�͖7�by㭖7����7X��F��dy�-o|�卷Y�x�u�wX�x�u�wY�x�u��X�x�u��Y�x�u�o���m4�݂�wX��N�eA�4>hA�C�c4�4���.~M=W�DS��X�m�1v���)�S��k�~�e_�c�o�.��@����B�U�����PK
    +Q�H����  *
  
  w/ew.class  *
      �      �KSW�OOw�n�H�����`�����(j'����	`�NS�+��v�"eeCU�E��8-?@v��d����Ow�T)�l�	U�w���ν�t���^Q]�HOu|^��Hu]��L
�4S��%���DN��!��� �����t=�Gf����	���jS�3�X<W��߯V�h�t}��Tfqji.sq�:�����Wf�H]��^X�����9Y��XX���e*�sߢ6���-�[�K���ě��q����Өs�'�Z�+5![n5#�����I�&	�V��b�H�����dHh�:%OX�Y�قAT�W���:�SpH�t5�n: 8(�R�z��R:JI�݂�(g�}�~AVpD0 �E�ҋ[=ys��f��Aq9��ɷ-�m�m��g�F�v�����=�5:�ɟ���:G&E`G��hD�zLM��-ίR�k�_���ÒK�5:5�����s���U�`eo���NԨP_a�+Na_vPϙ�ԧ��攗pT�c��t�rL�*�L�c`�<�:j6����c�������g�6{	O�(�ktvms�`�6l���_˔�`��`|!b^B/g[h�!�0B�^.{	3��r��Fz9�ʭx�a���$b�	3H�̈́�z[k�׿�w�c2՚���ސ�;�����C�.��/}Ox�H�1�Ƥ����Ŵk�f9��l~�J�i�B+�J���})��=�S�љɞzء�0��?2zN�?R^�#nJIϡ5��
[cE3V"�����z��a��QmV��Oh n�W�I버�Fí�3?�ԣ��+T��ŷ<+���-�����v�k�PPb������R��W������������y�{�q�s���JD[]�5'"�����6�Y�֟�i�ƴ��o	�>��.�|�X2x�X2�d���T�d��b��3�+>Z|�� 6�y0��m<��"�ȗ�&�6�; �`���p;�6~t�*�Γ�� ��%0���x
L�4����Y��+�n���s�^��������� /��|<�K`�o�]|��S0ͷ�n��p������=����~�f�s���q?x��� �x <�9p���#<�y�48ƙ�3|�/�P�� � ��/T���h�)�α�u��PK
    +Q�H݋��  �  
  w/ex.class  �      �      mR]OQ=��e�uAZX��R��e�V(��ć$��.e���6tUx1���|"�_ $�1� �:s�����gf3{�����)�Q�e�3$ȩ����T����Z^�pAX-�����i��z�$
+yrl	���io���m�?�n�^-;ĭ�*Q�R�Z�xMB�:%d�j���d���<�Z�w�R{�-y���!�C��ʛ�3�{+��bci��9�#o�T�P5W�����gKCDC��n����i�)	}���G�5U`�Zkn%Ϥ�$Ũ���Nɛ*�آN�B7f�@��$�#` �@'C}P�k3���$à7t�&��-��!�#�0�`1�0�!�4Ý�Qr���|u�n*t~7uz*T(��l�ExP�]ذ�AzNA\'���21�k�#�1f�?�H63LʠW�J�~���"e��2D-8%jc�J70a�40n��1d��0��$JV"�n}G���r�}��X|�����PŠ�\�K2~�t�.���E��i�	�H��%�7i��=���Kr���P�hlY)Rr6�?�Z�kM�2���-�9���a�M�s�L:f�'�}M��
ASeE�3q�gM�ܜ�C��f�X���-S�<C��n��y٥���T�@������I�`zR�;=���L���l��\��<��#�҉#<��ɃK���]�/D7�O�����PK
    +Q�HtM�
�  j  
  w/ey.class  j      �      ]��N�P�ϥ-,
*�(jmM�q�a�+�+]Ȇ�`c@�{��ݰ1�`�!�2�|u��hh3s������~|=��aY@�W
N�����
���<�^R���q�w��l�s�8O)OƢ�PT�k��YG-_�jշNj���une���A�h������ʡ]m�-�M��E־TRV1!ѷ�э�}���F���G�8dv
'Տ(�9�p�`� "��Lp����z�+�� $�y7ra��Ѡ�^��P_`��Ix�|F���C��0��D�C�S2�=,�!��4@�C��"˄Ȥ1����"mĻH	��=a�����(��!��5�;(r�|�"u�7D��h�xDj��W�\��[dH��Dy���Ձu�+I����1��q3���4J�.u�/0� PK
    +Q�H0����  k  
  w/ez.class  k      �      }V�Sg��.�$�����.Z�Zy��V� mQ,З$B0���Pb[k[ci���_�q�8��uF^�v�����_Q��ܓKZ20s��g���>����?��m �÷��z4 �[z�2�c8�0�p��(�1�H�(�H ��2)�) �A[��� ��=$e�6�khsw&���-�ڧ[zc2�h�V�~CO���TB ��	k֌v�鴙�q���5üi4N��*&�"A��g2zn�L�H/�6��4>�+��� �I��IZ�K�@��-��У5i�ґ�Fzm�
�������D�J�� {��H��Ϭ)ݘi�3X�=E�RY�����FsY+1���i��g+��E�p&�c	�H��f*�cZ[�W{YO|��������T
{$�5,�9�4
A���;:�]��˗p�L3��#�W�������Lc�ʢ�fk"g�[L\��Ŵ�d8,CX�4"2��M��pN|��C%��2Ic�O59D1Q�n)GP�ۭ4��0���,.pG+���KL[�2�h)�f�F3$���h��(�u
4 h&8H� �(��������S�v)�*�V�5أ�Q�+�U仗<TNA��!ۻ
��(�e/���I/\ ��G0N0A��`�����[0���AR>�|@�!�G1��*��,A����`��@�׌���5���֘�Z����z�xK]@� ���z��"�_��U�����z5u��p���A&�[��K�:"� tj�&�A� K`i�5Xд���ຽ�=G�sȴ=��{�'�{�X��
(+E�^�Ǌo­��	w��iu<f���1���'?��b��4���`�8��lg����#D�i�hI1<Ҵ�N�2{�
^�.�^��_`z�S'��.�}�g\u.LOg!ň��ݪ;�3�e��1܄�Y� eU�`�]��a������J����;ލ�XWI=�r�������^~i�UV�*m/	ǝ�Ԏ6	��� .��̇P��k��x~�O�����V�E��G�f3গ���l,˼^�dbNa˩�c!F݄/�=b�Ku�<��$UW�wS�{��{�� �LHS]�*���PB_��Z�q���r~�-�1Pxf���+Ԋ��.�������ƫ�����~},�q�f�h�1j�^�����ml��y�E���,=�V�!�,(]�;`7�'R��g1 .ƾ�9�	�S�}�Ex0�g�����$��[pط7!�K�)��*k`�1��w���ה�%��×W��۝�`���u���
M��_tT�b��=E;�s�^��y�����ǫ+6�f9�ig����#�-:�_~s��y��\Q?�Ӌ�p颱t����b�zI5Ņ�����/�����h|�J"��燝�s��O3R��;�Z�&�f�[�nG~-����C�0����s�N���o��ԗ/f�p�P錷�;��������6v�nz��b��&�lj5����O�]\a�+r����tk��c�=�� ��b]�&�;`G�PK
    +Q�H��gl�  �    w/f$a.class  �      �      �T[S�P�-�M�E�
^�b�+�D�[@@�xM˱�iS&Me�)>���ؔ�}�G9�	�Xhq�L�=����~������ F���Q�q�]�`�q��´��aO00
c�f:���67�m��'�О)Y7���/�Й����73ϓ�!@̲e,��e��*��i��M=�-�"�Y��6��(��<_0���z,����Rz�g(c�/Ր���g[���*�M�K��[�y�U�1�R%���2�*���3v�"�A�]��ؤk��݆�&ߩ%��]�(֏�gڥo�{��J�%�J8%�O�i	A	g$��pA�Ee��1ҟ8��)y"���p��1��簿V�Wmdš�k�o����_�����(":؄�	n��?J���+%���9>ִ�zL�f�X�+脤�>
"
��*`XA���Т���*8'` �
�qU�yĄcD���
�qC�I��[�q�w�0*`L���A<�q	q!�
ᑀ92.cF�&<0%`Z������2T�0)S�Y�8����W�ɭ�^,�"�5Uc��Vj�T���-��������Z
Yœ0�4���w�q��'�>Ԕ���e,��٨Wz"�:X��^:xUƒ)cQ�/#����
�Y�U��P��>-��U��"�q���^<d��Ji߰�G(U�*���Yv���Sk�
^'�R��'��m��2��J8؈~����d5�i(�?PK
    +Q�H�����  ?    w/f$b.class  ?      �      �R]OA=��.�@��(*�*�!.�Rc�$&��� !��t;�%�,�N!�+M�Ml��G�5�l��p��;��{�f~����6^1�m'�	C�4M��d��00N??�MA�a�#Ԟl2Lř��a��_p?��o���RK�SG*�d�m/��"����c*8��F���b?Ld�KS��ܾ�J�ONfW�Y�{#
�=�(��/����^���-E��Y��;�,0��6�`��{6U�m'K�};��B��u3��97�{R�V,�R�Y#��mgj��/�aa
�ܷ0f������9<�0��:|�O���bMC�D	u�cx�aC�c��D��У�Oڂ�
��~̻]ѥ�Y%�r�䀞kI� �Q���]�j�q���;D��`�
��]���1���~��t}}�r�b�9���n[D^/���x>���I�KB���%�|PK
    +Q�HR��w  s  	  w/f.class  s      w      uQ�NA�fǅ��cгƃD�ƃ��c3�8d�C��勼�E�$~�e|#c��}��U��-�Ϸw �(Eb��+��^��f���t�p"���N�Ɛl�;^��l���rM[2���ZS.Cv(]��)�Ӫ�����*�ۖ-��k�4�}����ǚ��U��M���q��^<��m�!���ނ������T�����qM�l���8�����17\�y��F@�$�����s*�XP���+*�XT��2�MŮ�DJ�T,�n�6}_��y'�"�:���_���Y�@�%<���u�� �B��>R�=��^��`[?�z�|�n�V�_�)z�åV��i�"a�,Y�.�<͟A�/PK
    +Q�H�L�){   �   
  w/fa.class  �       {       ;�o�>C.F�DF�ĲD��|}O׊�Ԃ���<F�hNb^��RVjr	#K�~Z";;3;#���L�iIAiIpIQjb��f#ܨb6Fv6`�bd� bN �H�20  PK
    +Q�H=f+�  �    w/fb$a.class  �            m��N�0�7NM�PZR�.l!K`GT�: !!��*q)łBb�x(�ٔ���w�}��w��z� ��	C��JOx*]�����}`
c1L1$��A������Jϭ)����la�{b+���n��\��K;�.+c���@G ��h��ꠏA�6�oZ^k���P3Ĳ(t5�Su�k�ݣ0��)N�l(n�m�eof�+�g���3�
�$O�r��Z]y���Ψ�/��jں���7����حD��Zd�PK
    +Q�H}zl�  0  
  w/fb.class  0      �      �X�s�?��_�eX/^[$�ʮC#l�Ie0n�u����[6�2i���3���Ng2i:i1��L��v25<i�ڙδ}�K��?�{�����Sƺ��s��W+���/��CPQ�9X�k�Z��zQ 1���7�T6Kgbj�f/+���",�jS���p��Hg-�ꉩ�B�PD��PC/���K�|y�����/@�|9¹�������
�7s�����<�]��:���[<UBf?t�6~f�sM���h�[��=�+�Ņe��㗍-�,�s�0;v�<�_(�~)�^(-�ss�:R���ĳ��L�h���5O0v�z~�T#B�Bq�V��Tʣ'y6_�!l��Y�������"�Ջ E\s����i;��tk�@Jak'�M���,��/��
$د��x^�
T�^T �@��V�W�>�Թ�jd����p4:����58�O��C���a�[�{
�6eh;�Y#���e��:�i(�H�����C~�-�:G��h����L6@d=_)/ww�3��jUm���|�FMr�nP� �Qh��(tC(
:�(���EK����R�,9
�i1A!e�T´DIo7���r���Ea/���4LD �#p���#Z���E`�"pފ�+�CZ&i���)x'C0A/�"p.��V|~�/��&�>�����5��J�b�bnv��{�,	��������R~	��ƈ ��x�A���/!�B�¨yO֬<�8'̿��<�3���������&��`�=@�]hށ��2o��1�@�}w|K=o�zXϗ�����B �,�'�6T�8MflKe��c�m+�?"z�X����O+�ڣf�&,\��?��g@�&�/��z+�;�$>����	�ǰ��ßA�����M����Ɂ���B�^�J$L	�����2{�G0�g��V� ��۟���Gx�,�{�c�GZ`{US�fL�iV�|�b��>Vg�ëdK"P��<i��*�3�MX��Dyb�QF��)���޾;N)���T{u�h[v��a�'t�9lT!�����)�`�<[�O�q�[�ü�/x=����O�1�����Ys�;��i��mV4�����>�qD�Zp_=�zG1�YiެN��ZM�(����|���?������R�u�L��l�J��0��-NYӼ��V=�2���7�7��4��d�p
{���.��Vs
�K,�%V���`���d�_�j��� ��C8�oN�if� hN�g�;8݇w��=�: �7�X׎��C������)X�R���$Nq8�8��4�4WU�XG���~ǋֹS*̟�Z��V��Q�I�&�Tm&}5� X7���K}S�A|�F�*����E�"��Ch�r��Zۀ�Pl���sgԅt�p�:J�7����;�*pR;���h'�>���L٤�d�&$�T��lR#�Ө�T��58*�^P�jxA�^Д/h����E��</�M��s��D�V8v�z,:��Ǥ�L��~F�3��a.��P�}�k�6��0�TC4�w�F�7y6��lT��ےF� �u1��7��{���~I�>�v]��܇=Q�NT��K?{�
��_݃ô��>�1䳔��ֹ��e]�N����yR���J���`Ed~3�8.v�jQ��Z�$X��m��^��f�Gp��uЀK���Z����%���c<@ɦ�!��e��0�����@T�	�>x�?M�BDa��ߒ�#F0��'3�KI���~Y�?�6�ش]Dx�L�~���#�#�t����r����G�#�#��g�jY�ucV���,�a��"��8/`%�Z�~�l +�<Ol�Kf|nR/�{��"�W�
��آl��8��*B����y�<�&�Wp�m� FÁ?o����.m��n]�(V%�ڕ�mZm��W�,��dXT��F�kx9٢5ɷ��~�*���+[�3X�X�.&b�����~�"㾑��4��AL��|�N k���1װ�.��+�
38�� S	1� H �N(�I�0���PȤ�%'� 5DS�^�]G݇�F�0�'>��j�x�!����TK��O�|�*���4P��"ሎ�eO_y]!�B��@�W�kͿ����_�®4u:�s��u�Yg!�_>�-���d>��-E4�8aEB5iK�`Z����E�?�Y[U���J/�g�4�h�PK
    +Q�H��6C  �  
  w/fc.class  �      C      UN�N�@�s�q�MD�t�E�A��("QЙ�Db[�C�h� jZ(�@| �ٻX<N�����|~� �A7w��iU���se=�����n���Tە��� �g`�3����s�����8	��/��d�L}o�P�x���<��i��Pͨ.���|���S)D8%e5u��}$���p�k�w]�����0�B�<���`���.�H �&��nQW'd���+6_����9��1o�|�ӎ�[�t�t엡_��W2c�?�5����u����m�q�j�q�����Zwr��
��)�ES����Z��7PK
    +Q�Hr�ŕ�  �  
  w/fd.class  �      �      �V�[u�{����E��̪x�)�����IH%;k�..��e'e��
jYt��&F��=ODCA��ð,�$������wf����S 6`J�C�R���-< ��-o#�孯g�������Z�Ȍ�)�6�����T�	GÉ-�Zc3�����]����߿]@;� وǍ��X� ���O��͐�IP�`�ؗ���]d2)�y�߈��"!�$�8	d���Dm�?$�H|����l��?b�<�wĢ��&�$�\R4č�nK� �f���r��on����/|���3gU3�I覘���F�1����Eb��0����Ѿp,*�8���qZ=[�l�=�p4����LѮS�Vv����m�P8j�ѾP,�#�3מ>��^@Y��1����M�J�\�'h�,�7���kY�f���T���P!M���9��Mg�� u㎘ѮM���ip�R����-'���� �s�"�&$��A>$�Ϡ��?a����(����X#b��u"*D��A�F�D< �A�"�E�PQ��{����o�z���@R��$e�7;$?SK���]�iȸDd�2M3)+�t)�2����f��j�	dﯺ�`��n�-]@?��X��e�a��~ٱ:�Ӆ���̎�A�#5�@��4k�d�0�o1B_`�TV����Cz[�Yd<�����/�d�[���1m���*J��b5�f�-�2܅�*�OEC!�ư�Ux�bP�N�3<İ.����a�*�Ab�բ���xBŽhUq��O�(�S*��iv>����Μ����N�TQS�*�T��KF-�1u8,c�a��؋n�0CC/��8CCB��GN0����)؎^fxC�x�)h��/)h�1���*�cH�N���]�g8��
�;
T��*x��6a������
���I���dx��iu��I_�{阀fH4$Z
��rx�l�VdQڒEi��e[t�Es)���'��H/��Q/�I��k֫��5�Ct��¸^(L�>��	��ğe8�pFϙ�)�Ӻ/����;�f8����Hk����a��'��(Ti�fb�m�c�����2���1|8��1|@=\fyxNE�=93�%T�Tts̉>�t1�p��w��{�I!Z���N#O�yb��p^�}����$v�.�;S����xW�\y�$q�b�;
򓸢{\I|�c���7I�Ό��DC��A�g���>�/��V�.ƦI4���e���,��$�����ؚ�W���������$��r{�I\��a��_Hb�J�=��-�Vਔ��&�|eQ�׍�=�|���&I�&7����h����(Vh��J5�R%���#����t�l�(���T�������;7kϵ�W�	���ǹ�("r��"r��.���z	_�R�8����f{bA)�H�s�a��?�t9*ݚ�+�����*EM�OD*%M�$[�V�>�:�O4���{��X���5WӐ�&1�jU,AM?�ˉ㟼I����\������PK
    +Q�H��kN   Q   
  w/fe.class  Q       N       ;�o�>CvF.�hOO�hO�hOF�DF��ĲD��ļt}�����F�r��Tvfv6F6V`dad`b`1PK
    +Q�HFca�  )  
  w/ff.class  )      �      �R�n�@=��5qL����P�vZ1�E%H��P%#�"Q��3	S%��v�~ _¦[ش<�~ ��� ��(���=�>��������&C��^0LՔVI��	�D�ɰ�]wű�>ׂ�A ��DR��,`(�e��'��m�%��0�'�8z��xW�U��	�,����W��E_p1H�EŐbXc��5����|�8�G�
5M��>;8�%NgP/Q c�[-����Bтcᲅi�z��	����7��%�RJ�?���bX�(͈Fv^�~�G'
H�Z�U�{CUo`h�&��	f�}�����G����K���¢�L���m�`��,n٘Í�u��<V�X�*��8l�υ�jk��"I�c���ʡ�<�h�(z�����s����ӭ�z~�(+ﰱU2<2+_0�l�b�l�a������Ƿ~�=u��C\����X��v@w:e.����~�d�'PK
    +Q�HX]�_       w/fg$a.class               �SKOQ�n�qg�QF��(��
�8J�
�:Z|D�A6L�X���n\�\�2qㆍF��ѽk5�G���s�@��&�<����wΝ����; pIC��u2H��U9��fP��	��0)�<:�{�+���A��x�|:9:y����)7���w��[�ݹ ���\�Z�3��N�y�bX	���V*��+AȰ���wK~����烻��t��c�J�����f
�SA���d��.�n���re�X.����R���l.l`����M�T�b�� �+��w���X�c�F�cG�f����8l��;8ڈ��i�l���h�Kd�W��D�Io\��������]q��{���i����t�j.�c�	I$͐�L7EJD=��<����щ^{�栁�8d`�0�&#̠A�#�5�wX�~]0Ѝ�&$p��nd�F@k\�ڙ^��H�� �~*�F�Z�`���z�~d�5���Sv
!@�I.�Sň��Tq�1���5�LUq��et���"��C����Ѥ��&B��y���k�EP'E�&��PI	�%�pj,%��Oɽ9��f�e	�U��V�[-���NJ�6[�^��+�~�3�[�����[%�Oд���U��4*��>#j����pl�"M���V�>_��I�I󓏮<4سm]����U�ԚE(�k�ؚ���ULyaL^�A�O��]�ѕ��]�jK�n�H��I�f�%�ӓ�J$�[�Bc��:T�1���2FK���c0�'���؉v\P��PK
    +Q�H�]#�h  �    w/fg$b.class  �      h      �R]KQ=W�mu�վ�L�r[���cыBo�|]o���k��
�>���h�&�Kxa����9��~|��8�����K�wWLP4)��x<�ă��C�>�MGx�v;A���R����>��C�{�o�fG:#�nK�}�I�؈ߵɉ�Rs�w�}��h�k�4,jHhHj04,1��y-\Ъ��ME��K�d��	���8�Pw�-�q'��5��/�Xg3�t�<�bX3ź������ ��v&vHc7��t�jТ#�Nn�|�jO��qB4��2� �T�H�b��u9���)�2F�~ƞ}<F��ч���`��a�~B��Xy��+J�f˔�4��2��y��M2�����PK
    +Q�H"G��      w/fg$c.class              �RKOQ���ێ#���@ FL�����CE�CA�V��a�NZ�D�pk�ʕa�&@Qk�/�׈�4�&�I�w���{Μs�����&�Vd$x�ؘ�K��1c��f����T[YK���2c)�t:�S� �(�êdњ���P��e�|�Z��'O�2�鴕5�񒕠��@�L8�����J�zd=�k�`�� A-	s�;cM?��;��¼��T�'gθm���X��b��J�s2v�o����8�оo�x�)J`M��S6����hڏ�w��|�8[U���D�8*P+P'AO�v���Vqf�i�v�g�c�ܼm���9���b���Fi��U>���N�o��E��j�D���z
�
�2�1�L[x�U��)���(�������Z@�A��w�ጂCg�^����.�p:�d4⪌&\���C���ze��c��pSF=	�R�{Ѐ��lzszb�?^�b�d{�|�Σ�7A�����0wI��}�ʽ��9��1��=��W1�qG�b@߀�$6Y��U�ͫ�Tz��9��
�R�s=��ٚ���_�޼ŕĒE��W0Ԭא�����#���d�9��[�9���0��j4ì��5�8��>ś���8郴���x�S��
��lW5�Hvd�jp�k0��e�����:5�-^K;uS��jPu��g����^�.y��[?�<��6�%�E��a���҄5�z����i�*M��B� PK
    +Q�H��r  4  
  w/fg.class  4      r      �U�wU�&�d�A�ЂY�$�TD
.�V������N�i�,&�qE����".��`�����x����꟢�;3I��y߽����͛9���� ,�Q�0ׅ����f��@G#��9eEidŵ:ޗL'�[ɶ�R�qm
i�J��F\�W�zN���e�$�3�H>�n�"���֕T#�LN�lNvi����"ҼI���:�j*��R@��	�?�\J�ȗ +�d^��Z�r�A	����d��L���1kK�U���'���&Ȑ�t3Z�*��B~$��F9�ˉ3�o�ji3��j�OM'"���ZVOf�Z1aUҺ����'l-�۴�^���ɾ�z5�ӤfL��s1cıg�i��<�waG|�U�x��9��pT޼��g.=Ӧ�i*SP����8�&���b��t���H���4��{y�Tȕc�����?���;�;���ݧs�>;����?9��64>>����J	UfJ�%a��%�J�V�,a���n�p���$��p���n��������f}dtF9+R\Q3=R�ʁ襟Y"F���?��|�f�J :���U�ܨ(�Լ�VʁR����='�c�f�5�i��*��%�v\IibWԊKq���(_��V_*e���<ϩ�Ѽ�Tj>��)D'ݪZs)n�^n�N�^QsW�S#�ȡ��Z_�w��*U�e��P�P���aC|l#�
�x:݇��Ķͼ��m������W	�1�A��ף��{ٶ��,`��}��~^x�!Π1t�DoK�Q�Cڍ(r:C���e�c�0<Ȑwc�1�2d�؈�𘇼<��z<ꁂA��ɰ˃&<��]xƋ����!�3<��ÓO1�f���4���2]�1(�������u_�e�)i�u}j>���������:C��ϱ��lH�8�
Z��6���v�e�a����`�	�;
�}I�FC�5�J�f�Hz�Ǳ1��Gi�'�Ṅjq6�'I�9�|nCS�/pGjN�D}�}�X%�O@��J\���GQ��8�W^exmo���C��.��+�J�Ө2��T�1�~�x���E��jE+$�$׍�16�w�CcX��C�1���v���͟+��uxM�`�������c�"Ÿ�F[���P��� ���'��
A�b��m���p��U,�Rr�)�P���Y�:��]-��6+�����i|(9�]�s`��G��T[�4I��B�g\��G�"�'���8���]Ӆ�o��,���u�E]��"��i�@�%/�cW��v%�]~��`������ˍ�t$ǰ׌邻�v���͗~��앨m�����5���1g%ִ~���Z��ZrPO��+r�DW��B4�,��
��V��;m#���g���_;�h�y���/PK
    +Q�Hv�!p�  �  
  w/fh.class  �      �      u�][W�g]ޤ�fcbU�ƚ�mJ��IL+��	H"�j_\qE.�\��_��Л\���F��<�}?J?D���n�����ߜ9sp9;���"J�A�F$�c�D�X�x��>�b�x�u l#͕�5�fߔHZ��j�[P��;6M�Y�N��h���t���l��v�a]�ƺ�fF�iZۀ-��De�h-� N��T�v��'�̞�5uê&���Y5�K�jgߴ�l�b6m ������gV���ۭ���co�ҝZ}�l�GPڇ�Oj@M�1��mMCv�U3�u�<����t=������L����t�$��k:������:_ʥeM�JltY���ʨ[XÎ�r�Ⲝ+.�eS�\W��b2��`o1�B�E^X�Ħ�G��RN�ʇ�n�M;H�4���4��Db�7��u�Fq1N��7�7��<nT��>��vWN����
�hH��$��)4F~��B�p��Bh�������i+L:�lv´θNU656{aڠ
\J_���{y&Ӱڶa�e��1�6m��M��s$Q4D_�G�~G���q���	�o�"�O
�	8*p<%��]�?_����_���3�/�?x	8�|<+p<'�*�#��?x��K�U�?�^�\ kg��g�a�����V�>#�-�����
\�ߠ �?+Q�HZ$"�����N�(�E���yX8o+�32�yjx�e��+<>�ϻ�gy���9�y%�w�G4w}�g
{+����N)���L��x�8���{uE�n�������Y���f�8�o�WCux�*U��uzpB�Z׏�1"Q+rD���yL�~���<J��(���G�D���h���ڃ�d�*���.E�����$;5�ی:��ۜr�������y�/��-���h����& ��W;F�[o��2|,�<�"/F�?��\4����O�������/�<!]�;&���1��>�?{L�_�e�PK
    +Q�H`���  �  
  w/fi.class  �      �      }R�n�@=���-�n��M�C��,i�pmA$$G�x@��"�ƭ\�����@�G!fm�Ҧ�0g�9k��o? 4�Āa��b�a�y�=����/��u�й�*����S�St�^��/G����#QO޿�H����>�)($��A�$5^��c������(=���Y��c�0��t�ut�2�݋�v�������I�W�Z���W�����aR���ly��t�l�{���̱�Öp��X�XA�Ä*��(�ʱ���%�4Q�-	nK�$�,�AX(��)�.ᮄ�E�;��_�!�e*Y��Ė��$�Y&7��4DY#f��.�֡C�\n�+�(���)v� I�I�T�JL�̅[�+��Ω�L�B�t����`1���["��h
G��-�jg�Z�_�\Y�,���w\�4EҨ�����%�O����F���7Sܷ�&x,�<���7%g)oM�������d~PK
    +Q�HI���I  �  
  w/fj.class  �      I      }TKS�V�.�,#D�#J����
a���i��<P	�<	e�K,1�챯�tX�O�Mg�a�ݘL�а�"�M�Pȹ�������{�������v\�bd��Z"ְ�c�^L�q��8���W=�����j�T,7�p��K�l�-ǳ�r��8�d�K%��0��|���˹b2�+
JǛ���^?���$O�^nY0��y�ZHs?S	5�yEH+j���ڳ�$_I��sn2�f)1�S7r��n�{C����}��	��w
��y�璷֞�%�}�����n��o�sՂ�ό:FsK+�S�v�A=e�ϥ�^>#�R�����9z��˩�1Q�YMf�p[�pJ��ᴆ3��pV�9_k��Ч�^꼵��=���`
z���V�N����G[E6�6��I ��6�Ѧ���!��	~�*H��B�)��;0�~/�w�9q�����`�w�Ǧ�䃤t b�SB����/�J�JN3�#a�K����H�����^|o�c.��Ǆ�%\�p]� R:qU�y� �C���~�pC�%O�nI��c7u��Y��#W&��>�É��?���_�T�8Z�@R*1@|��؉Wx2���ف�@��;�6���i)`�6����`��B�]���fg{�@[�k��E��ޓ8P��,YMѺ�<��o�ۻ��tSy�oB��� 3/��ؠ�B���	�F&TS�w_�¨�����N�od"j�j3�k�1��s�U���aS�~ע��\�5��c�/�E�R�b�	��Z=Ξ�����X۸��R�#�ѽ��`s�e��	�CsÂ�U��o����PK
    +Q�H-�"  w    w/fk$a.class  w      "      ��MO�@���SZ��~�j��4��쉄ăƃ=-��JhRH��<��ă?�e�%ڂ	�lfg�gޝ���z� p�>Au�[�����'�?���88K��� �`�"Bw*b��l2�
��}AЖ��'.��X���-����6��k���|�aec�X���[-�.�I6���=�����6����Z���͢�`�Y�G���8���m�R�=��:࿝2��7�B~<�2-q�M��5R~��^"�^V�*2�˺M'�T�
R�h�����Tj��)��J�x�C�{�r�x����PK
    +Q�Hv��l   [    w/fk$b.class  [             }QMkQ=�d:�8�&�֚1�Zu2i2�o���XHh)E���6c��Nj��?čn��&����J�G��N&-:p�}����}�ޯ�_���m����8� ��]���PA�+�c��pq��;wƗZޮ��l�z�����Ue<axz{{~P#�`l��?��mc�ko/6k��Ď��s^��n��������V=غ�_o���u�ÊB����-%͊�+�:N�8�cZa�^>�Px�����,�r������K�a��M�i"%�Ƹ�$t���)�ML`F����r�� p1�,.%a� �撔ؼ��՚� �[�����|��1�|�Rr�0��_�� �$�S�1g�.;�J��Cٙ����DmD��1f��Z�n��E���)�g��Q��F�5�C��ş�bݢ�Z�[���ېGnEv�1�I��LR��}�FX|d����ÿV��z4�|�H�ů����p]�Z�t�F����q��+��+���c4�1ɜ����PK
    +Q�HO Es        w/fk$c.class         s       ;�o�>CnF�D Nfd�J,K��I�K��O�JM.ad`)�O�fd`Q*����,����>@�Lk�0Fϼ��"�����b6F6`d���	b1pI.�;' PK
    +Q�H��_��   n    w/fk$d.class  n      �       ;�o�>CFf�0FVO�hOF6�h'�(F�D N�d Nad�J,K��I�K��O�JM.ad`)�O�jQ*�0F
;;';;7#���BgHFQ~ybRN�5�Nd����̼t�ht{�Jm�S��*ϼ��"�����b6F~F>`p� =���� ��� �f����T�g���j����,>^66N�-��l� PK
    +Q�H�$	�   4    w/fk$e.class  4      �       M��N�0ƿK�$�)��7;�D�A,Y@Bb@*�ۺ�Kp���s1!1� <�Kz�ww�;ۧ����0A.�_L�u��DQ3jNi�p٨}��YyA��'��+�x��TQ)g���Z���������܅3#��H"�DFH����G�Xg�R�c�^p���]��SU���;�tSV�mu�2�zȩNHv��-�[��,�����ɀ��'�>Й��>a����PK
    +Q�H(�~  ]    w/fk$f.class  ]            mRkoA=��][J)
�GkU������4��M�&�͖.��ۄG�[v�X����?�xgX-M:�9wνgn����?�ȣ�BS1�BWqCŬ�$C0�yϠ�����2�E�T�o��C���[f�u���(����gZ�z�fT���d��&kU�lQ=���9����)00���6C��?v����0{d�ع��vs�;�DmN��ةSI�M�פ��97$��e�d�����.c��T�~p�G������h�s��?�L:3�<u�,sYޙ.W��pX�N�^AGwt�s�r�qX�ǜ���Ʋ�[XC�9<���հ�5)�sx�Qn��r|HO�����-gH_��u]{48�<�R�[ȥ�P��cԏ1?.�IrktB"c���9�8E>4�_��K_���5�Ңr��^@�h���\�� M@ɮ�αs*/�H�JS�� ��[�`��ΰ!�$	�$dS&�$����$��a�$9��i�dy��xزΰ}�;�X���dE�m�K��PK
    +Q�Hk��    
  w/fk.class        �      mR�n�@���BZZh��m�Kښ�b%�Di%$�> �<-f�L-���5���|@��_elp!K�s朳��G����pG mW/2����9�$�%\�Gh�Ox����@�������ƿv��fhOm��^�(�;~t�5<����%`E�����n��@'A?����"�V}�'Q�X�x"�T�$�L�DY�"�B�bW[�;�����@�iz�Ӑ�����i-?�V�)�c?V�L���ڞyM�8�հ6-��h�����깫�g,���ب�\�`�!��},Pl��55k�|��Be&#m	��kN.�-d���>U
/���A-ٕ�M�ewp�d+�+j;��b΢�����x��x����3�jqj��N�29��L~%S�ǥ��?������r�.��Kޒ���;r����g��PߺPK
    +Q�H�	���   �   
  w/fl.class  �       �       ;�o�>CnF�DF��ĲD��ļt}�����F�r��v&vfF!M��Ғ�}���k� ��ob��f#��J�I��v@h:l|��e�[����d.gpfz^bIiQ*#+0� ����\ '���s00  PK
    +Q�HcE(!  �    w/fm$a.class  �      !      M��N1�O��q�V,��3nLL\��/P�d萶0�\���|(���8mN{���ޓ~}|�@��b$P��F�[!�15���h��ZƩ4��i<W/Иk�� �c+�+�M�R&�K��|R����n�>Kvsm�Y�Ki��I�Xf��@��d���Z��@���ז�/Yb+D�b'�n�0�v��@�����[mf�u� "tУ�$��S#Ɍ����LW���1�&�tN9~F���*z(�'���J���j��ȵ��6f8��i�F�s���7l��)׈{l��PK
    +Q�H/4�x�  �  
  w/fm.class  �      �      �SYS�P�n�iX�"�KE,)4�hY�*��M��[j��0M��+|�� ^x�)v����G9���0�'3s��󝓳ݛ_��~Ѓ�:���&�?ֹ��2C �,�Рi��0$5c�yCX�"_4�{]w�Ŷ�g
fvM�2-=of�i#k�q�he�k��\^��va�!�b[�0-g�ء�Y��VIrT<g��5�)���r�X�C�	7�Y3V��]3�O�ݴ�`h8�l�u��T*�W�"y�[:l�����BR���mU�SU�U���DhԬ��$��1�i�����h�8�q����"�%��W8�r\��q��5�>;PR��?� )O���ȺXgZ6�d��W�Z���&�q��3��S�/���%k{�����*B�G@�*�AB��&	$�T���㞊:��h�i�*��!Q(��~�:�H�c	I	�
b��R�ɐ��.	�V�@w0"a,��xBG���t;�I�2
��p��C�����[,��Ĩ�|4�}0,�!-� +c���*ݽ�y����^;DC�K�x���6��eL�0SƋh�Z�|(����L�b���%4Uн��<1#Zi/��b��>	��1���D�)c��p3��O(q� �}�W}K�C�磆�Hˆ5��w�W>�������������<�Q�{�r=$�S>��������^�B�t'-�~�?PK
    +Q�H�����  �  
  w/fn.class  �      �      }SkS�@=m���X��@+֨���-|T��N�X���%-8���?��'g�*�P����z7���L�ٜ=��ݻ�?�|pV�����/��&=�7Y5̊Z��f�����002H��D�V�^t
��$�X44`6oϘ]Y{Z����L5S��)5o�s�uB��K�P(ʢ(��:y��)���y��SSN�*��V�0K;ܙ�c���RI�Y3C��	�B���(����R�l*���.�V+"����g�tƬ�f�V���@����{d��4�Q�#ۣ�G/<*SsfU��i�F�f��;9vq��h�h��˱�c?����83���#��h]���2�N<z�ag$���>��lVݣn���4��o�kYK��ݸ��ga��I&����U1�J�%�z���ƶ����m��ę���l���[j .&���H
��&�pZ��:�Q/F>2�(㬂�)؆�
v�WAqa�Z��@�8�� �1�)1����#0*`LF��	�.�WdD��K��qC���2N`\�[KZ�Ѕ����ݶ@��t�\2��?�1��uĒ�9zk&f���U� ~�d�����.��
�Й�x������񡆎t�Z�2�/��2���Wp��/䛇��W5t��I�?�[D*�_Az5��j�JB��H}�����	��h��D�5KUd��~��:L.�ɿ������_��n
�V09���-�������3w���PK
    +Q�Hrl��  v    w/fo$a$a$a.class  v            mP�J�P�kbo�Fm}�]i�ru���J���4���@�w��?���7.f�������.��x*�xH��z��H�K��V���s��Q%`/�kθCF�ka���C-ѐ�M���#��b��"���%O�*.��,��(�`�Ks9�s��?���{.���b��z�:h�7O�Y,�>eY\L�,����� ����:z���]�݀����W5��N��'�M��w`�?'�ٶs�Ke��C��PK
    +Q�H���3�      w/fo$a$a.class        �      ��]se��ٗdY$A�Rߨt����ږ )��-�Ԉv�n�$IZ���p�+n��Lj3T:�1㵟�!��ݶ(�d�w��<������[ Π)3ӳ��.�Yx7'��Bo�����:���8�Rd[��S��,0X��V�]�����X�����*������R�tX#�\����^�B{�Riym
��~Pn�h]%����fknc);]�ze6�E��u�6T_n����R��j�7�5spW7���]#O�w����MW(�Y�E9+=Q	(8�:��^j��WE\��␊���*���SqBE��7U���m���+��R�οj#��p��;aZ(:�	i�o
/�N�m��2��;9bN������F/��N�;;��t�2vT��l�ܣ�W���)s��Ѱ�=<�������!Di�pԑ��Cc�g��H2^g��8�P1�vC|�>�e�YwF��� $1���|�!��e|��>a�Ou�HO�r���|�e�1r���'`��&�%��eƕl\d\��.�`\e|��$
%�������dX�dL1�5���^��`�����������i�p�>�}��F�d��&��
��6��, �ʬc�����'�:�<��$�6a�o�֤ݷ�����o�Y,<�5��Fβ;���:��Y)%љ�u��$��l�)�a������2���0c���W8�B5�|�EeD�)i��eȆ��`&�2F�+�/�/j���f�z���٭b.C��N܃,r�L7������#�P��!�i�7|e$e���a�O�'��3�[!p�g��bcQ/�*���ű�__<g�I{+כ[�}�vJ�=���K�r4�.��^�Z���q�S��E}n��;��t��4�;a�L�{�a�7PK
    +Q�H��+�K      w/fo$a$b.class        K      }TkS�@=�ʦ�b���*ji�*�T�ZEE�WJ�6P��ķ�?�_С����?��ޤ������>��ݻ)?}���dl��$�U�Q	�º6L;l͗Jf�ֲ"�)�%�")vؐ�xN7t{@B�HY���BK��B���R�Z*i�HZӴ�k�r�9�6F�$Ⱥa���y��g�5QT�|bxqZ+ٺi��֣)���ZY���ؘ]֍��^�rF�M7B�}�PU��t 65�rL�����L��.����v�lN��n"-
��%�[`�@�@��>��a�	t8B�i�}$�Ԫ����&�%іHg��KR�5�1�/�F�!S
mk��)s�>ϛ��3��Ѧm���o]�#��	��f9�Ȕ��L�j�ښl���"�6f����=�q���3LG�L�����Z�� ���B�Z��).9�p��l ;������`�8v.���g6��g/�� ǆؽ�0�G#��~�q��]��G7�ݸb��@u=��8ǎ�*�M�+��-Q�f��p�aR!Q�%0����S)H�Ä�^<�O{���oO�~q���C+U��,����p4,��	�؀`�D�&��랧��䝂�j�X4V�\4���PC|����tVaV0��<���'�� 1��H�G6����2�t�WA&���/x[�B?�N/!���
�j�V��{�
r5�����L�B-�i��P��vx�tp�Zǟx���=&�HN�]��<wB+x&�x����7��/���\EdrQ�c)��
��(�|./2��W�t�wwRoh�h^Zo�'�H�Q��Mz�cd9�C6H��C�G<�f?�	�4�PK
    +Q�H	�p�D  �    w/fo$a$c.class  �      D      mR[S�P����QʽR�F����xW
Z�h4�����>�i�	S&��'���� V���۴�:��~����=�����/ ��T�-�x���pE@dY��X��]��k������zZ�}˭:����!uM`���!0�c}��������셮�	�N��*;�
��=�*�~P���^��^����GJA��'ݲ:�����G$kG�0*�ٚI�,!)ᜄ��Q	c�%LH�$��'�����Q:KtR�ޛ��L�	U�'�&\�N�)�t��.�y�t"��>�T{+q���N��~�[V�R0�A1\f��`W@pH�<�,\Sp�$���*3-���E!�9�`�)c
w��HC�qwedpK&]��>���I\B�a��6�-�~���C��dx��6�f�i�HC�$���R|�Ni��_P�!>H~$�?D)�Or�C,��o�N��������kWCoq����&ʚ�4��#M�����t����Xkc�����3�(���bm��x��3�y�P8ާ��(���_�ie�w<���d&�R��3Ĉ��#E�v���_PK
    +Q�H߫ߵ  "    w/fo$a.class  "      �      �V|Sg�I���)�)�ti [;h�Ԍ�l�R7�G0@�HW����&�rK�v0�17��5u����MT��MW��k������-��_���{�$m����?��}�9��n{恇 ,m��k{6Z��l����@�X�@�mhw�kk[D�m�ֶ��L"�cB�*"$�[#]�Й�$�����P ��U2�U
0�w�)5�-�['�I%�j֨rR�U	Ĕ1uH�/Z�%5��-}!'�b�R!b� ��憒Z���i�Ù��^%<�Vc;�I55��p0�M�)�:-eEq4Exh�r2I����F�$UJ:���'>>��&��iy��AQ�Y�.�����:ߧƲ���-&r$U���uH)	9��)�LVΎfV�u�Bu;�19�j឴���fӊ���MʩDx��!e$�j)�ڢ6��*	%Mg(��T��e*ʧ�h_�U�G�dlV|�LV�Y|4�&�7��򾨚���ZCQSTl�G���:ڤ�N����H��U� ��!o�h���8I!�\D�2d��:�Za�Ҙ�U�P3l��e� �Qi����N�5�d����2X`b�A3d��S��!# kd[�&a�$�$\%a��k%<_�$�P�
	�I�^$���%a��u�K� !"a���J�J�$a��-z$�L��%�J�*��I���0%�ԼhySH�ܵue�؂�������ٺ���=J�u��J�#jԲ�˘L\#�-T��E��b���n2-�w":gH�P_n0�#�H��@d�����
���\��(-h-]���YyL������^��T~���D�x[�e7B_�O|�v�9/g�:�Bq���l�n����M~`u��Q�T���E�:�G�Hds�H��=3"g�奕:T�͋���{��2ͮuG��]ƿ�x�˕�(��i�����J;0j8��C7S��KR7�������Y#�5�sW��C�&��V����V2�/�J�B�*��Q�Zs�U8F�q�	W���!����°����������8�5��Z�^�Y^�p�!��un7�2�fh@�j�e�|7�dh��Ej�h���:�n�or�of�����-l��S��ܝn�ah�[�x1�ոˍN�͍�x�a�����F7���{X|/��8�nN�a����a��|ʉW��N(���~��0e��q��p���	���wBeQe��O3��p?ea��F�9�c�N0�&\�G��!�/3<��=����va �r���7�^�︰���&�w~��d<�B?pў�%�����\��(�c�`����1�p���.��4�N2�ą4~�B�t�|������#_��~Z����U��ww���_3?���RJzMR�d��j"E���
��P`xy������V��&���:�F���yK���*ɵ�����I� �D���9<��`U炖�EO1\d�'qS����ƞ~ro$�q�}�X9����V�+����ȹ<��I�q�r5���J���ʖǿ�(����L
'-l]����uӈ�O���M9��Öß8�~ӑ��~H�TǔX�w�Ey�QJ�� 7o})�/��-�~�q�uk?g���j۽�)q�$���N�r�Y��a8�l^xr8�t i�B]�?/jV؊1�%�8N{��,�J�O�
g�s8[T�sx�(I9�=H'��y�I�����$M�EA�B���+�g�Ko�XJ`�F���q�&|��yd��^�ʶO�Ķ0��F�Yl�:�'���`�?�Wl�F�?�ޑ�I�;V��>�7��NHD��N'Dæ�)؎����vhJ4[���􊲒�YQE�S����WQ�i>.LcW?���S�*���~+�Eo�-�ۯ��N�y+�������7ڧD��Y�1�|-�At�Q�?�E��#<�q��l��_}F���f|�$.�M<�Sb�@���0���iJ,��$���s��+b��k9�y~��w���>ӏ��C�AGYK���+қo6+B;�y���BtM��p�	�z;�Zؼ��?'��k#��L1�	A�S5�g�zZsNn��{��>J�s2�w���v�ƳF�㠐�5�3C��o;�zn���?J\dnι�yIEsI��V#=�c}�����i���f>Q��R�!��vp������$�2��c����	H��Ο9�dЗdD/l�����c�"D~��	1J�2��PK
    +Q�HU�(,�  �  
  w/fo.class  �      �      �Q�N�@=�ґReuT\PڂV�1�HH411�@iJHkJ�~��0��~���Llr�2�̽gz�ޟ_�A:r\'8f`&�Eh��A���~��KI�g^�F�tm��m]��2�<�6Z���g�����1���u=� \ɜ��$J�����q�q�c�c�#A�3�kKj�[�i�g��ZCk0dU�Ge"��q�9T�.��,g�D01����ĸ����7_���}
�XQANG^A�¬+�C2Rؒ���0�����bG�"J�/�^Ǣ}mb��4\���}s0���Q���k�}�vIA�|^�TQBaOA�R��PB��s$-7���8D^�O����?������*�cU�TY�p �P�,i�%R�bX&/I�PK
    +Q�H��z'      w/fp$a$a.class              }S�R�P]���(P@� VE)M!�(*�
�T+�(xK�PRJR���?��'t(82�>�Q�{F3�W��}�ɯ�߾�_F����q�����lǏy�R�q}3'�w��qZ���e[��@ͨk,�1�Z3c��Aa�T2m:#2$Y�����{�ƪ�g\+WЋ�]^%���V�tF7���S&ɂ@d�ɧ���<�"�% [�?m�䮲��_$wA��`�zѰ���j�,��c�({ޔ�y�h��M��e��V1��DB|����;}�D3񫍆��U�A�g;P���;���5�[�P+ᔄ�Z$�$��p^�	m.J�$���O;n~g=��h��D��r���.�������)~���%�:��31;O���7|kŜ�̬��_�&��2[����>ο�T��.�S�v���5�tm{���<��Tq��:�z�(C#C�q��gZ�\c�Sьj2$gq��*T�Tq��r��AGq��w"�B:w�Epc�z1�p�a�a��>����
:0� ��
4�+Hb�a��	�3�
=e�V�'�Q��]�a'Gw_ٽ垀��m�.�gz覎.C�!Z�~�(�����>��4� e�%�a���V�|B[��h(�	'�������
f��1����DdL�q���zg7QJk�
^1��똭���*0ؙa�j�����b�^j_�0��	=[H�n!IdV���̲��h8��X�o�����]��f�LЧK�n$����B'uZV��heݨ	�ں���PK
    +Q�HR@q*�      w/fp$a.class        �      �V�wW��y$eH�4[���Y�P��ء4�DAq�:Mb;����3��Q���
Z��RЖB�I['�lQ��lm(;��e/~�_ �of\9����y߽��w�w�}#?��G��
�!B$�%!�TA ޽W�Ow����i�鱊��U��>�ʛ��c��Y���	+k^S���)�N�2'�X��:ղ3�T��͓��F5��&�bΞ\pV��j�M������(I�lFde�y�bJY����#fj�l��Sy�X="8��k�L��.g(+Z�E�y�j�+鱢]6�t�����l��+����9`�|L�!Y��-;K�2���qc�H��X��#Y��XvQAgS�.:�Y�`Mٮ�q3�\$�[%�ꅢ�V>G{�YU-����P-���FHH�<��{�mIP1Y֔�{�%O�ǖ���aYY{.	��@�0�Us��C�L�J�v���9&�)J޾�%�	yY�O�t��1�:0��\,�h��Xuq�ţ�u��b.װ^��5tiHhب�U^��5^��u���z�hآ�GC���ޠ�Zo�p�t*��B[$��&(L��aal_�����	��"ޝY�,��/��I��)X�B���E*$�r߮�X��N��Y+v�5�ǚ0�i�B���U�\l8��͊���6� �Œxƛ7����&�^�gN�{<٪���-�[���U�a/�q���m��n沬���٫��gq��clu��Z\�UB�aH��s�y�v�OH_�E�*-u,������������p!JXKx�
�+I�+	)�U�mX��M��� -�� ����F�7өA�#��e����:.A��K����q%!�Q�1���tt�ұ��؄<����(��aj�:����:6�ho��ø��I8N��c��>A�$�S�O>�^���1�q��>�>��~�+�A����0��y�m	9�>�>�w��Cx/�v����z|�p7ዄ{��J�Z}8�v�A_�`��<�K��D���F���#؍�NFp#�H�rx�0D&�]���f��.��Ϙ�.��b�,o���)���5V4����i;܄%2A�_�g����ҕ>���T��R�Ke
\*��R�^A����C�?����d�]��=��u<���/�:H��q*��1E�!�!�%<�#���x��'o��K�*�KU�3�DM��Bh�'tZé�{p�,�g�cp�^�L�w�O�����~����������5̞�~�&�������=��b���d��o��Yԓ�tD���)'��tb��s�D�@�����ʵu<�rx�����>}�T.�C�/���7z��_$ �λ�,�E�W�5��H+öE��"�3^sW��YÅCtR�wu��u�����^�G�e�Y����'}�:���x<����I��c��7�~ZK�6����Y|��j8w��gU���5�i�����R��}��;j�8&c��õTh�ʔ{��#"���\��/W7N�Wwc�,nL�a�``S`��x����Iu��������q9v��?�|�y?���xV���ͽ�EΫ�c��ؓ��q��Kj�])
w�W����5w,�_3
�l[מ�z&�Ǹ�@�b���å'k0��i�g�X|�n>�����^�D|�H�~��o�T?��Zu�Ī�[u
�U�GN��NL�Pצ���nF�|�v�'�'�����e�a�c�^�=�_#�]�_��PK
    +Q�Hg�7X�  �  
  w/fp.class  �      �      mR]O�P~�=k9��l*�N�vӊ�Z�f�d&$$^鶒�.]3��M0���Q��t ���~��<��s����� 6�^�܊�(�  v�]" ��.��{a����(f"�ˇ�8�A��?��,Jb�$KI���������Dq�Ƒ�r�v�`�g�<�u/R��/���������X�X��.Q�X�(K,K�PJgf�/��p:���Y�ot��|gO�ޘ홭���U��/.���.��|�;<��ջ����E� 1�`is�y�W(b]�����<R�����hZX�k��86n�ec��yj��FOx��� �5�����ډ�0m��(�?Xe�~
�``���1[�_��N�x�oN�_*��ݼ!��{7��@_u��	6O��o�_�|r[gxs�W���R��u��=�s~�m���o9�O�Ili>�V��`|��iZ�C/M�PK
    +Q�H���)  �  
  w/fq.class  �      )      u�]oQ����ª��Ԣ�j�.PE�V�VM�`� ��^-t![7�
[�֟��h^��Q�wX��-�yw�����9g����o e<SЬ�k���B^ɪ�����iZ��Gsh-Z[aa�~o�<�o��l:��{�+��Gw<�i�^=�g����N3`���[���zc�4�N+$����0u��qR�)s:N�'W���h�k������m�8L¥kX!+�L����	˚]�[�.����bEM솱���:
\���>��S�~֭���l���!L�8gB���I��9o"!b���$Ve��%��rXO��d��U�k"�H^� R��.rC�$r��}��fH�.��`�������n��Qw۾u�X���*�K�l;����&����҅��U(�@��d7#���g����}��&q�`�|����A��0���Q �Ut�G�d<@.�Y�5�J?�F�5�e?�%�d�xJ?�5|�K�������J�������&Rŉ
�n�S��Vt�8�N�^���f�N����06���a�L�|�0��y8Y$��?PK
    +Q�H\A)#�  �    w/fr$a$a.class  �      �      �U]s�T=�?d�jQ�:��+��.�
��.�N��Lٖ����r>x�����0�dx�?�î�Ԧ1��gtv��g����<���"�H�����, ��3%&��T��Iެd)�\8Ig�+�e������P��ջf<�a;k�Y���I�& [�:n�ы=��s3u��{e������3��������4���-K���me����mk��Zu�zKmk5�f;�ju�[�uͥr�]�窷�r~#ݧ�Ӵ5w]�����H����S�����E$��:������
P���5��ht��ni��jjVS�[��dEe��-:݈�[MwW�9�y�
�m�9,u�6H�T.�8�ڪ�Tnӱ�\���{[F[��Qwh_3{T���b�ޙ�Q���\��������L�.�9��i3".�H�xQ�K".����"^�D�"K�I絝e�/�����K[8�(J�O��~���}�#�ǒ'����E��ˣ����X��(�M���a%�WF3L]Q��LM������	�+�g�!��W'H��'�O���ɲ�V�h�I%U�Œ�81%��2� (�B2�GX�Q�ޑ1�we����<��2�-â+��}�V9�ʉU?`��a-�7�.�
6���-!���HH�c�M	W�|�pK�5|"AEA�/u�a��s�2�6�;_2T��py	o�>���]�Y���'gj�.wz�K�]6�F���,�v5��%�ii�F\�گ�_��(�B�@s�e�}�f)�"+�����韱��G"�"�k����.-����>j��B�qw �w(C�8z�?AoQ��o='�	'�}T��JFL�}|}�a$a�h"HD��h$"�� �1�<;�Ӗb,�`m{�4���)sp�#���B������u>yo��7���F���� � /��7vL饝��P���|�4@w�q�������~뎼&�pH6F�|��W�8K怨J.ҽD���,��PK
    +Q�H�ٖ  �    w/fr$a$b.class  �      �      �S[OA���n����B��d/�E��j�K	��m�͒v���*�͟d�����2�iq1���|�6�;3{f~����<v��c���1��M�+�B� )����vCw��K�Y9�FY/��?}{7g4���uN˚w]^�3+���D��*/R�i[ԱB�I���c4x��L~�Ɖ,lZbϨ{<4>zݰj��Q�7E�|�<���q�b�S;�e����\l�G����U�	�%Op�As��ϲL����
��{�Oz��CR��'��F��M�nJ���Q�
n(QpS���[�� +3�P�R�9O���Y:�eA��x��	2rdZ�Om^α�w���,ÒH�g
�s���d���L>��dw~�����l'/2�iV��¸��WBw%��Џ��0,�����٤EB)�Қ�p�� �"��1/aA�Ccx�b�%,���#����VT�x*!#aY�3	�*f�Ɵ�+t-U�2ʫ��,����
s�d�^_ Qy���@@�<�=�B���m���N%S'XO���e�o�J���l��	��t�wr_!?�]T��!�	#�>y��6޵�km��?Řt��T�$���6dPF�x�fS�бYo�}�ݎ;$��I��Q�?E-D#�&K!=�BA�PK
    +Q�H�QF�N  U    w/fr$a.class  U      N      �W�w���-��z[N�M��M��iJ)v\�!�ZcS�6����:�V�V��gz�Iz��gz�ִH�C�@ ����>A_gvWZ-������7�͹3��ʗ��� �ƿ�h�%�P=A�DTD��Et�x��[ԇ���Ǻ�1�X|�� �zV���S�3Z��2:����Hi3zR��;�kVGR�YS�г��%��_j,[,P�����5��)uF�f�l:�+1�%�>�)�2ATS��㲑�]��j5�1����6�����M͓E�V��&�1�cOҘ��գZ4aꩩ贚�&S�f�ё�m�茦�ɏ�p����0M�B�_S��g���5R˙Z>�����fTr�,��)s�2��B)K2q���M%��%i��C�FV�?�U<M������*ROS4�)����d�@�f�pA��c�,�2�r�	M�:�ݭ��I����'�d����5I�i����cɜNk�&ӛ�G�Zβ����i}�Ѩe�Y��>*Xz&�S͑��h�|	Ӵ�K �9H_(-��v�S�ƜC�5�1�y������Q-3X����m�L,��_�[�i�)d�vMy��U�����l�Mo��
�r�Û�|�b1�p�,G�Ꜩ���E<S�"nq����$�y"6�x��"�q���E�D�PċD��)bD�.�D��ui�m�sm��;B��.Mߝb2X3\�!:m�!WJE�h�n�R��}�����k��؞v�yZ�s�MH����p��;��p,��J�k�>\{�oº��6�����
�畫�*w�6���sTyjsku�^����}����>����q4��E�d����E,��.ª*KqX���	mr���5���f/�r���>]�m�F/_��?��PF����[ֳ�3#���h��~�a�N��v��^c@��j�b����O�1�W��3>	R�}ڊ��F�|����ސZ���Q���w�y�S�N����&�9X#�v�-��Z�X/#���6L�P����:ݘ���pC+�ю��Րeldb��Њ��d�U�c��̚��d6/#K���1�#2�ᨌA�V���~�{%;xSo���I���x��.�E�ux���Z�6��q�bx7�{���>��3|���cd�Ç>��Q	{p\¨_b��� >��E	{Q���`�$�q�y��$�����c^�/H8��0Js�xT�A|��s��&A�W$$pR�N4a_m½�çf��=d��WQ�����e��i_N�m�8���*��g�(V!�]��5B�:����N��wj3��˦Z���,���Ӵh�l�v{�!��-.O�c�4W@s3ύ���x�߉F ��oU"E<����)��D����J�����J�qF�XP�8��EX�=E�S��x��O��G�����J�(���S�׉����+���EO(��h�X��%j�ǟ�@\���WlY���J��N�qZO���;ڎa�)����9��¢2~
���2�W�E
��".�����(Q�Y��TJ���i]5�x��@{�k���Q���*?�X�(ջJ^�'i��u��ߕ�mvP���j��V�j6���A<@�{�ۙU���0kk��!:a�-d�}�0Z)�g�p�q�{�����٫Bpk^�V!�M�G�,\D�D��{a��1:9��x%�H����_h\O��~���\�se�)�=�������CY���<��5%|�:?�X�D٦�ox+^嚶�Φ+8�lU�W���k$*Шwڮ�p�Sx�O����������J���=�|�<{��z����B�C��ɠ�������W��x���Ҭۺn��/A��_�)�f��C�����vI������F������PK
    +Q�H*LKE  �  
  w/fr.class  �      E      �T[s�F�6�Vȍ�@�m�(PzqHKlN�	���-е�Q6c�F��7���8�v��3?��YI$3��ft�\�=��j߽��? _A�1���F��f�	Cj^z2X 垐�V�0�.�`��qr�VKx5zm�n6�v��V͗ζ��6�|aym��v��Z]��Ȧ���s��v5�3�L{X�x+���,v�-.&e�e�*Q�R��9\5�0j�������s�M�Ig��ul4�e@�2
2��q�0��w�U�k�ye�V8u�� ;��	&�M����)�v��_Wy�Z��	�N�`G��7�ڔ^�J3m<�m������䋎��^Z���R��� �����;���0�ᘆ�F4Lj��0�ጆ/4|�ᬆsW͕Ϡ���˄�]9� j�H����J�r8?���O�������2+GD&�������6��04�'��@�7Ch����]2{�����B��TƧ�x(��G�fi	.���xܣ>�t��/��6�F��m�*R4p��n`7���N+q
7d���1|���TEX6o@�-%����m`�:.�'%금��K���=&�ȡ�Ē�XՑGY�e�QbY�%�tp_�T��+5����[��`T<O��:o���5�z\}{�w/S�zRt��fd�b}��s�"���_�XO�]��ų.~��C����.�*l�򻰻�oB�>EI�^D?h�&p~���}�3{x2ֿ��.~�]�������B��G��c��8�Ӫ�ffw�G�&\�ƨD͓��&����C��g�w|��5���2����>M-��F`����:���PK
    +Q�H ���  	  
  w/fs.class  	      �      �TISA�:$2 K�A\A�.�	�@��A�*�I�8fpf�r�*o�՛��!�TY��Qꛉ%�,�����u���?�|Ѝ'�8#���$�:�ᨇ��^�Н>Z$�f���'O�|�fhJ�+���7��h��em����i	Ͱ��d�e�M���r����b�4��E�/mj&�W��%Ś�-Ǳ���'�a3g����C E?CU����c�FfZ,�-mq�8%A���DZ�3���Aэ՜S�GM��v�4�r�C�2_�Z�ѳ��nB�)BŁ���?Pd�L��j	�&�[�!֟2������1�b��Ҵ2� �3�:�L�������Ӎ��ُfS�$ֵ�lAXaDNB�EB��:	�NJ8%�Q�Y	�$��p�AM�7��I����A���f9��:�H��Qm�C�>���1R�&7E�|�l��EF��Q�7��pU�,�����D�umq�3��C/�����b
$h
�(QP	�� 
�\�KA5��pE�i\SP��
TУ�7ȸ��n�ALFn�0,�w\��C��.ܓq#2Z�'�qm�wᾌܕq}e�������%����c�'���t-��j	诊$#h���m�C)��5��e$�|��.f��2��db�c������74E��l��@IOP����u���W���<վ<f��j��዆�P��B�RyL��a����i�CǼ���g��0�2ȶ~nwx��y���
}�u~PK
    +Q�H��G�  �    w/ft$a.class  �            mPMK�@}��S��������<+^z
�^<�5)-%B�o)� �8k+���̛�y3��_� αO���O��l\\�w�I�G�8E7�I2,.s8�)���!OQ� ſEjbńe�nb���1�-f�l�梧�\���r��U}g��q��p	���[�GBYXCK��6���t���βd֝�y���!$���*�@WY����3���˷�F/<.��a'<)�	OK�_���}ͅ�a$�Z����<b�n�i���oրa��0��PK
    +Q�HG;UƑ  R    w/ft$b.class  R      �      �S�R�@�6-MB)�J�4m-��*�Z���0��JӀ��t� �;�C)��� >��٤�
cf��9���mw����� ��VBDB������~6�RSk]j!�^`������{Rf,���bkV�t����&0��z�j�e2J������&1�&�k��wH�,�[�G=g9�eײ��5����Vt{3�T�2"� bY����U)���ʧ�g�4�������K*rv)Qo5��۫�n.�H�f�<'HN���6�i�%��R^`{ɒ��"Ή1,⢈K".�q�a��a�<U*�I�p�#e@M�OI�z�73܎�黢*�i���!|�x��}jV퀟�n|����|������\�ű���唜
�#� ��7��pq9��䎛
zp���ܼ�5܏"�\�e\�C㘑������q�2����=��LoL)ض�.T�Zͬa��`HA@�7��'��e�%�L�(1B��j�}<��\��c�+��x��ڻ��XL����Ij�b�s����Ć�Ƿi�¦�j��IZ�+}��MF���6W��^[�p�7�=����h�,�%�?�uh8�jX��`L�GO|Ó_H�;@!!�QL�J0�:^��g��j�Cr�UL�7��@_������PK
    +Q�H=]��J  �    w/ft$c.class  �      J      �R]o�`~�V`�1����P˗ݦ�}�qE�1Qㅻ*��L,	-�'y�&N�1ޚ�����p����y��>�+��~�`��	�z�@To�v�3zsw����z��z�¤Ӧc��$̷��3�}�I���<�J�zݞa�k8؎g�^�M�2���޳�k�Tе)Fq��e��@���{M�;��7�{EKAB����
�$��Z#m�TL="i�u��:���?5���<�u�\��=�]g��{z�5}T��������0n�<�����g��BAN�.��Bb&�/`2CD����4~И]a��5�l����8���PH ��.@O �[�,�(2\g��p���Pf�0Tj˴�F�C+W��c=�um�T!Z$�4�L��UΒ?����t�H!��+W��Z�����V>��g	�YJ^�����	�"9-�ٲ,�|<���q�{�"�� )Ȑd�㞘J���BX9V�K ��k�ϸ3�+�����z��X�SzZP��Q�ܴ��ؔ��XUED�Oꑪ��Q$L|��W�I�(on�wK��$rZ'E<��~�W;c�Ǜ�!L�c���,�� PK
    +Q�H�����      w/ft$d$a.class        �      �RMo�P�g'q>\��кu8NJZ�!�C{���CsrSR�TJ,��8P��?������B���7;�v��>ۿ���`�
�[���v��vS!�6��#��ޠ�QP>W�똫�`��_�z����vN��P!u^���G$��QFy(y6"e�@�@�@��i`��5�Z��T���3N��������~А��nev6�FL���w�78i�[�N=����F�޲����e����Hc�D
J���)�t[�la�����J�)pK`;�e�.��;w���<p*�@����(��� ���(a���PT�.��_�dl��dh�&�)l_1�f]g,y�1z?P��5�6���Q<�����1�}G�[\���&�5F���zD�	�i��Tj�r�L�Q:<�0�S�h5���*ad_eT��ɼ[f��^�ȉ56_��sjĹ��	�V�Z�S�K��f/S���^$���TU�u|��Ztç�6��(�B6��
?z��D���PK
    +Q�H��o��  A	    w/ft$d.class  A	      �      �V�S[U��fy���@\Z��y�P,h�bXm0P-X���B����R�uA[���:~���4t���Lgt���F����;����Y�Y��N�~�� ��r�JI��g8�V&.%)���Ƣ�.�%�zB3���TZ}��iЊ���5$ wX�T˓�/o�鉔&���mWur�o(N���u���	MS���-~�3�zltK���tj�tt���<�������j)=18ӐL�1=AE8�ʩP'�5Ƥx�f,�n�:<&S�ںA������]0�;\lrc̈���'b��|O�xZ�3"��8 �YE"�qPD1��~�rL儞Hҩ���5�%��,{IQ�Nہ
$�r��M:�tB����YO��)%�v�&O)�B@��e�|wʶX�0Tc��f)f;�A2fw��3�.U�\�:���������4r����)�B��Jlf�ipsVe��>��#�\�Iew���F(>xd�ᕱ�2d�ɐpBF�̐��c�a�PϺ��%,�{d��68XG�$�!�����P�lmb���f�Z�����6D8^^a]����ËJ��p�����/���i�N�.����3�)��m�>�~	/�-	�I��C�a\�1�2�C	��Q�!��N���a�!��k0�@��)5@o�ѴX�)��������L�5U�HǨ�j�F@9<�����y��{����d:w�yl���&h�����D����8E{o������\
�Õ`�f��B�`.���B�w�!S��.�2�%属`����`~�x�̚^�Nr��D���]��1����p�@��i��o��{cy��PYST��!��1��#���(yp�.���Fq�˸~�5Q�8���Ş�?�,��E8;Bk��j���B�}>�9{%?�M'D���h7(���Z���➲=�_���	���)�\�5��o�`�Q֗.�S���|Խd�kn���m�'!��&o�d~�q�r�h5j��^)��i/]���+��z,n_��7�1B��l]�� [��"|�P��/�b?���ao���H���q�&����"{�yIm����ERl!�r�I������_Z��WW���}5"K�"����<<O>���a�U|Cu���D��!�?5��E?�q�b��3�+����B��Bv�-�
�[��.����>�j��~�U�q{�#����Q��v{�PK
    +Q�H-!��   :    w/ft$e.class  :      �       MOMK�@}��IS��~��A�ϊ ��P�P�}�nJJ��dU�_�$���G�/"�]��{ofg�ϯ���
�˫��{����+(!Ē�,de����*��Y�F3��f5�m�o�E�B�:yZl��V�5ɘ�&]h��G�C���C�I��W3[�f}
��9���ziij+�Υx���UZH]�߈��gPQ9�Q��1u�@��9�2�!��t��1ء9
cƀ9b�E�PK
    +Q�H,Z���   �     w/ft$f.class  �       �       ]��
�PF�I�Y���Е�n-��EЦ�UT��W�gk��P�آ����a�y<ow s���	$�����0.�Y��TY���ɩΏ��}�mT$qM0/aʲ�RK@tl�����a�?�r�q�|.i��V*����:���.�2L~�m��v�4<��l�r߸m�~PK
    +Q�H�^�L!  �    w/ft$g.class  �      !      mPMO�@}�kA�á�o&5^��$^8m�m��J�E���<��Q�iЀ���y��fv��?>\��P����1a���Й��$RE���8���YZ���5�xu�'�����p&eB�\�Å	�K�.�h
l
lڶW��u�8�r��5l�,X�y�+��QY⻄���?�C��*r��m�^��o�W>��՗?��wJ�M"�,`j�HI=O��E���
�'���c��#��C���3ˊ��In���S��9��.L�B;�r���sô~ PK
    +Q�H���G�    
  w/ft.class        �      �V�W�֖��z�؊s��-�n,K6&mC�IC��BB�B�:��BV�Z�D���r�p���J!� �2����R%��@B�>K)�������������y3�yo�����g lſ�hrCvc�����&76���F�;x}�6���O}8�ft-�"c�O��Riݗ�g2鬮���8.��eq����EC`r��0 �q����]�Ԅ�k3�/���R�i�TV�V}YEW}3J2�
�ޒMgԬ>���9��մ/��h1�K���D���0_@@G�0'є�vJ1��UԸOIfU%>���+���Uuu�BA��(���"�(=1zX���)z�I��=�#�x�u�=� �����E
��?��(�I%����vOź7�$��#�D~ZM�UNݫ��:QX��R��Մ��\��=�ƨ�MSX�j��h^K�W8:�T�L��I%����k^ג�ԟX>��Z�==�ņGqP�R�ㅟ�'I�4qDLkS�#Iz��1S9]ɒs�XL��3=m&`�7j�l�PL����:DSO�.B��Ȣ/j+1[�ۊ媛�z�b+Q[��J�VT[���GQ4��d+������!"("$bPĐ�W��j[E�!b��{D��z�E���G�D�+�>o�&tм�W�nG��$��C�o���V�wN��9��&��JTU�*+�3rK�W/���ֿ!��ʟ��������S��&�e�8����o�)-Q�ْ��t4앳���Vp�`�a�j׃�Tʨ�y�a�=��(Xe�>T��#�����L��D7�e�N�L�]��C{�*☒�aŌ�-V��↭�\]y[����v���N+���4P9U�7�5*U�9Ui�V���ڽ�������+�f4P���JC�h�p\�'d�0 )�N��:���i�����;d�FF+���b�f�3�3����hfh����9ۡ˸3�$��2|�e�S2nǻ����}l{��l�Ç����}��� �O1|��3�e���O0|��c���C�=�0���K_e���#�z�f�����0/a�&�M�o1|_��D��0|���8+A�9	S�2Óg�b�.��~�?bx��=�8]vk��St��H�t#�{S)5�'��r*�z�Z"��U��S���$��'H�;݅ux+��aҽ�d�F�$9ʽ5$����Ӽ>Yz�s��]U���Nۇ��pQS�K#/��8���,�jPX�e�å`	��"~��u��^$�0�W�-�\@�q�����rx)�Fv�l��V�X�-$�%<��Yk��q�h?�[��dEo��ˡE�T;F7NYN~+�r*]��i����/�h��)�������V��qkJx �uqe��^(!��OE�F��Hp�
���4���s�K�������"�:A��p���
�/�D׋x���^�c�[��0a��0�}����ST�I��\�(5�7f���[=�q�q�:���:hgm�t!z��f^�Z�t��U��9�V������yz��8�l�x]E,3���\)�E�9�k� �-�e�P��?������W��`���9���Oghmy+�Uo�9sΟ�}o&��Ǭ�wP^���u����t6p��:���,�j��u��7�Cq\\ %�H�x��Bd�Y�d����-�#�u��r�R:���t��Y�"�����ъ�~:�XȈ�H���_\�Ѿ��2���"��V�O���N���+�n��y+��$y��i7u��1^���c�4Ј5�i�ؚ���u�f�k�k����=��;�:oy��&���������ǟD�`����l�s����Ac�ϱ�[l� |�6q�%~�8�fĖ�"�V�N�c�n*��ߝFci��qx���G���ֹ�!>��C7u��2���/ٟ�N�	G���5���zv�!F7J�K��,J56Ӎ�\�tmE�,6#Aҏ6#�C�4��$�F���v�ݍ��PK
    +Q�H�����     
  w/fu.class        �       ]O9
�P}�Y�&n7��6�NHHc���!��蹬���O!80��ޛ��y� �1$���`E��*&� sqA!�,X��t��-8M�l6La�'�[)Y+q�Y��f���m�E�Y��oc��h����������J��KjL�0D�����N�s5�`���B�)5�i�h���PK
    +Q�H`&�i  2    w/fv$1.class  2      i      uQMO�@}+�,R��Ib$�.�	ƃ����5m�������h��x�Gg$jt7o�v��������:�1M?gXlڮ�X�`z��]ߘ�Š�̉i8�;4N{#�2��8������3H����	U�M��ԟ���#���Hq,q�G����_���j04�G��P��tt��G�=��;sڜr���	1q!���b-	�BRH��B����7��d�ݾ��;<��Ko� w\��ێV��<����}�T��2�@�@]hY@��G��D�ٱF��R�	�a�R�!O%O�CRD�B��ꬪHMD�t���Fx�v�F�]����~t��Hg�R��!�+�PK
    +Q�H�j�M4  �	  
  w/fv.class  �	      4      }UkS�G~6A�b!EhDl11�,E�� J�c/���`|�&o@z�w{���C�_;�LM;v�L�~����������.��m2�<�=�9������+��rG�G��}��aw��K$y��`��<xT�
���)��p�;�hR�Y�Ḵ�����F����y��xzXZ��d����P���v�R-��e���筼=( hߦT>kCٌ�	�%3D!������gJ%�ʒ2Mc��&��4r4.��Ә���e�+�/�\�p���^2-����d�������9c���&�r��W�Y�˙��/��.��IޢH�Di�E�M��?AQ^�E
��kZ�sJ��H=�̹E��eAx�@�@��>{��k b j`����G�����z@`����[�E�����Ӳmk�"0R���pi�5|�̥R����e��/<΅��q]����Ծ�E�?au�GX��U�|�@��v�Շ�h�>�&�m��&�%)��g734�����a7CC/��8���x�Q��$Kc��8oz���b�b���	�8�+N��1$N1$�8��1��!�&Cы���0N3�x1���8����1\`�3�2\d(0\b��Aڋ'p�!����S�0<����t�F�Y�p�;w�B�[�Y)d*����|���ղI����/�$@�s�~!�׃����4��Fcq�k�h�$s4rfJ�R����U�c���c)e?�yBs"�)V~�hT�z>���:��L��\Ts�����h9���D�����e&bAHe":T&���w��D��H��e¯2�}ڟ�lf�0���Zbz>�6/3-*s�k41v���	�	�?��TED������'�_B���zRsJǩ*%ZT��_UJr�9ض���3~ �C��K�z]��~�W��ԴY��/TMqU�Wx^��I}:L}*���`��0��i�.��.��.Z=��|�O
�:��gڤ𑃀>vP�rq�?މp\w���#�_:�?h�u��u��Uױ�#��#]Ց��.��e,���[�U�T]�-�E�R]�:�U���pUg�*��AV
o8HK�-I)\q�������=?���z�z)�Wz�V𶃎u���W���݅��&ݺV}�7��Ʀm��
^\\�5���n��[���[���͡�9��/Z�^2D�"��Α���|�^ƭ�A�Sn���P�j���������&� �700uG����2�Y����fѿ�^0F�L��Zp�T�%\.a>POBۚ���FV�Q� X��2*���eȂ�y����&z�a��
�
���EO;<x�T��PK
    +Q�H��bf�  c    w/fw$a$a.class  c      �      }S�R�P��M����X�`.�����*�Mo�m�M;i���| ��02����w�b3���~��wvϜ����;�a$exe�e44��b��;��f���#%��D�5\�F��yߘi�θ@ӌ���z���NH@�NA�N��B��H@��%�(��[)ɐ��i9Kzv�h�з�XV�ұ�OI���y�Z:d�c�[����wl�JOn�����dY�I;yw��.�R��5�N-�؅u7�r]ɥKL�n�%�I8+�]B���%\��pI�e	W�(�ңn�^�@N���F��;&�-R��%w�%׭�OHe�������l�H��چ�tjj'�����<���`�rF�N<S�(*�-�:ΡQ���ð�V�R!ç�4$�����&\W��n��m^���U��#�Q�1�{�~�����0� �G
z0��f3<Q�!���
����;�ʧ�9*�����,Þ��ŢQ�Ik��4А4+�,5�3�x(����|��W���W�|�ӿ�7Z�g�'z�xU��W�Gg�G�\�Mu�he,��}�(Z���
�s�8F�Ge<?��f�fs�����˽��F���{�]���`C��]�JPP\�K?�>u2/u&[���&��ꥷ�~�t;� PK
    +Q�H��X�  �    w/fw$a$b.class  �      �      }SkOQ=���vY��*E��>PAP�Z�REY��e�tK��������-��?�8�U��ɜ{�ܙ�w�n�:�`��R�UЬ�@s��V�	���|��O(���@�i�θ@�LA�2���*i
�J�|ް�O�P�R��qy��)ߠ0�r��6I-��=�խ���Ϊ�w̜E���	�1֍�@{MK;�Z��6���)���ɹ;R1�)��]]�:/A�͋n^�\qI���#�M�9�2�dt˸ �G�E��+ɦ�.Y+Q�n?��P8��9InW�R�C���梶��_��@�Q�\�3��i�:U�����{_͞gbi�*9�ǍN|���P5��-�:ФAC?� C\C+5(�5tb�ِ��f�k�n��M���
ƽ��;�cw��bn1�f���Tq_E&���#�R��#z�S�}z��G����,�0��m۰1H�a��xh*�����|>���|�c^��k�F Q-�D˘�DK��{b�X��<�?��ys��t����?z0d2c�2i��K����X.�q	O(��EG���$�i�&rU�Z\R�je]��N�6|J�����4��Ç�]<D��>^�*xō��K.O1�+X�G��;�
���xK���#�4IНGhJЕFq��PK
    +Q�H�֩(�  �    w/fw$a$c.class  �      �      }TmSQ~����Z�o�fT��(jo�f�ZeEi�����.�����ѿh�əj�؏j:�-�tb�>�9Ͻ��{����/_LbKF���.W:=z�c�LOq'��L-)`��B5\�{C��@۬n��@�JA��<E���Q��'�+l��G@P���B��j>��$6i$h0��)��P�\���D��. 놹�fwh]ז�����.�%�����kC���
}-bt#���g�<#�����&k3g�RC�`�`�b-�hm�U+ߵBɒK,��V�$�I8#ᬄ!	�%x$\�pQ�%	�.Sa��g,�*�Ö�n�/��I��W��86�K*k��u����Y�H��斖0knc'=�?���=���xM2g���L.�+�dp3t3�002�CQЁ)�����M���Ӑ��uNo(8���7��6���Ĭ~,;0�{��KL`�A��9����A�	/8�C���c�U'��̉q<t����t?sI����夫��C+,f�bQ+ҲI���3�O��GP�n�.wIy>��oA M�U�(N�G+������m�#�ئ��[ś
���������z��	�ș�cŪ�����xN,ZA�I�U�I� Y�z�V��f��4�2�3.9[���i��0w���!|�}�u�T�ɅU�n��cGx�� ^Ż}��f������7%��3C vA'�n��m�N��PK
    +Q�H@A~��  w    w/fw$a$d.class  w      �      mQMO�@}KB61.�P�WKZ'moA@TE�@E%zr�&rld[�q��T�j�C ?���X�43ov�<��<����>�!%^d��@n��dG@�4O`��uN|O�_���Mx�f����ܠ��_������0�8�����.�!�b�F��}�u>^4m*�t��i�O���)�x	C�����$�%��65�An3%.��Ǿ"���z}�U�R��Tħ����@�<J�?Q8ju)��kD��"ã���8���󼆉q,h�hbK&rX��ky����me�+`/�j`��P5x�A;�O�z\�1z������zn��T(q�²���pK�7\7�D�a����^�ߣVk����,ʰDSW�c�v�� ��Ӱ86��� NZ�%q���x�e%��xV��9
�2G��PK
    +Q�HE� �D  �    w/fw$a$e.class  �      D      uT]se~�f�7	[LK��j��	m�U��Zi���"��@7�7ɖe��v��?��xí̄���^��� �݌�C���9�y�9o�{r&=�m�;�$N
Č�fTU����(W��$�m�V�. �U1�J�2i&1�����Ig��"���a�q���`���Y:���-s�,9��.]1С�'�n�����V�g���
�8�L�-U<wG���3�����C�dE���V-��|j4�c:��vK�oCcu#�Fy�i�����Ɉ�DJbJ�U�9��%ސ��8%qZ�M�c��ް$p�eu��B���ao��C��)%Q����K$Y��%:ej�^on�̀�1�
#�<bD�4ʼ�n���(6~��ې��'7��C�]qL�_���~K�,)�4"�-X怷�2���H�d8�p�!�#�y��3[`x��=q��8���	h:2x_�49�W|��"]�cY�Q|�B��P�*C���p9�K��0��S�ç�4��"��Qc��p������4�a=M��d��p����Y��z�uU7����]ߦ�y�6l�n:j�u���e�X�n�]3��RY<�-�����������W�dx
!�d\ �"o1R���g�_�V1�G��=U�P�>GI���N�=l����j���}���Ԁ���z��S$ę�������dD�5��-\�"n��U�~�?�������ag��I:�������b"�(�2��yꠑMd��Y�x���Fz������x���'���TN��}�����>�{����&�1��4��t^S���$��i�,��i�s�^�%;�3p/��PK
    +Q�H`�=�  �    w/fw$a.class  �      �      mV|g��%��Ŗ���u�6��D��P��$v��8�6��8Y'�Yr����RZf�{4���P(��U�5�%:��*{Cٻ��ww�b����{���}���O�y7��$ٵs'�E��^tx�,/��b��^�y��S���o\��wo�/j-$k�e2*V!��J��A	���� {x�9���y�fd�d�����r��ɤ�ѻ��Ys��w'Ƽ^���jY�͂�ϯ�aVKY�4���rK��FR�Y���ycJ��E=�F��`�=S�)�PA�L�v��d~A�7)�h��H�`$�#F.�5�]P���|�OJhNf�"ߞ|aF3IH���UsZ�M���[$���&�l��TA��/эt�8��F�k�,P�w�NHEcF��P�4m!�s&�z�%����HV˥#��gM#���Z�Fs���6We�4�
�'��@N�R�s�r�͙F��f)�Az���Hh��v�	�R��@ޠԔ�7kQcyJP����"mz?uI�ײs�r/D3bI��h-�XR��P%^z���ś=)�H[�ykY��=4^��%Ur�J&��.�,�2�-�<�˸@�sd<W��e\$�2v��1$c���e��B�Ȉ��+�E2�e�1"c��2^L5��m���M�M��P��b�i�7qx͙���^�������׷�w�\��m�
똄C]9�㝵��R���ճz�D��:#$B�z��A��P�MGk�	f�U��-6=9���%MBB ���ǯ���N���j���8J��ʉKC����WXN*,έ�¾�"	���cs���y�(Ԗ��f҅X�\�~���:J޴�Q���Z4Q��>gH[j����~��W��	��[����%���U�}mg�p��v�Q�sjr����w����{�<z�x8ڊ���x��-[��p!�6�Ɋ�TD�FNE'�*����.\�bC'
*B(�8*+֩؀fV�0�Z�U�d�9f��c��=8�b��Z^Ή��2�e�W0\���1�J��^ž�Q��z���x��~���oax+����w�x&����}h}�Gnb� ���!�nb���V�1|��c�8�Q����1,*x	�)�'��	/EI��P0�/3|E�˰�PfXf��a��_e���k_W�\
u9�8� �O3|��ni|����0ܯPU�1|J��/)�f8Ȑe���M��MH�v��2�E_��|���J��L35J?�
CY�X�_0�Q#���W�)Ct(�X�O� O�<!b��+͎�Ӽ��K�[m��~?�-����"� ����Jx<���c8��Hp3q�?]�A�^\Z�CAW	����p	��Jx�8��>�.�.���FZ}����$�����V���"u��]N�(�����[�X<а����r2�U�&~�R��K�=���ˉ�h�?R����_�O�nX�?C�a!P���J;���@( [,�*����pj�\ĉ�[�p'�ܷ��fi�'l��]�IG���T���{�%|�����]�e���_�D�$n��5&y��7P��mI3iX.e���c�a�e�H��O��
�x0����`�[�N�I�*҃B���-)5-+��	m)���N/R��vq�щʴ�l�������۾���Um���?�����}���&�4�d?�ָ�+�m��Cf�������������x#�]�Sy:<�.���s�ó,54�:��]vq�>��YA:�}&{i���Gv������������?�� �N���â�?�K7�w3E�3�TƏo�	���N������Kż�vj���}>t��>l��SD9�(U��j��Lqt��/��	����:Y6��u��r�l�kרi���:ޏUk|��P�\�G��>�n\J�ZWb��G7�B��������ݫڎ�����5C����P	~h�߅$�����PK
    +Q�H::�  �  
  w/fw.class  �            �Smo�P~./-�n267eȜ�� ��S�-i��&$�>u�]jK���KY4�������� ��<�9����폟_���~	0$5�Ð���CZ;j	(�8��20��5p�&pL�%�|�v�����?|oD���d��O�Vӵ�~s�c�����ٷ�����Sǵ��!�C���=R�D��~'qa�q��@����$cYƊ��2Ve�1.>�`X��b���n`��ɰ����K�9���R9�DcbY����s1��X�f�g�Y�87�����M��ǈE�De�,њI*NTHH����
i
6UpCE7W-Uu��TdQWP���	�%���VPFC���5��/�#xH_��ۜa��{����V�\��jz�]k4�#��e7���SlJ�
C��1۔�(Vk�P<��q��xV
�4ē����zi�W!^|�V�3�c��&(J�z����͙��v?����2��^�?��Ϣ��d):u�y+VZ�H�*ҵ;Q#��"���2�%�ʂ��5��R�PK
    +Q�Hfl  >  
  w/fx.class  >            uTKSA�&YXX��Q�Lx-/���@�CPC2����f!p���腫Z* U�g�Ojo�l�tO=��u�������>�*�M �� f=U8bX�;��fȈN�L.N��i��J�i�1��}W�ȳ�P��)�N8Ʈp&D*�Iװ-����������6#���K3�mlנ��~J�.C5�9�R�!�in�M�PF���V��j��r��]-lo'mKX^l�qSs��)B�rh(��$�9۴	ʯ�bW�嶓8�;Nr��2�,؆�
��!�my�f�V��)5Ev�)xʫ %܈a�v�,��քȨͬ���U��#bԤ��N�$�C�W�3;(@�;��ʨ�Q)�JF���2�d��h�qMF���2n04�W��3�=F4�������3��)n~cK�_g�	/8�gD������π�?�y��9p%1�]GWR��<%k��P>�� S�L>Oo����%�/żz��
����C������o��p�h�(D�
�*$�T4xB�_ETaPE9�hİ�b�WQ�ޒ���#�G���c��TA�1���x�i��PЅ��o����c�w@�]
�q���a�J��rW��Cvq�HX��q�1z)��>4AF�_�e���U@s?aT�u�*I3�GX�����<p�x�vJ�#��q����*v�5���1�����l���&��ء��m���G��X8E�����#ɪ9��T+U(�0X+uU⠛�1�ޢ������:>!B�/X<��	����Fb�����F�� PK
    +Q�Hr�c  s    w/fy$a$a$a.class  s            mRkOA=�];��eQ|�V���V
��P�G!�IH �Ok�m�ԥi�(~�'�@�?����n�VR6�;眹�̝�����/ K���`h�P�t)�{�u���A�phThT⵶���v�z#��l���
�!���AC@��`�ivI�:p��\��빭O�x����H-��[w��x�ܶ�i�qZ#-�J�K��#�ީ	�s5�<��>?��c�Z0�0�H\�HHLJ��$�%�Kܐ�)q�����U�eD��R�<�9-�V�\���IkT���n%S�ָ~A�$���K�ڞ_�x/1H:�9<0p��(.1�pY���;�y,ĐB��#93X��X�,�t$�L��eO⸃�t��*���w����b��t��+I�P�ɽ2�= ���G��zHC�5�����k�+f${��LVY���
��g�ꐬ~�Gfl�I������'fߞ�y�6R�߰���ۦ �:�n���X����m���%q�*ߣ��+�hr��?PK
    +Q�H`��   v    w/fy$a$a.class  v             �W	|�o7��N&$��&e���B��dI`1�$CT�d'aa�vg�����/{h��ƣ� �E<��R�eo{ߵ�m�im��������6�_���{�;���k�~�G`�(B��D��F��EX+�:�D�D��"\*BP�"la�"l�Q�m"�E�.�"��'BD�� ��f^/�8$��U��x� o�-n�ʰ�;M܍��3�%�C*����������@pV�M`5�y��	���ψk��ֻO�3*
B�N-��ElJ�:P">�'��1Ft �H����z�/
%u2nO�)=nhF4ߢ����!#��⭺an�#�A�N�B�t�CzIҢG�Z��>9P�*v�M�Gbf"I�aP2���'=�Z�!R�p;կ9ѷ���4Y��7�d�7m�)���B�ܖv$��>}��E�dS21h&h	*�cT��1����}١�� ��RKS�޴I����4��Ҹ���kG�qO}g�pCWg㞬����a��ggxK��}�֮��|N�C�qv����I��D�I,���+t�cV]��Jz��i�Z ����ڀ��i	���%�m�QԈ�"���Չb�l8n ��Ws">@���lOD㆞D(�!�P�iCCz�|�4�%����` 5����hd_`$Ģ�sfM�."�JF�����f�'����ӂ��+��"�D��i-�
�I=��X�O��Oj��6=:��j�1�:�דV2�]ш���Re�:)"l�Zo����X�G�07�d��1eB����>�y�]c'��IA��>}ȪL����hfç�h�E�}e3E�h,��^S�6��@(��3T���E�Љ�@��3(����m�����m͍��ޤ�����c�Y�YY!ehI#M�#Q�Lj4H4��a-��ۨ99#��$}�,2h��EX$;$e�"i�[�I"#&�-/�Q���Y��f"�°���~�����QK<ZI�L�f%���h�M���	p@�� )�0"�An��*��x� ����K�w�n��O��S�f�Ɇ,s�f��Ld�q�00Yʉ�R�Țg-/Rx�+���.���l_{>�vG��a�n�=[�wzlk!�����򓕛�t���M��o�f�. ��o����[�<k;��2�A�����N��0��d���X���8�K����}��|a��'	��,���`�W������0�/:5̩�~��ų��2��CP'#
[����пii�bZ*���A�SK�JW°>1+��U����+�:6�X�+�-d��9*8�W��X�g�h��Mf=7�gfs$ph�S��֡H�V:X��)î�3���l�d븲}�ma�W�v�(C7�n�L���,� �����I4�A�S24AF����i�he��2Ge��a5��a���v%CC�P#�k���0~��Ge��!g9+����2\�a�ge�O0�9:���]��y����)N�)N��"x�����"×�����5n��s��ߔa|�=�d��a/�>�6�=ˁ�e�;ߕ�~ C��݂1���'�~��2����x����dx��W�f���~��	��$� ���7,��CX)�G����Hp����]�b�eP%����W�0���

"��a�B�r�EK$�.���X(��01(,�e��r	�	�B	�,�=(1�3�g0,�`)+���R�'�2�`�K��?�I� ����1x%8�+%8NdX!�����χ��g�W	�,>����	�;��;%���cv�qI�$9���C>?�G��#:׌tR�
��a@�4�Rx���p�z��0)���61)���V2)m$�Ү(*�C��]_ă��Dz7�`U�I\_u
/�x	C��k�1�f��
��'qMU�I�C��$��g�3��>Q���1�bܜ��˪�2�^�`|S7�Rf�-���g�5������3pW�)�W
�qK�	�ch�ܜn�`�.[�mg�nˏc�q�ǫ�;�9j^/�j�86�	�:�'�����'��#��J�񉷌c؎`�B��OQf�됈c�>��X�2ءҼ���)��AQ��z��L���i�����Tf�%X�\�d��yδ̉�XY���8��8�*�8��x�Mv1u�6ϛi�V��c�9eϔ�Tm���*���a��a��\ �:ŪY�O��㶹<i� �>�v�#U����Ҕ�˃^�<.s�J�~�4��=A�m*�e��L�aSw]��u���Wv��m=N�Wj{�4����)),	�W��ԂƂ����|u~w����zkʏ��L�#p53�<��;(\�9�B�OU�S8d��=�\&����9�@-Ri�\��P)-���j/�!�^i1�c̩k.�͆�����/�P��U%N���J�t�ku����|G�a�.���l=J|޹zS��ڽ)S˸7�fo4�,[�mV'��R�D���ϡ��==	yc�9䥪�����jH�i��ɏ����p�Y� ���2���,��_3x%��ˬݮL��2:�R����j1Y�c�,K1����jۤ0�c��$���&�t�Q�:�?�7�7���f:ￗ�C�I�"�K/y��X�Cp��d�Ct!�*��P�L+��讪9�Z�k3�x`z�6y���Z"��vh����R�V�=��I����O\ݜ4�����y�Мjy^�m��w�8��j��/e��LDs���m'̰s�$Ѭ�Qiʝ�����
SRZ���xT9���;K2�IcV?	L�I�!P����{w�ya�r�-��:�sxXG7�lM����a��G�`��tF�q���uċ���m9��Hm��Ͻ�q��q�)���N�3���j5�4��`Z�����IT��c�b)���"��V|�)��/���KdEveVӺD�K�δ��Z��#�Ў
�L�'����Y����%]�Ϣ��j�l{�Rbk�y��(:B�5�}�����g��p=�Tz���y�1�IЉ�c���xǉ� ��?Ez-��oPK
    +Q�H�rkT�  P    w/fy$a.class  P      �      �R�n�@=Ӧ�5`Ғ 1��:!-�.]P���E%�.�ĉ\EN��G��,H*�� >
q&6T�4��s�3��?�|��}Xt���{Q%�"`a�fpLiQ�ߡtVN��A�������p�D�X�|�=L�Q�}�&�á���ӌ@�]��p�2v痓�i|j���:v aH\��$aJ\�(J�H����j<���<����I�J<���:��߬Xo9�l>cKx�i��<u-�4"�d���N�ͨJ+m���p}Π���m�^#�2�@7�h@Ú���i �[�����n���T���G)W��Re�ӉV���Զu��A�
��k��8��(a��e~2a����t��m�]������g�_Q:��~Q������<f�:r�	�����ajl\ˆ�����v?d����Mf��kgx�Q�؛R�ByN�Q��e��Z�*����F��/�PK
    +Q�H��q      w/fy$b.class        q      �S�R�P]���Q�E� 1�`Ļ���:�#HG}2m5XN:I
��E�����	
��yؗ�u��;;����� ��Y
�)�)�U�aP��ٷIÖIO�n8O�b������x��EE/�����"ָS-9��:g8�����-B�;�5^�N@sN@A�A��p�s%�ap��r,׳V}BJ�ϝM���;�f�ZA�	����U���uxx��4V�۴�7���5e�Y�.�S�ܶ*ۑ[oш�M�U\P1�bX�%�U\a*�t�����!t�4Z(v�.?Og��bǘ!���r��m�/cd�v2����Tg�������i�q���↚1:�WN�n�úq��w�v�ː�"-ȣ�#Icq�c��B�xK��������IA�t�`RG��H�G�E��1
SG?n��tc��F����p�5\�iJ�H�8�я��U��܏��隤KnM8a��D�H�4I�a9ʦ"D�X%�� �HY
E@�������9�������w��
��e��2�����{x�N���un�zg��G��u���?P�}�8�wcU�Xt�a���ɫ�ox<��pL�V�U�%7q�Mq%'�QO9ఓ�,�.ɷ䳘�o��PK
    +Q�H����S  �  
  w/fy.class  �      S      �V���֖�����JHb �d�F$�b7ԇ�HN�����V]Ig��Y��(�4@��Sh��Rh�7�
n)�R�Un�r��3Jgve;`�M~?}3�ͼy3��>��<�,����~Vx�҃�<X���=X+�-�#AZ+�>Ъڸ�Ɲ\�w@U�Yqv�v�Q0��N�-j�lL�GL]��|�nu�rŴf陸e��{������"��`2��;N�՝a	�Ϻ�C=��m�+�ǴѢ981Fy�~	�X���)q�E�SeK/ц�H�P������/��4�r,�S�2��u��/�#�uh{o8�=8�]�Sjx�/�HP9Z	�NY��������{[rː�'A�u��$���`�LFB�V��Z�$,�������V|��u���1�@����M�R^ۯ�R����P�H�bz��"�r!�YF�:��m9��]4��q�{�Z��Z?�S�nB��%���9f
6$���i��V	9tO��e��嶧l�P�ijQ��I�X���4��9R�������9fv�s\zl��mk45R�fNP�����%te2������U��ӵ_*jJ�,ʹ�c<Vq��8%�Ez�yG8df������f�N���Y�ޝ]�r�#ʎ�p��(��Ok��k��/Pme���J�
��l���
\$��^�>��@D`����@��eQ��� Dt�0;��(�E�'��BjS�5:w�[S�z�"��_������4Ό)|E`>�r|3�9�\�{D�|3�fo��w�m�&�i~�v�Ӷr!��K�gF��\c�ϮS��'i_������7u.�� sH8��MzsZ�Թ��k�/2��3n�;bV�q����Lٺ��Q�;�x1������#�|{Tidх]�%�vvQy��)`����������3�60|��b�M_vc
�q���r,Q�ŰK�\�p*�O�y��`*8%���Rp	C�
��>�_�Z1��	W��`5�b�j���FA'���o*8���b�N�`�z/��wn�"�[nc����;��B��^��A�����&���R�N��� Ó2v�>�G~�pX�8$�k���$�e���!��3<��Ï~�pD���~���Ge4bRF
�3<%#��e���d��Y<��S9��_����-f��W�BA7������#�*�:�U�VK0�W�Non���@�?ȺnxH�5�*x����'Q%��
�zґ��?}��
N�YpP{&�(�=���t]���S�3'F��A�Y���&l��`��F4a�,1�=	��/V���#�g��_n�+��j�J/"F"�6�� �� D.?<�_�Zq�~5k���I|IkY|�,�`�>|j���א�����������`��t�38�<��AV�{
�5V�O���XoT��&�Ͻ�U�x >�3Τ����Lb���l����VQ�o�Z��历i\��7L�M�����G��S�����?�E/�$�*x��/���ՙM�'�t;�{���F.����צ��1|R��U�[s��x瀐��F����q��٨�����i�q���r�x�ߦ��������Iz�Z��DW9K�2�I��/PK
    +Q�H�ᗨ3  �    w/fz$a$a.class  �      3      �T�rQ=�`�1A��]Ԩ�G�.j�,J�5�Hp�L���ʓV���V%$e��g?ʲ"h\U�>�t������O ��	b}���!�MQˋڎ�jժ���(С�2k��@��Ɍ5�y˶��F]�"��5'���w��ib&5�ժ�IL��QRQ>��eO 2���4|�.�:n��B%���A��'�r��zf��Q6�1� ���شw���}Y��@W��u�@o�0]J׬r�[CejX���-}���YU��T*5�*���V�Z6l�Td�2���ʂ��8/���!���\9,_XI��H���OG������4U:9���|���ql�╂.�lW�C�N��Q�O�~�)8H�Y�I�l�9Lt��mu��,헊M	l�c���n_��K��޿�8���L"�K��x�.�Ǳ��?��v�+\��.������8����:�˳F�G�~��5�����kspM�6A�a��F�8�pBC/:5삢AE�!�a3Nj����5�qF�V�հ�x,�p�?��l��.1��kn$����FU踮"�+*⸪"�C��ø�$n2�Rя1�k*�SI�6���dl`�)ҿ_m�Lt�iۖ�P��<��(}�A7o�N�'a�\ �a���uxCG� �2e�4�A�L<��|<1��HGr�x�c�bu<\��x2�Jr��zJ�u<Z���K�v��Y�:���џ����<8N-Bf)�0����B�(\O$�~��e�e$r�xYW�S��Ì�<�\���"|f���M2K�i�/8�k��Y�በ_D�&��v3p�A���A���PK
    +Q�H��ew  z    w/fz$a.class  z      w      �W�W��-��Xǎm�1ĉ�Ȓ�h Sr8������Qz�����,�:�Ĝ-	Z
-�r�R7Զǩ[ �r7P���>���ە���/q��~gv�̼y3��[?��s \��8��ċ�x��
�}]!��oV`����$s�B!�}
��1Ѿ�
l�A���C�|�8v)#߫@!ul�Ҧ�`RK%�����v�h�Hp�p���rE#N��¬��)X�%�阖��,ّ�=1�7�L�t�I]!ڤ�QВ�P"�����W��j��^�HL�q�|ۯ�tcJ'C�|�Ӥ�\����7�����pĈ�'�_��K�$v�����ز����Hy�5Ŀ�8�'˪-$�2�t6�[��L����1�9D����p4�g�F:�`mUJ�����y��p:E�6-���H>k��9A�HyU}��qv�*�������I2��6T�CZFA_J��,gd����d!eP��٠1�ISzzR�Z0.K��H	D��L����)#F�߿z'�7e��1=;�'�u���W�\"[:��rY����zzrz��ە��ݖ�tM���I�M�v-gR��{�Y�qSZ���δQ�&9L��{���́����/3	s`�$Ӧx��v��d:5�3�O�E�U�:���x���z^-p��k�	l�#0 p���7	�	
�V ,0$0����#�u«���yun�
�}ot�|M������E-t����_$m��1Zy����Ր�)V���y���9�A���Y�/�~}%�Ui��!�c��Ζ�lj�����r#����7����"Y]�v��V[��W�<������1$�h�Ѿ]j,��̋..���7ڨ��ŷ^SU�][�ojݡ>_�����u��:M�f2�?���W&��"/?"6>�b+_�/��+7�J�2��`W����`��_k�a�R ���ъ��MhR���eX���hUD��vRц�*^����T�EJ�v[v3\�� C#��2�`�����7s]PU�kT�#͐��;T�C�Ur<%�F�U�DA�zL��Gx���^L����*����Vx��Y�*�p���`�=.L�}�2����1���A�>��a7ހϸ�F|֍|э7�K_f��Q|���0�0�e����8���q>�� �G>��i7n�74~�i��2̺�����Pr�@уQ�b�ü0���xȃ1|��a�G���O��C�]�
�o���=j(�ҳ�I-��_�#��x+���~
t���e����R�%�����F���֑�GR�"������=��"�;��E=�;��Y|�?���Y<���c�V��9�k,8�p��,a�,�ݳX:�ѭ�c䋽�ѻ��G�4��K��!;&�?��.�v6�l+�OuX��.��;͊��������.�Fc��>u����n�`	2����GϚՌ���(��-3��Iў�rp��D'����>q��o��c��{�^��ص�kߺ���i��8�tt/@e�e����<~^��0rܮ�yf�����+X�V�밄����8��) cN��!e��.0���@��Q�c7��w�o��ںm�vk�"�����`]s�i� -�Y�R�og�����k�Gi�N�Irw���Nv�'�q�E%��U�{lV�{�E<��X�m�^��`�(�/u ����6�&؅�A�Xįm���ա�+���B�i�ɲƋ�`i<�L̃���E4Yh?A�?�"�⪤��"~���^ķ���p	���g���'����;����Z�'��&��c7��v�D�9r���4�K����3"#nrҚ�mE��Z;X����n�mRGT��G�
w�T8_U����⌕�n�����6�k����F�����p�y�f�	r:�&�6!N�M��PK
    +Q�H���   �  
  w/fz.class  �             �S�n�@=�\6q������KJ�4�(��")�C%�>n�M�*�-�iQ��xI*�� >
1�*H`k��������o�� ���f����o���U�3&(�/�dY����;2z%z�a�P	�+܎���#�Hy.��iv/
����nK;���1*�v�^��*GD^`��ߵ]��dK	���D�[���ݫ?�rW)��D�d[��ݎH�J�NL&�$8L�s�9�8.r�8�9�V�T��C:��(7�r��2jE�1���#���h�{�5}�VsR�8Z���Lg�̍3f�I���9����]:K��~HG�H"a"�e��j₆4VL�p]�7txS{%�򸥡���a��",K�(`Mú�@��	�^����ٚ!��p]Ի"eH�@����7��5�'m�����g��G��cC�+qw����G�"��_���x���sZ�o���@�R8���1��§�J�_��<�0Y��^"�&�
�,R	)�/S!�t�rK0���PK
    +Q�HNqg~  �  	  w/g.class  �            }R]o�P~��R��c�HQ�k;��nS\������U�$�a���x��.f"`\��G߷�L7b�����뜜���� PC+	)���(	H��J a:�Î�i����8�\�0��Z]��C��[�A���c�#d�U'���7H�k/�n��2�A_`������8?��#��	�#/�]O@9
>)�hxVA�P�XTqU�5i+9�z~���������X6/�]�a:��gSR����7���E��r~n<����؉�z�#���+:�
�Aѱ���%�ԑ�-J:r���Z
�1�gX�p4�aj������l�2CU�`K@�{�)�2 	���[=�2�pMbo� A��ܔZR�NWҥ	��b�톜���7<l~��P�̤5#
�vLNa����'Ԙ��V�e�U�A�6����[X����ܠ�	�|L�F�vF�D�1�����k��(Q�lΞ�]c�6ƨ��1�_f�<̟�m�d�S����<�.L���u�'x|��oPK
    +Q�H��#��  ~  
  w/ga.class  ~      �      �T�R�P]�i@(���"��D���V��(U����z�M�$��g�W_x��(3�o�����O�S��vf_V�^�ge'?~}�0��z���82�ٗ5�L��n��q��s9��(ʛ.C�Q���ms�\Y�a���[Y�A�l�l��(��9�B٥D��\%}\(m������ܼ�����Ł��k+Zv\����AeW���ˆp��i���4_`���#$.}A���^&)
%N�Hg�	�tu��z�T,�-��n��Eq��[f�h��s¦�8oJK�X&�-�7m�\�_��;�幂
��(*hUpRA��S
:t*)8�4�JgHǙ������[��U��h��r]���{2�%hRګ�G^��ԇ6��'é�A$���d�ߔ��ګ�J�o�I�8tD�D��՜I:�1��P��&�ȨVC=�hhD�Lug�i�&�A�]Ӡ�7Ő4�Ut!.�=�qGE7�����=H����Ҍ��`4�K�@/�^��r��6dD��Rk��D��!�iV�������y�e��3���
F��ƣd&V!�z�BVvS��|[l5��X�����l�?�ns�k������j�磟1�}]��W�Z��4����`�@��:��u<�!d������6+x��'C�͏���@d6V��+�}x���V~���t`���PK
    +Q�H�5�e  �  
  w/gb.class  �      e      �XkhU>�3sg�;;;3�M��QkI6I��N�$m���6m�Z��¦I�jl��6Ʋ�P
*b��X�HkK�6�C��*�HA�T�bAK��̶��hۅ{�c�9�wϹ��$��>� ��3�4�<��4|e�.�ʪ��4B庪u�KW�T��UlY�A��!7u��Z������!����p��c��օ� �n�|�=�z��a��@��8�Q7�q��nK�>������:����:�&����d�g�|l�B?�����ơ�^%�WKOT��Md��׿w�3�|�i���KG�<��4��m�H�'��~1~�4�\���߆W�հ���5'%P$�J� !AR�
	��@�����[��e޴��Mc��P�K�DИ�AQ@�([C�M6EQ"�&1�Ȧ�L���0���A+�XUˡ���axօ�qXևq����Ll`b#O0�fb��ŵ�]�:,G]�$E%K��"�8xg�1O&��§-�����_���[yS�B�<�THVL��9������\�h�C=	���s��ib�ۖ^S��`VWP!�T��IР�Q�õ��g(�*�Z�HV#Ù6�3N��yq����َ0�p�$Ք���c[Fl*�p=��SY�e�����pIr)|�R�<
G�XR�1
x|Y;��tD�I�3ײ�H��=���p�%�{$^tH<Hb�<I��Y���Kø�\_H�/�$�Y}Q|�}!y��l_x4·��|A=]H����@�+z3��G|��g�>v	}���8�"��D~D1��Ct;[��Ⰽ�6��P>���s���98?\( �I�
8�w-+�E�ꏠm���i�-�fl����3;��^?났��s"��n��Y��_� +��d�ݏ[�gK�K�-�-	Ma�й�ބ&�����L�
�P/����hJ\6��MbG�����9l��6�smn��a�"�m
/��r�XW���o����Z�o 58�jp*�ഈ7üaw�T,����ZM0cl&��X^Xě:թ����q���{��4�Eq�͊i1i�,��ʎ�b&3&���\���8��ji$᰼�ђ�Cj������1^�L�]����JN�w5��f4�w5U_Sͩ��f.��tn�f9������P�*4��Tu����ߟq���#�0֣b�{T���EG���乚�R-(5*U���Q�Ԩv��h�Z����נ1�	�<'T�=��������7 oc J�c�\/��a6F�o*��f��<����1�suV`ܒ�Y�qg���"�����v`��f�
��zY�����{G����=����NF�����ut|�
UY�0G�d�:�&���
��d�O�M��˒�]�鍮3���g���S;�~���?(~�:�m�!j�!FkY�N�n�ki��S�=�E���%�E�9ʻ�W��{��|KC�|S�y8���%P�u]'��Ý������Vk�:��XC����U�iK�L�Y5Ϫ����i��e���6w�Ìm�a��k��̪�P0�Wv!��,���=������]-c�sǭ� �	x�,���y����/PK
    +Q�HŢ��   =  
  w/gc.class  =      �       E��N�@���Z-�P �q�q�q���B�1�j��h
!��f#F��2�Vgq���������
8��(��k�vǾ�1���3Z>��8=R�@���{��w�F�4�$������8
S�3��Iz����,#���E�_x�aj���h,͚I�Y&�w�㾍��1�aP�)Q��iX�S�ؠi�)�'�a$���Cv
TD\D�'��?���8��vo�.�}g���|����H�NS�3���k9�Rw��"O�PK
    +Q�Hܰw|  �  
  w/gd.class  �      |      �W]lU>�3s��v��i�mW���ݲl(q*`]i��R��ԢNiK���+��l0n$�����И�E�MH,�CbD��E�O����/������R�6�s�����|=������ ��J ���@�KַH@����.����Z:w]WK���c���<90<0��RRG��0��!���'Nt�������^�>��h�hi��A	����������#�}=�s�Rc������chCh<FA;����_9?: \/����[_�S9B�߸}��q��$._��}g=I\��>$��x�G3'�&�oqc��$��:�&�ܭ��w��o}�m�����/m��o�į7/o=�!��.��yڲ1�VQ�����Z
�$r)�y�۹�Ѻ����=Yd	A� t>P$>��A�k8T����nx�{���V����
�.�@���s|x�/���#�}�/m�5��� �+8c�� MmZק���ȏ�����B�}!P�F�TN^3-��0%63�1��F��TN�&��ܓF������k~�ʢ��9O��܇��qN������U�)Q�q�*���bwDe$m���Q��b@>kj1Fp�X[�,=���j���gc���F� �IO�5����%Xc�)E��
�_+���~�UO3M��4k��^��ĭcb��my�0௬[��֡.\��Ց�:4�m%���v��C���	����I��\�V$���4Dbrlf
	�j�V�����Hx�MX�%�Î�}����e�FLͮ���L�i����������.e�A)M2w���y��;�7��d��K<���D>�>�
�	wbc�O�hf�jU�Vfh��݂+nƕ��=��
8܌5�^c��Y���,{�G����~O�K�g1)��ʹqX��3؍�E#ʞN�rIV?$�Z@��"	�36�T��e�P�e8��ĥ�k##�ĕ�8����w��ca؎3͙���_��삮[S�i�{WE.�xq>ƿx�Ocٔ�p�i���:d��Zf`#l2�X�Cg1���+�y�r|HcA^N������\ԓ��K@Q�lc�:�z���09�ȏ�����f]����e���Փɐ=�҆��S)m�o�a��t�@���Dz�aD2�,�6�:J��+p�r52|'9�W�!�QD� �B��B�g_ \�V8�XH��%5�'����E����tHS�.j�1[̆�w��iT�t]�F��"�*�Q�&R2(��YR�D�D��h��|*�(��&
��}��Q ���W�L�͑(
�*i����{/����}�����+��Q����Ҧ�JC*j���w*��pd-���r�5-թ��q���>���МC�� ���p�f�PK
    +Q�H�x	�^  �  	  w/h.class  �      ^      e�;S�@���A�,�D��q����}x��P5%�?��J����r<���윳��=ٽ�ϯ�":�SA�Wk	2=߯��,��W	�8���B� � jC�����!4$G�CИa�q��:�����Bh����`��t��5��`�le�K� �(g�N�Li���*�萎�i�e���.
¨L�{T�f�g��8�����'.`�v�k
�i����K�u���Y��`�p��ě
��K�n-����/�x'�Vr�Ȭ����>~ך�*o�#���,Ů��YQ�g�')���_Z�I��0ۺ�&���OJ����e%a�&��Dr5�P�PK
    +Q�H�ݘ  �  	  w/i.class  �            E��VSW���b��Q�yH�"Zgj+X���*jm� 	!�$m���й�
z.~��^@/���n����>�y�w�}N���?镗F�9f丑FN9e��ȇFN����F��72`䬑O�O��iL�����M�|�4���Fp�G�����82�L"9d
�Ff�<R$,d�l��-MgF���v�"Ed)!�@Zʕ��x%?Y��#�;��D*HOS�/�Fy^b��E,`13�w,8�:�K�eǛ�Ǫc�q�1r\��-�%�e����z��AV�bFv�c�#G�N���Jn��eg.-��N�G��&]Ii':�N���H�����b+���N�$v���&������ �K"��q�h�uI� ��a�@F>k�Q�����H\".c��*q����������N� �%��81AL9b��&f�<Q f�"1���RJ��$�S)��fl�<�`�@�T�eK��lq!�e�������$��au2�m�qlw���ޤ�Y{��V�m�۵wj��ޭ��Nk��ާ�_���A�^�Cڇ�����i�i�kwhw���?>/V�����+��r�ܸ�����ĸ+�'�b6�Z~{-���b5�Fg�ȭ0jT�cE���ص~�Fq5�n�Q�h��2w�F���Vq�=�Ɇ���	UL�B��z?�M�b�#��6��Oе�������Bשb�j���!��?{m�	�Sh�m���n�>�v����N���gh���/�6�ϬB���֠m��UL���'� PK
    +Q�HWS1�    	  w/j.class        �      }R[KA=�j�]Ͳ������l�P��Ө�6b���F?�'!�Џ�άEQK��w�|��y{~PAY�)�#�J+s$ j�$�D�hqC�ĭ�tG��ە�wϛ�e
A��P�;�	{-�5H�e������p'l6$lplHڐJa�$�Oc"�)�|�[�"P�xaU`�ǩ��=C�s~��n��ſ*����������n�T�\�;q+q��qm�1��Y,bˆm��IЦu'��7R�����˞6��k�{��z�ZFE�@�J�Z�^�aK�F��]`ߺ��ԏ~��H�ُ1��5L3��9�Ѹ���`���Hz-"̳�$�b�k�3Xe�#��"�ŭ���E��(U�N�v��e����`Ζ�,�;�?a� PK
    +Q�H*�#�    	  w/k.class        �      m�_OA��t�.P�R�
�����JC$&�&��m��)ˬn�>�O$&��P�3[#k�&�s�̽�s;������ �p���|S*�w�i�tI��I@>��D$
,��}5��u�AOs����(	��x�uc�zm�{�_�g��d$�;��1�r�zGg�a$c�1�5�3�7��1�h����Wqq�Ų���� �#�t�/�v}���8�O-�od���y�K�u~{�:��a]i�r���-qؚ�ä�a�m�[�����<2F����S��~��.�Gj�}�;�.+-����n�*i_K	̶�@�zXG�m�"���a�4�����_�wS�B?����)�I_H���sS���/L���_���E?���\?�M�%d/&V��kE[��U���s���0^R���߂u<0�C����Պ��m�k����-�ax���������}K>�~DL���3��Z�����Oj&C?� PK
    +Q�H2�=@  M  	  w/l.class  M      @      m�KK�@��4����6Z����]�D
�B7�&�P��	����\��(�ND��9'����������>ZN�3c�J%����I��椐$�K��~��¿�b��8Y�A"å?�I:�ߠ��QJ=Γ9�c�r�cyE%���g��X*-�C��*Wʿ�"
i�k[��x��=xV۷�{�D��T�3vTB��N��qH�6�S�壘ɕ"q�T����Z1�r��N��(�:� ���2�G*��CQ����Rl���kU�m��A21��eOt�����2|H2أ=r��n�y��g_5��:�>PK
    +Q�H���  o  	  w/m.class  o            m��n1��ݜ���RH	�n[
9 Kř��4��*�J���&Y�C⅍7�w�W���x(�?D-p������?}�AD��R�S�teRI�#H�C>ԅzP
�w� zIh(�0���7���{�=���C

�h�u#�z�:�{�o�G�A��bh*(=�G1�u>{c�Jl�m��aK���2lY�[��e�e���[�-�V`s)M����3Y:����Vڧ�&�JQ]�c�W�kF�l�%�Q�[���h�6m�X��˖��X*��Q�߾'�ۖ�F�mo>��t��V��}zƆ�j�}4~���������6VZ������(h*j_K	�?���8
h�`�"��N��3�5p�`�1x�5�8g�M��ep��
x��*x��x��[���^6��3�.F+��	?��*F����O���H��$��?EkE[�EX�%�.�%[b�-q�-���"��&R��O�zBϿ&o��O�fr�FD�j��N�NhwV3kL��7PK
    +Q�HZP>�_  �  	  w/n.class  �      _      mQ�JA��&��ķ��~��x�D�@.�f�u����:���I��(�f�(��������{>>_���@�i��N�V�% �D���O��DH�	���"�C��}#P����5z]��}�m�e���y�þ�$,,9���J.�.�\�,v~��Z{*�Mvi�2�b�M�4��y�M��;�ܓ����N� �k*(@XZ+c�6���U�c�`�6�Ѡ��Tu�ԃ��L��H��$0�U��&Ml��k�qj�Kص;�,�_�On�1����m&
��b"Ϙ����$���EJ%Ϩٍdء5����G/�z�ߜ٫��k�Z�����7,�`{�����|PK
    +Q�Hf�ѽ�  0  	  w/o.class  0      �      mR�J�@�mZ����U��{/J�EPAP
�����mc�R7����SA����T����gg2K&����
`{N�P�(�́�8%j�$D�hqM��B�����nW�{��xM#���T���L�k�/"q/�=�8���|�"l�����%����%1��T3��o�_i�e���Rk�0�c����-�o�w�T�����x��2���lR�(��7�P���������B}1[6RX-��c���Ə}}g�6�A��=mԭWWw������4�"���jkiz��5,�Ha	f.P��#�y��<�9�����6�K�G�s��)f�RX�d7���,W��4V��
⌞��F�X��("�6��"�6E��C���W�W�>v�e�u����K���4���> PK
    +Q�H^ȁO  r  	  w/p.class  r      O      mQ[KA=㪛�J3���=yyX|V�a�H�Yw��m6�Y�]=	A��~T��J�眙9�e��ϯ� }\1�Δ!?R�8�%��g�,����s��]�3�`���v#�-쉊��1r+Ĕc�����&�)��Д5Q0Q4Qf�9���C!��N������Λ���u�ȴ�)��4��ٞ*���{N��Զ3-#��QD'�N�7�G��x��O�T,���R��+�%Ca"撫8���!�9P&=�%�J��4�.I.��#ɧ�$f�Q!�A�.�ҿ��퀪(�Y�dE��q���4��	ڶ�I�����8X�|����PK
    +Q�Hʃ��X  f  	  w/q.class  f      X      mQ�JQ]G'/�fN�݇����"TE�/>��A�Lgh<~VOBP�GE����3�/�������z� �D�!Y��Rm!��0�.'sɆ�	�s��rl߻o�� �n(F����P�Ɯ�3�$_��$�C;�]���˛0Ml��0���C ���C�O�Ki_�!_��o�珨~���v�K_/���Ϫƌ�O�����#n3��n8����~	0�3(�H�c���`D�*?ΤO^_L��{WR�+�)C�'ƒ�Y衂=j��NI�B��)PV"$�E�:��a�2#jѤ,�R�B�T6��jdg�0�K��F�O�z��-OP���w�8]qV���oPK
    +Q�H���G}  �  	  w/r.class  �      }      mR�JA=㦦�����[Yn^,^+AA!	�t5��2b���F�Օ��P�7�a�,�sf眙��f>��> �`3X�͐h)��&p�K����H��=>�N�K߹u{^G1��w�Pt{NK�Î�1�#��Z��	-�MLSL��iNS\S"��cH"��BK����w�����_�\J�<��a�Jx�.͗���h�r���
C9��d<4��"���F�in�����i�O��M�s�A��W�J%�����K(�D ���%W��C	���;ZI�f8���a��$q��%I��\tc�d�d���L�I[tĊ�}�F�uMyl���
��)��F�JN�8z�����.P�i��j�cc��$3�T�PK
    +Q�H��VMM  D  	  w/s.class  D      M      mQ[KA�F]����]�!�����B���O����6����I����3ka��˜��̜��|}��C��3�{B
�g`C2N�0|�-�˹u�,ܩb����r1[X#�S�+�.�=[�$iC;f`�2&�&LY����x��Tn�e���r)�A�uL�V�ތ�W�Uz���k�v�ī6b��7〉��������YP�渀�v��q�]�!u��hF��P*���R8�;��W\	_.�#1�\���K��R(Q<�v�8�X��LHf�t2�C�2���"R��7)�hc8%�e�����%�%W�4\%��\��|��'[��
5�PK
    +Q�HS^#�U  i  	  w/t.class  i      U      mQMO�@}�
��*~�C�BBLL0M4�pᴅ�YR�I�b�Y�HL�����E��6yo�3ofvg?>_�t�`�6[�\_H�lD��0c(-�����}�.��b��ȷ�H��XE�L�$�b�Z>�*K���i��|u��]���mt
����P��R��(��)��s�7�w�;�C�(�S�I�mO߾���:��h�i;N�NhlkRDL�Ie�j:cع紫�C,�x�&b)��J*�D(����%Wq䡁C*��ʄ��o�l��%���(�ɡB���!`%�c��8�����	.IVN<�h�q����N�j��h`�l��ɾ����F��T� PK
    +Q�H�5Og0    	  w/u.class        0      m�KK�@��m��>�Vm���]��uJA�PP,t�j�eJ�@:���UA����DD�,�9�{o�$��� ��$8�ޜP)�̘@�`�+$4Vb#�H�w����q��D�+of�ta~@i#�T��g/u��F�
�;.*.j���w��ڻU2
}����c��L|�d/<N�o��sjG�i����{�(����h���	�x�|��C��z�s�VA$����0*�kBe��Z�4����Ep'_�p�O5�CVu�:G)�r�������g���	(����O��#��m�Q���[�~�\�_�_PK
    +Q�H�̖��  )  	  w/v.class  )      �      m�koA��p�B��j��^{㢮xW�ML��h$ዟXqp;��,՟�&&��Q��l�	y�ógfOv~�����Z�RP�V*t�V�+H�>�`F`�L���TPu*��������`dp�#�!� ������8���?�� 3��0���0��=�6�|\_��,�N�#Ñ��q�9
�G��ı�Q�p,q,sT=Z�hգk�V{�v+��_� ��5��&R�q��Ww5��N�&]�r��4{������L�Kt��r`3��h��T�#=3R��ɬ��&ڨ�`�fj{ZGF�E��}5��$q@� ?C��O���GI����[p��m���;����5���ux���by�d�Mx��[��o��X���Z~~��|�������~1R�!_�ۃ�\9�(]�M�K���eWc媫��r���E�p5j���ꢵ�~áhS����p�'���hfнczv�f/}�'D PK
    +Q�H�V�f#  �  	  w/w.class  �      #      mPMK�@�mLcc�Vm��x��!��RA(�x�$K�7�n��� ��G�o#�H3�-��1o?>_��q�`���D*��lF���3t�|����Կ��"�^^�~T�d��uQ��G��<+������3�p�8�u�2��_?Wʿ�"KZ��#<�RiQ&۠Nx
��f�5��QX�8������c���vn�.9,���b!W2�čR��Z�j�К�Tq]����KΊ/�G�Kh֮ͪ�T�u¾�U�R�ԭ:�nq�b>���F�hG��;Yo8���{��|>N�/PK
    +Q�H1L��  4  	  w/x.class  4            mS]oA�����V�Z*j+�V��+~+ؤm4iC��K�Xqp;[���>��|21���2��;���{Ͻ������??~Q��9�J[P���2�bh� ]�x�{�| 0��c��R��ם��5(|��@ ��}����m�p�5��G�' ��R��a/�{����$�LS�)Ŕf�a�1}	�E�R4~J:���]��<;ś@i�uAy��R_�w�-Y5�����4��Jy~���ͳ����_�s�%�qМn��x�f���m�=���Y��#�ǂ��A�^���Hm���ߎ�Q�^[U�����4
&A�-��ҌB��/O��QԠ5��5����;���|c����*t��%�K_����謥7��,}z�ҷ�,}���yr��[����C�!�.�a!�>t�Fd�E�ed�+�rr@b���.���UV
q�w9n��%JN7��q�u�������2|/���ɷ���}���b1�Yu~<OǞ��|H/���/PK
    +Q�H��^�:  7  	  w/y.class  7      :      m�KK�@��4mcj��Z���X��S
"��b�W�f(S�	���?�UA����DD�Y�s�{g�e>>_��q��;S��@*��lD⤀4#�$�P[�5�"���]�3�Ќ��$2\x��3�
k���<y��c�XΘc,�������ĕ�n��B�.h���TZ$���c���#f�}K�7���������2��2v̐��Cک��*-�b*W2�ĵR��Z�j�P�ȹ�:M�p@m@�I�3��_��A���MQ�����R�6P�ز��Y$��z�ECu78y1��&��&���,w{��68���0�#�PK
    +Q�H�t>*�  G  	  w/z.class  G      �      mR�JA=�M�c�n���?͏���`�P-rӫI���YY'
��+y%� >��̆�`g�s�|s���=�����]|�j��@���2�␐D��}""~�P�P�2�2���_�èg8}B�A��n����Ȥ����P����y��/ǃ������Y�[*X*Z�-U<�O�}<�1�cA`��o�o��&J�'f����}�/���j_�g{�4��c-M�e�h?���w���j��ap�z�����VQ�T�$}�4{��s#��C�~i�N��:W�8��ub�Ql�>R-�(����*�*��<�ض�"`]��_�.N�/X�����z��u��?�"e�e���xI�q�(e�Q�̺�%�s������O�)ח+6�[��oY��+{3{��v�5r�R�����5����?PK
     .Q�H               META-INF/services/PK
    -Q�H���!        META-INF/services/module.Server                ��O)�IՋ700� PK
     +Q�H                      �A    ACvqqLVUSwkYm/PK
     +Q�H            (          �A,   ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/PK
     +Q�H            	         �Ar   META-INF/��  PK
     +Q�H                      �A�   _004_/PK
     +Q�H                      �A�   com/PK
     +Q�H            
          �A�   com/smaxe/PK
     +Q�H                      �A  com/smaxe/bridj/PK
     +Q�H                      �A9  com/smaxe/bridj/linux/PK
     +Q�H                      �Am  com/smaxe/bridj/linux/lib/PK
     +Q�H                      �A�  com/smaxe/bridj/mac/PK
     +Q�H                      �A�  com/smaxe/bridj/mac/core/PK
     +Q�H                      �A  com/smaxe/bridj/mac/core/ns/PK
     +Q�H                      �AH  com/smaxe/bridj/mac/core/qt/PK
     +Q�H                      �A�  com/smaxe/bridj/mac/delegate/PK
     +Q�H                      �A�  com/smaxe/bridj/mac/lib/PK
     +Q�H                      �A�  com/smaxe/bridj/win/PK
     +Q�H                      �A%  com/smaxe/bridj/win/lib/PK
     +Q�H                      �A[  com/smaxe/uv/PK
     +Q�H                      �A�  com/smaxe/uv/media/PK
     +Q�H                      �A�  com/smaxe/uv/media/core/PK
     +Q�H                      �A�  com/smaxe/uv/media/java/PK
     +Q�H                      �A#  com/smaxe/uv/media/java/swing/PK
     +Q�H                      �A_  com/smaxe/uv/media/java/video/PK
     +Q�H                      �A�  com/smaxe/uv/na/PK
     +Q�H                      �A�  com/smaxe/uv/na/lib/PK
     +Q�H                      �A�  com/smaxe/uv/na/webcam/PK
     +Q�H                      �A0  module/PK
     +Q�H                      �AU  net/PK
     +Q�H            	          �Aw  net/java/PK
     +Q�H                      �A�  net/java/sip/PK
     +Q�H                      �A�  net/java/sip/communicator/PK
     +Q�H                      �A  net/java/sip/communicator/impl/PK
     +Q�H            (          �A>  net/java/sip/communicator/impl/neomedia/PK
     +Q�H            3          �A�  net/java/sip/communicator/impl/neomedia/directshow/PK
     +Q�H                      �A�  org/PK
     +Q�H            
          �A�  org/bridj/PK
     +Q�H                      �A  org/bridj/ann/PK
     +Q�H                      �AK  org/bridj/cpp/PK
     +Q�H                      �Aw  org/bridj/cpp/com/PK
     +Q�H                      �A�  org/bridj/demangling/PK
     +Q�H                      �A�  org/bridj/dyncall/PK
     +Q�H                      �A
  org/bridj/func/PK
     +Q�H                      �A7  org/bridj/jawt/PK
     +Q�H                      �Ad  org/bridj/lib/PK
     +Q�H                      �A�  org/bridj/lib/darwin_universal/PK
     +Q�H                      �A�  org/bridj/lib/linux_armhf/PK
     +Q�H                      �A	  org/bridj/lib/linux_x64/PK
     +Q�H                      �A;	  org/bridj/lib/linux_x86/PK
     +Q�H                      �Aq	  org/bridj/lib/sunos_x64/PK
     +Q�H                      �A�	  org/bridj/lib/sunos_x86/PK
     +Q�H                      �A�	  org/bridj/lib/win32/PK
     +Q�H                      �A
  org/bridj/lib/win64/PK
     +Q�H                      �AA
  org/bridj/objc/PK
     +Q�H                      �An
  org/bridj/relocated/PK
     +Q�H                      �A�
  org/bridj/relocated/org/PK
     +Q�H            "          �A�
  org/bridj/relocated/org/objectweb/PK
     +Q�H            &          �A  org/bridj/relocated/org/objectweb/asm/PK
     +Q�H            0          �AZ  org/bridj/relocated/org/objectweb/asm/signature/PK
     +Q�H                      �A�  org/bridj/util/PK
     +Q�H                      �A�  w/PK
    +Q�Hc=��  ]  1           ���  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/AUX.classPK
    +Q�Hܧ��!  y  1           ��9  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/AUx.classPK
    +Q�H�:�k]  (  1           ���  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/AuX.classPK
    +Q�H�]O�*  �  1           ��}  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/Aux.classPK
    +Q�HqpCo'  �  2           ��
  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/COM1.classPK
    +Q�H�H?�  Y  1           ���  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/CON.classPK
    +Q�H�9��a  -  2           ��  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/COm2.classPK
    +Q�H}w���  �  1           ���  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/COn.classPK
    +Q�H�}"�*  �  2           ���!  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/CoM1.classPK
    +Q�H�����  ^  1           ��v#  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/CoN.classPK
    +Q�H�w\�i  �  2           ���&  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/Com2.classPK
    +Q�Hb��K(  �  2           ���)  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/Com3.classPK
    +Q�HS	R��  2  1           ��,  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/Con.classPK
    +Q�HmzK|Q  �  1           ���-  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/NUL.classPK
    +Q�HCQ�$  �  1           ���1  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/NUl.classPK
    +Q�HQ#\Y�  
  1           ��24  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/NuL.classPK
    +Q�H�u���  �  1           ��B9  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/Nul.classPK
    +Q�HB\�%�  I  1           ���;  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/PRN.classPK
    +Q�H�Yq�  �  1           ���>  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/PrN.classPK
    +Q�H�b�Y�    1           ���B  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/Prn.classPK
    +Q�H�ms�'  �  1           ��F  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/aUX.classPK
    +Q�H�9_+a  z  1           ���H  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/aUx.classPK
    +Q�H���  �  1           ��RK  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/auX.classPK
    +Q�H.�גy  �  1           ���N  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/aux.classPK
    +Q�H�eN�  U  1           ��eP  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/cON.classPK
    +Q�H���9'  }  2           ��PS  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/cOm1.classPK
    +Q�HO:��)  �  2           ���U  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/cOm3.classPK
    +Q�H� �  u  1           ��hX  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/cOn.classPK
    +Q�Hϐ�=#  �  2           ���Z  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/coM1.classPK
    +Q�H��ߤm  �  2           ��n]  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/coM2.classPK
    +Q�H�B)  �  1           ��?a  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/coN.classPK
    +Q�Hw��  

  2           ���c  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/com1.classPK
    +Q�HA�  5  2           ���h  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/com3.classPK
    +Q�HִLn�  �  1           ���k  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/con.classPK
    +Q�H@���  �  1           ��o  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/nUL.classPK
    +Q�HL��}�  �  1           ���q  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/nUl.classPK
    +Q�HR����  0  1           ���s  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/nuL.classPK
    +Q�H�W�  �  1           ���v  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/nul.classPK
    +Q�H��7�  5  1           ��_y  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/pRN.classPK
    +Q�H����  t  1           ��U{  ACvqqLVUSwkYm/qjoNcDwEuTGzEptsMFEywgGCK/prn.classPK
    +Q�Hq�l�  J
             ��Y~  ExNativeAccessWebcam.classPK
    +Q�H�~��  �	             ��G�  _004_/SendCapture.classPK
    +Q�Hh��aj  5             ��m�  _004_/WebCamCapture.classPK
    +Q�H=�;/Q  K             ��"�  a.classPK
    +Q�H���  r  -           ����  com/smaxe/bridj/linux/lib/VideoForLinux.classPK
    +Q�H��\�+  �  )           ��"�  com/smaxe/bridj/mac/core/ns/NSArray.classPK
    +Q�H*}b�$    3           ����  com/smaxe/bridj/mac/core/ns/NSAutoreleasePool.classPK
    +Q�HicK�  �  (           ��1�  com/smaxe/bridj/mac/core/ns/NSData.classPK
    +Q�HSہ  �  .           ����  com/smaxe/bridj/mac/core/ns/NSDictionary.classPK
    +Q�H��@�     )           ���  com/smaxe/bridj/mac/core/ns/NSError.classPK
    +Q�H�U`�  �  )           ��6�  com/smaxe/bridj/mac/core/ns/NSEvent.classPK
    +Q�H�:X=  P  )           ���  com/smaxe/bridj/mac/core/ns/NSImage.classPK
    +Q�H�_��  5  5           ����  com/smaxe/bridj/mac/core/ns/NSMutableDictionary.classPK
    +Q�HR��  �  *           ����  com/smaxe/bridj/mac/core/ns/NSNumber.classPK
    +Q�H���;  �  *           ��(�  com/smaxe/bridj/mac/core/ns/NSObject.classPK
    +Q�H,5-4�  ,  6           ����  com/smaxe/bridj/mac/core/ns/NSRunningApplication.classPK
    +Q�H����  �  *           ����  com/smaxe/bridj/mac/core/ns/NSString.classPK
    +Q�H]QToo  �  -           ����  com/smaxe/bridj/mac/core/ns/NSWorkspace.classPK
    +Q�H^�9_  �  5           ��z�  com/smaxe/bridj/mac/core/qt/QTCaptureConnection.classPK
    +Q�H9�#��  �  B           ���  com/smaxe/bridj/mac/core/qt/QTCaptureDecompressedVideoOutput.classPK
    +Q�Hf�ےp     1           ���  com/smaxe/bridj/mac/core/qt/QTCaptureDevice.classPK
    +Q�Hb�:��  T  6           ���  com/smaxe/bridj/mac/core/qt/QTCaptureDeviceInput.classPK
    +Q�H6�\��   $  0           ��Ӷ  com/smaxe/bridj/mac/core/qt/QTCaptureInput.classPK
    +Q�HV�@5�   %  1           ���  com/smaxe/bridj/mac/core/qt/QTCaptureOutput.classPK
    +Q�HC$���    2           ��5�  com/smaxe/bridj/mac/core/qt/QTCaptureSession.classPK
    +Q�H?��~  P  5           ����  com/smaxe/bridj/mac/core/qt/QTFormatDescription.classPK
    +Q�Hb�� I  M  0           ��x�  com/smaxe/bridj/mac/core/qt/QTSampleBuffer.classPK
    +Q�H
5;�  �  K           ��#�  com/smaxe/bridj/mac/delegate/QTCaptureDecompressedVideoOutputDelegate.classPK
    +Q�H1�捥  �  ,           ��R�  com/smaxe/bridj/mac/lib/CoreFoundation.classPK
    +Q�Ha���  R  &           ��U�  com/smaxe/bridj/win/lib/Avicap32.classPK
    +Q�H��>��  �  -           ��v�  com/smaxe/bridj/win/lib/MediaFoundation.classPK
    +Q�H��хN    5           ����  com/smaxe/bridj/win/lib/MediaFoundationPlatform.classPK
    +Q�HdU=�  �  6           ��W�  com/smaxe/bridj/win/lib/MediaFoundationReadWrite.classPK
    +Q�H�ا}�  .  $           ��I�  com/smaxe/bridj/win/lib/User32.classPK
    +Q�HRA�3/    (           ��W�  com/smaxe/uv/media/core/VideoFrame.classPK
    +Q�H��͘�    A           ����  com/smaxe/uv/media/java/swing/JVideoScreen$AnimationOverlay.classPK
    +Q�H3��S  <  =           ��"�  com/smaxe/uv/media/java/swing/JVideoScreen$ImageOverlay.classPK
    +Q�H�,���  �"  0           ����  com/smaxe/uv/media/java/swing/JVideoScreen.classPK
    +Q�Hf�i5  �  5           ��,�  com/smaxe/uv/media/java/video/VideoFrameFactory.classPK
    +Q�H¶t��  �
  #           ����  com/smaxe/uv/na/WebcamFactory.classPK
    +Q�Hiv[�  V             ����  com/smaxe/uv/na/lib/Lib.classPK
    +Q�H��:1�                ��� com/smaxe/uv/na/lib/jitsia32.dllPK
    +Q�H5ߨjE�   R             ��?� com/smaxe/uv/na/lib/jitsia64.dllPK
    +Q�H���$  �  0           ���+ com/smaxe/uv/na/webcam/IWebcam$FrameFormat.classPK
    +Q�H�>eޣ   �   .           ��\. com/smaxe/uv/na/webcam/IWebcam$IListener.classPK
    +Q�H �#�x    $           ��_/ com/smaxe/uv/na/webcam/IWebcam.classPK
    +Q�H����   �  ;           ��-1 com/smaxe/uv/na/webcam/ScreenWebcam$ScreenFrameFormat.classPK
    +Q�H͂���  �  +           ���2 com/smaxe/uv/na/webcam/ScreenWebcam$a.classPK
    +Q�H<S��'  ~  )           ��5 com/smaxe/uv/na/webcam/ScreenWebcam.classPK
    +Q�Hy�{  �             ��< module/_004_.classPK
    +Q�H��Y��   ^  X           ���= net/java/sip/communicator/impl/neomedia/directshow/DSCaptureDevice$GrabberDelegate.classPK
    +Q�H�MA��  �  H           ��0? net/java/sip/communicator/impl/neomedia/directshow/DSCaptureDevice.classPK
    +Q�HC�L  �  A           ��+B net/java/sip/communicator/impl/neomedia/directshow/DSFormat.classPK
    +Q�H����y    B           ���E net/java/sip/communicator/impl/neomedia/directshow/DSManager.classPK
    +Q�H�J ��  �  $           ���I org/bridj/AbstractBridJRuntime.classPK
    +Q�H���R�  N              ���P org/bridj/AbstractIntegral.classPK
    +Q�H�R&��               ���T org/bridj/BridJ$1.classPK
    +Q�H��|�J  b  !           ��W org/bridj/BridJ$CastingType.classPK
    +Q�H9���
  D             ���Y org/bridj/BridJ$Switch.classPK
    +Q�H�\��>  ��             ���d org/bridj/BridJ.classPK
    +Q�H�'��Q  �  %           ���� org/bridj/BridJRuntime$TypeInfo.classPK
    +Q�HX`+Vx  �             ��-� org/bridj/BridJRuntime.classPK
    +Q�Hj�s�  L             ��� org/bridj/CLong.classPK
    +Q�H��뚞  �             ��ܪ org/bridj/CRuntime$1.classPK
    +Q�H��T�  #  "           ��Ʈ org/bridj/CRuntime$CTypeInfo.classPK
    +Q�H<l��  �  .           ���� org/bridj/CRuntime$MethodCallInfoBuilder.classPK
    +Q�H�ۃ�A"  �M             ���� org/bridj/CRuntime.classPK
    +Q�Hן�l�    ,           ��*� org/bridj/CallIO$GenericPointerHandler.classPK
    +Q�H*�|H+  S  *           ��� org/bridj/CallIO$NativeObjectHandler.classPK
    +Q�H�#��  H  %           ���� org/bridj/CallIO$TypedPointerIO.classPK
    +Q�H"BY"  �             ��� org/bridj/CallIO$Utils$1.classPK
    +Q�H��)6�  �             ��t� org/bridj/CallIO$Utils.classPK
    +Q�H���  �             ��L� org/bridj/CallIO.classPK
    +Q�H�$l�  B             ���� org/bridj/Callback.classPK
    +Q�H��;z}   �   !           ���� org/bridj/CallbackInterface.classPK
    +Q�H(�7�  q  +           ��R� org/bridj/CallbackNativeImplementer$1.classPK
    +Q�H���&  �&  )           ��7� org/bridj/CallbackNativeImplementer.classPK
    +Q�H|O�+  �
  "           ���
 org/bridj/CommonPointerIOs$1.classPK
    +Q�H)���  �  #           ��7 org/bridj/CommonPointerIOs$10.classPK
    +Q�Hi���  �  #           �� org/bridj/CommonPointerIOs$11.classPK
    +Q�H[��a0  l
  "           ��r org/bridj/CommonPointerIOs$2.classPK
    +Q�Hh�g21  �
  "           ��� org/bridj/CommonPointerIOs$3.classPK
    +Q�H��/�)  _
  "           ��{ org/bridj/CommonPointerIOs$4.classPK
    +Q�H	�zZ�  N  "           ���# org/bridj/CommonPointerIOs$5.classPK
    +Q�Hj�z�9  �
  "           ��) org/bridj/CommonPointerIOs$6.classPK
    +Q�H?c\�9  �
  "           ���- org/bridj/CommonPointerIOs$7.classPK
    +Q�H2u�4  �
  "           ��!2 org/bridj/CommonPointerIOs$8.classPK
    +Q�HD���  �  "           ���6 org/bridj/CommonPointerIOs$9.classPK
    +Q�H��&��  H  2           ��
: org/bridj/CommonPointerIOs$CallbackPointerIO.classPK
    +Q�H@�2^  �  7           ��> org/bridj/CommonPointerIOs$IntValuedEnumPointerIO.classPK
    +Q�H�nC�  d  6           ���A org/bridj/CommonPointerIOs$NativeObjectPointerIO.classPK
    +Q�H���U  �  /           ��MG org/bridj/CommonPointerIOs$PointerArrayIO.classPK
    +Q�H����  	  1           ���M org/bridj/CommonPointerIOs$PointerPointerIO.classPK
    +Q�HݓZ�0  �  0           ���Q org/bridj/CommonPointerIOs$StructPointerIO.classPK
    +Q�HW���c  O  6           ��ET org/bridj/CommonPointerIOs$TypedPointerPointerIO.classPK
    +Q�H>^�N�  v              ��Z org/bridj/CommonPointerIOs.classPK
    +Q�Hkt���  �             ���^ org/bridj/ComplexDouble.classPK
    +Q�H8Z�  7  #           �� a org/bridj/DefaultNativeList$1.classPK
    +Q�H���[0  �  !           ��Mc org/bridj/DefaultNativeList.classPK
    +Q�H92x�  �             ���p org/bridj/DefaultPointer.classPK
    +Q�H��qM�                ��$r org/bridj/DynamicCallback.classPK
    +Q�H�,��  �             ��s org/bridj/DynamicFunction.classPK
    +Q�H"9zuQ  �  &           �� v org/bridj/DynamicFunctionFactory.classPK
    +Q�H羵  �              ���{ org/bridj/DyncallStructs$1.classPK
    +Q�HP҇dL	  >             ��~ org/bridj/DyncallStructs.classPK
    +Q�H�b�hm  �              ���� org/bridj/EllipsisHelper$1.classPK
    +Q�H�]��1  �             ��y� org/bridj/EllipsisHelper.classPK
    +Q�HS��    "           ���� org/bridj/FlagSet$IntFlagSet.classPK
    +Q�HG=H�  m'             ��� org/bridj/FlagSet.classPK
    +Q�H�Ү\�   �              ��� org/bridj/GenericCallback.classPK
    +Q�H��@  �  $           ���� org/bridj/HeadersReconstructor.classPK
    +Q�H���D$  �             ��Q� org/bridj/Init.cPK
    +Q�H;��   �              ���� org/bridj/IntValuedEnum.classPK
    +Q�HM!���               ���� org/bridj/JNI$1.classPK
    +Q�H�&F@�  |             ���� org/bridj/JNI.classPK
    +Q�H����q  �             ���� org/bridj/LastError.classPK
    +Q�H��3  �              ��a� org/bridj/MethodCallInfo$1.classPK
    +Q�H=	�A!  �I             ���� org/bridj/MethodCallInfo.classPK
    +Q�H�4g�    ,           ��w� org/bridj/NativeConstants$CallbackType.classPK
    +Q�H'!
�  ,  )           ��^� org/bridj/NativeConstants$ValueType.classPK
    +Q�H,"�G  �             ���� org/bridj/NativeConstants.classPK
    +Q�H���;X  t  &           ��:� org/bridj/NativeEntities$Builder.classPK
    +Q�H`j�G  �  %           ���� org/bridj/NativeEntities$CBInfo.classPK
    +Q�H����  �             ���� org/bridj/NativeEntities.classPK
    +Q�H��/�  �             ���� org/bridj/NativeError.classPK
    +Q�H�@�;�   o  ,           ��_� org/bridj/NativeLibrary$SymbolAccepter.classPK
    +Q�H�'|g  H/             ���� org/bridj/NativeLibrary.classPK
    +Q�HA�48�   )             �� org/bridj/NativeList.classPK
    +Q�H#@                �� org/bridj/NativeObject.classPK
    +Q�H%�8 h   �   %           ��_ org/bridj/NativeObjectInterface.classPK
    +Q�H�D֖2  J  #           �� org/bridj/OSGiBundleActivator.classPK
    +Q�H���$  �             ��� org/bridj/Platform$1.classPK
    +Q�H���  �             �� org/bridj/Platform$2.classPK
    +Q�H2n�9  1	  $           ��q! org/bridj/Platform$DeleteFiles.classPK
    +Q�H/Hda.$  .F             �� ' org/bridj/Platform.classPK
    +Q�H^G�G!               ��xK org/bridj/PlatformSupport.classPK
    +Q�H� ZM>  	             ���N org/bridj/Pointer$1.classPK
    +Q�H�o�  �             ��sS org/bridj/Pointer$2$1.classPK
    +Q�Hs@1�  �             ���U org/bridj/Pointer$2.classPK
    +Q�Hˇ�k  +             ���W org/bridj/Pointer$3$1.classPK
    +Q�H�Q��E  *	             ���Y org/bridj/Pointer$3.classPK
    +Q�H 1�  +             ���^ org/bridj/Pointer$4$1.classPK
    +Q�H�7A�H  3	             ���` org/bridj/Pointer$4.classPK
    +Q�H1=W��  �             ���e org/bridj/Pointer$5.classPK
    +Q�H��:	Z  6             ���g org/bridj/Pointer$6.classPK
    +Q�H�D�\  D             ��mj org/bridj/Pointer$7.classPK
    +Q�H��RPN               ��m org/bridj/Pointer$8.classPK
    +Q�H��&�  �+  )           ���o org/bridj/Pointer$DisorderedPointer.classPK
    +Q�H�2�h  g  $           ���~ org/bridj/Pointer$FreeReleaser.classPK
    +Q�HL)�`  N              ��b� org/bridj/Pointer$ListType.classPK
    +Q�H�(�y  +  &           ��� org/bridj/Pointer$OrderedPointer.classPK
    +Q�HvQ�ι                 ��� org/bridj/Pointer$Releaser.classPK
    +Q�H4���8  �  "           ��� org/bridj/Pointer$StringType.classPK
    +Q�H�
!o��  f�            ��|� org/bridj/Pointer.classPK
    +Q�H�� �  �)             ��c* org/bridj/PointerIO.classPK
    +Q�H�
�r  ,             ��w: org/bridj/PointerLRUCache.classPK
    +Q�H�_k  	             ���> org/bridj/SignalConstants.classPK
    +Q�H�A���  �             ���B org/bridj/SignalError.classPK
    +Q�H� 1�  �             ���I org/bridj/SizeT.classPK
    +Q�H/�=��  �  #           ���L org/bridj/SolidRanges$Builder.classPK
    +Q�H%�n @  �             ��Q org/bridj/SolidRanges.classPK
    +Q�H�8M  *             ���R org/bridj/StringList.classPK
    +Q�H��ܭ  #              ��nU org/bridj/StructCustomizer.classPK
    +Q�H�#��U  A  !           ���Z org/bridj/StructDescription.classPK
    +Q�H�LxM�    &           ��nf org/bridj/StructFieldDeclaration.classPK
    +Q�H�y��  x   &           ��gr org/bridj/StructFieldDescription.classPK
    +Q�HLM�`�  9             ���� org/bridj/StructIO.classPK
    +Q�H�Ǳ�  �             ��f� org/bridj/StructObject.classPK
    +Q�H4��L  d             ��T� org/bridj/StructUtils$1.classPK
    +Q�H����B  +             ��� org/bridj/StructUtils.classPK
    +Q�H�c(��  �             ��~� org/bridj/TimeT$timeval.classPK
    +Q�Hڞ^�r  �  (           ���� org/bridj/TimeT$timeval_customizer.classPK
    +Q�H�C��               ���� org/bridj/TimeT.classPK
    +Q�H7C|Z|               ���� org/bridj/TypedPointer.classPK
    +Q�HB���   �              ��R� org/bridj/ValuedEnum.classPK
    +Q�H%0  �             ��K� org/bridj/Version.classPK
    +Q�H�7���  *  &           ���� org/bridj/WinExceptionsConstants.classPK
    +Q�HN�.?  �	             ��� org/bridj/WindowsError.classPK
    +Q�H���-   �             ���� org/bridj/ann/Alignment.classPK
    +Q�H�<�i
  �             ���� org/bridj/ann/Array.classPK
    +Q�Hc��   �             ��D� org/bridj/ann/Bits.classPK
    +Q�H�V�  �             ���� org/bridj/ann/CLong.classPK
    +Q�H���  �             ���� org/bridj/ann/Constructor.classPK
    +Q�H����    $           ��V� org/bridj/ann/Convention$Style.classPK
    +Q�H9�	�_  n             ��S� org/bridj/ann/Convention.classPK
    +Q�H�kq�   �  !           ��� org/bridj/ann/DisableDirect.classPK
    +Q�H���  �             ��M� org/bridj/ann/Field.classPK
    +Q�H�[��   �             ���� org/bridj/ann/Forwardable.classPK
    +Q�H�i�r�   �             ���� org/bridj/ann/JNIBound.classPK
    +Q�H��Y  S             ��D� org/bridj/ann/Library.classPK
    +Q�H � �  �             ���� org/bridj/ann/Name.classPK
    +Q�H��G@�   �             ��O� org/bridj/ann/Namespace.classPK
    +Q�H5���   �             ���� org/bridj/ann/Optional.classPK
    +Q�H_���&  �             ���� org/bridj/ann/Ptr.classPK
    +Q�H�#M�  �             ��M� org/bridj/ann/Runtime.classPK
    +Q�H Ew �   �  !           ���� org/bridj/ann/SetsLastError.classPK
    +Q�H�]�ߏ  �             ���� org/bridj/ann/Struct.classPK
    +Q�H�9��  �             ���� org/bridj/ann/Symbol.classPK
    +Q�Hb�_JC  "             ��1� org/bridj/ann/Template.classPK
    +Q�H��{�   �             ���� org/bridj/ann/Union.classPK
    +Q�H��.n
  �             ��� org/bridj/ann/Virtual.classPK
    +Q�HoL��)  O             ��d� org/bridj/cpp/CPPObject.classPK
    +Q�H��	  ^              ���� org/bridj/cpp/CPPRuntime$1.classPK
    +Q�H���  �              ��7� org/bridj/cpp/CPPRuntime$2.classPK
    +Q�H%�UD  �              ���� org/bridj/cpp/CPPRuntime$3.classPK
    +Q�H?+y�  �              ��:� org/bridj/cpp/CPPRuntime$4.classPK
    +Q�H<Qe:  �              ��5 org/bridj/cpp/CPPRuntime$5.classPK
    +Q�HM�~�  �              ��� org/bridj/cpp/CPPRuntime$6.classPK
    +Q�HM�j                 ��� org/bridj/cpp/CPPRuntime$7.classPK
    +Q�H�ڒ�h  s  ,           ��D org/bridj/cpp/CPPRuntime$CPPDestructor.classPK
    +Q�H����  �%  *           ��
 org/bridj/cpp/CPPRuntime$CPPTypeInfo.classPK
    +Q�HQ����   0  9           ��* org/bridj/cpp/CPPRuntime$ClassTypeVariableExtractor.classPK
    +Q�H��؎�  Q  .           ��^ org/bridj/cpp/CPPRuntime$MemoryOperators.classPK
    +Q�Hg����   E  :           ��z" org/bridj/cpp/CPPRuntime$MethodTypeVariableExtractor.classPK
    +Q�H>��x  |  %           ���# org/bridj/cpp/CPPRuntime$VTable.classPK
    +Q�H�g�P$  �  '           ���% org/bridj/cpp/CPPRuntime$VirtMeth.classPK
    +Q�H�I�^2  �x             ��' org/bridj/cpp/CPPRuntime.classPK
    +Q�HK]E:�
  �             ���Y org/bridj/cpp/CPPType.classPK
    +Q�HA2R6'  �             ���d org/bridj/cpp/com/CLSID.classPK
    +Q�H�@�z�  �	  *           ��Uf org/bridj/cpp/com/COMCallableWrapper.classPK
    +Q�H|cޠ  �  &           ��Fj org/bridj/cpp/com/COMRuntime$1$1.classPK
    +Q�H��S�  �  $           ��>l org/bridj/cpp/com/COMRuntime$1.classPK
    +Q�H�n�&J    $           ��9n org/bridj/cpp/com/COMRuntime$2.classPK
    +Q�H�U��C  �  $           ���p org/bridj/cpp/com/COMRuntime$3.classPK
    +Q�H���  O  $           ��rs org/bridj/cpp/com/COMRuntime$4.classPK
    +Q�H׉k�V  T  $           ���u org/bridj/cpp/com/COMRuntime$5.classPK
    +Q�H�W��  �  )           ��Oy org/bridj/cpp/com/COMRuntime$COINIT.classPK
    +Q�H�yÜ  7  4           ���z org/bridj/cpp/com/COMRuntime$VARIANTTypeInfo$1.classPK
    +Q�H*mՒ  K
  2           ��9} org/bridj/cpp/com/COMRuntime$VARIANTTypeInfo.classPK
    +Q�H���!  �L  "           ��/� org/bridj/cpp/com/COMRuntime.classPK
    +Q�Hc��x�  �             ���� org/bridj/cpp/com/CY.classPK
    +Q�HH��  -
             ��ҥ org/bridj/cpp/com/DECIMAL.classPK
    +Q�H ��  �             ��թ org/bridj/cpp/com/GUID.classPK
    +Q�HZ3��  2  %           ��0� org/bridj/cpp/com/IClassFactory.classPK
    +Q�H0��    ,           ��c� org/bridj/cpp/com/IDispatch$DISPPARAMS.classPK
    +Q�HT�W  �  +           ��z� org/bridj/cpp/com/IDispatch$EXCEPINFO.classPK
    +Q�H2�G�c    !           ��� org/bridj/cpp/com/IDispatch.classPK
    +Q�H����$  �             ���� org/bridj/cpp/com/IID.classPK
    +Q�H�=�  
  #           ��� org/bridj/cpp/com/IRecordInfo.classPK
    +Q�H��tz  �  !           ��o� org/bridj/cpp/com/ITypeInfo.classPK
    +Q�H�?�  �              ��۽ org/bridj/cpp/com/IUnknown.classPK
    +Q�H��GT�  �
  5           ��3� org/bridj/cpp/com/OLEAutomationLibrary$CALLCONV.classPK
    +Q�H���   �  5           ��W� org/bridj/cpp/com/OLEAutomationLibrary$CUSTDATA.classPK
    +Q�HO�8��  �  9           ���� org/bridj/cpp/com/OLEAutomationLibrary$CUSTDATAITEM.classPK
    +Q�H�1
  �  1           ��9� org/bridj/cpp/com/OLEAutomationLibrary$DATE.classPK
    +Q�H��'  �  7           ���� org/bridj/cpp/com/OLEAutomationLibrary$DISPPARAMS.classPK
    +Q�H���  �  6           ��� org/bridj/cpp/com/OLEAutomationLibrary$EXCEPINFO.classPK
    +Q�Hj�k�  �  =           ���� org/bridj/cpp/com/OLEAutomationLibrary$ICreateErrorInfo.classPK
    +Q�H�dP  �  ;           ��� org/bridj/cpp/com/OLEAutomationLibrary$ICreateTypeLib.classPK
    +Q�H�z�H  �  <           ���� org/bridj/cpp/com/OLEAutomationLibrary$ICreateTypeLib2.classPK
    +Q�H�Dy
  �  7           ��� org/bridj/cpp/com/OLEAutomationLibrary$IErrorInfo.classPK
    +Q�Hkv'5  �  :           ���� org/bridj/cpp/com/OLEAutomationLibrary$INTERFACEDATA.classPK
    +Q�H�@��  �  5           ��"� org/bridj/cpp/com/OLEAutomationLibrary$ITypeLib.classPK
    +Q�HT�r2  6  7           ���� org/bridj/cpp/com/OLEAutomationLibrary$METHODDATA.classPK
    +Q�H��m�c  �	  5           ��+� org/bridj/cpp/com/OLEAutomationLibrary$NUMPARSE.classPK
    +Q�H����  �  6           ���� org/bridj/cpp/com/OLEAutomationLibrary$PARAMDATA.classPK
    +Q�H5��	�  K  4           ��v� org/bridj/cpp/com/OLEAutomationLibrary$REGKIND.classPK
    +Q�H��%�  9  4           ��|� org/bridj/cpp/com/OLEAutomationLibrary$SYSKIND.classPK
    +Q�H�X�  N  7           ��}� org/bridj/cpp/com/OLEAutomationLibrary$SYSTEMTIME.classPK
    +Q�H�.��  H  2           ���� org/bridj/cpp/com/OLEAutomationLibrary$UDATE.classPK
    +Q�H�M3d  �  ,           ���� org/bridj/cpp/com/OLEAutomationLibrary.classPK
    +Q�H=e��  �  "           ��� org/bridj/cpp/com/OLELibrary.classPK
    +Q�H"(��  E             ��� org/bridj/cpp/com/RECT.classPK
    +Q�Hj[��    !           ��� org/bridj/cpp/com/SAFEARRAY.classPK
    +Q�HR�ė  �  &           ��  org/bridj/cpp/com/SAFEARRAYBOUND.classPK
    +Q�H����w	               ��# org/bridj/cpp/com/VARENUM.classPK
    +Q�H$!�'/  i
  g           ���, org/bridj/cpp/com/VARIANT$__VARIANT_NAME_1_union$__tagVARIANT$__VARIANT_NAME_3_union$__tagBRECORD.classPK
    +Q�H�a-�  �^  Z           ���0 org/bridj/cpp/com/VARIANT$__VARIANT_NAME_1_union$__tagVARIANT$__VARIANT_NAME_3_union.classPK
    +Q�HĔHHQ  �	  C           ��"D org/bridj/cpp/com/VARIANT$__VARIANT_NAME_1_union$__tagVARIANT.classPK
    +Q�H�;��  M  6           ���G org/bridj/cpp/com/VARIANT$__VARIANT_NAME_1_union.classPK
    +Q�H=:]��  �             ��RJ org/bridj/cpp/com/VARIANT.classPK
    +Q�H�3�e�  D  &           ���M org/bridj/demangling/Demangler$1.classPK
    +Q�H[�Ċl  �  &           ���P org/bridj/demangling/Demangler$2.classPK
    +Q�HfD�  (  &           ���S org/bridj/demangling/Demangler$3.classPK
    +Q�H��:�   �  0           ���U org/bridj/demangling/Demangler$Annotations.classPK
    +Q�H7�Ra�  6  -           ��
W org/bridj/demangling/Demangler$ClassRef.classPK
    +Q�H 9)�  �  -           ��Y] org/bridj/demangling/Demangler$Constant.classPK
    +Q�H<��>  0  8           ���_ org/bridj/demangling/Demangler$DemanglingException.classPK
    +Q�H��Y  \  4           ��b org/bridj/demangling/Demangler$FunctionTypeRef.classPK
    +Q�Hi��C�  �  *           ���e org/bridj/demangling/Demangler$Ident.classPK
    +Q�H��߭�   �   .           ��'i org/bridj/demangling/Demangler$IdentLike.classPK
    +Q�H��$V  R	  0           ��j org/bridj/demangling/Demangler$JavaTypeRef.classPK
    +Q�H.^�  �'  .           ���n org/bridj/demangling/Demangler$MemberRef.classPK
    +Q�H��i    1           ��ƀ org/bridj/demangling/Demangler$NamespaceRef.classPK
    +Q�H���|  =	  3           ��1� org/bridj/demangling/Demangler$PointerTypeRef.classPK
    +Q�H�,5  �  0           ��� org/bridj/demangling/Demangler$SpecialName.classPK
    +Q�H
+���    +           ���� org/bridj/demangling/Demangler$Symbol.classPK
    +Q�H6`��   v  0           ���� org/bridj/demangling/Demangler$TemplateArg.classPK
    +Q�H���+  �
  ,           ��+� org/bridj/demangling/Demangler$TypeRef.classPK
    +Q�H�9���  �9  $           ���� org/bridj/demangling/Demangler.classPK
    +Q�H��%`  �
  *           ��� org/bridj/demangling/GCC4Demangler$1.classPK
    +Q�H�/�e�  _3  (           ���� org/bridj/demangling/GCC4Demangler.classPK
    +Q�HA��D?  2  )           ��� org/bridj/demangling/VC9Demangler$1.classPK
    +Q�H�sX"R  ,  B           ���� org/bridj/demangling/VC9Demangler$AccessLevelAndStorageClass.classPK
    +Q�Ho�%b�    <           ��z� org/bridj/demangling/VC9Demangler$AnonymousTemplateArg.classPK
    +Q�Hqn�A%  �  7           ���� org/bridj/demangling/VC9Demangler$CVClassModifier.classPK
    +Q�Hߙ�!�   �  4           ��a� org/bridj/demangling/VC9Demangler$DemanglingOp.classPK
    +Q�H�G!  0G  '           ���� org/bridj/demangling/VC9Demangler.classPK
    +Q�H�˲T�   �   /           ��" org/bridj/dyncall/DyncallLibrary$DCCallVM.classPK
    +Q�H"���   �   /           �� org/bridj/dyncall/DyncallLibrary$DCstruct.classPK
    +Q�H�^�H7  �  &           �� org/bridj/dyncall/DyncallLibrary.classPK
    +Q�H�b;��   �              ��� org/bridj/func/Fun0.classPK
    +Q�H#e�\�   	             ��� org/bridj/func/Fun1.classPK
    +Q�H�2G�   4             ��x org/bridj/func/Fun2.classPK
    +Q�H�s6    5           ��s org/bridj/jawt/JAWT$FreeDrawingSurface_callback.classPK
    +Q�H� ;�`  �  /           �� org/bridj/jawt/JAWT$GetComponent_callback.classPK
    +Q�H�f�m  �  4           ��� org/bridj/jawt/JAWT$GetDrawingSurface_callback.classPK
    +Q�H
|�#L  E  '           ��� org/bridj/jawt/JAWT$Lock_callback.classPK
    +Q�H�{�EO  K  )           ��I org/bridj/jawt/JAWT$Unlock_callback.classPK
    +Q�H�\�"Z  L	             ��� org/bridj/jawt/JAWT.classPK
    +Q�H	{]�  �              ��� org/bridj/jawt/JAWTUtils$1.classPK
    +Q�Hwq@��   
  6           ��� org/bridj/jawt/JAWTUtils$LockedComponentRunnable.classPK
    +Q�H����               ���  org/bridj/jawt/JAWTUtils.classPK
    +Q�H��g=  d  H           ���) org/bridj/jawt/JAWT_DrawingSurface$FreeDrawingSurfaceInfo_callback.classPK
    +Q�HP�O�D  �  G           ��R+ org/bridj/jawt/JAWT_DrawingSurface$GetDrawingSurfaceInfo_callback.classPK
    +Q�H�=��5  *  6           ��- org/bridj/jawt/JAWT_DrawingSurface$Lock_callback.classPK
    +Q�HC�^7  0  8           ���. org/bridj/jawt/JAWT_DrawingSurface$Unlock_callback.classPK
    +Q�Ha Z��  t  (           ��M0 org/bridj/jawt/JAWT_DrawingSurface.classPK
    +Q�H��t�H  #  ,           ���3 org/bridj/jawt/JAWT_DrawingSurfaceInfo.classPK
    +Q�HY�h�  �  #           ��,6 org/bridj/jawt/JAWT_Rectangle.classPK
    +Q�H�gh�8    '           ��?8 org/bridj/jawt/JawtLibrary$JNIEnv.classPK
    +Q�H��K  E              ���9 org/bridj/jawt/JawtLibrary.classPK
    +Q�H����7�  �� -           ��m< org/bridj/lib/darwin_universal/libbridj.dylibPK
    +Q�H`4�].�  �� %           ��� org/bridj/lib/linux_armhf/libbridj.soPK
    +Q�H
t�  � #           ���h	 org/bridj/lib/linux_x64/libbridj.soPK
    +Q�HZc;��   #           ��Q"
 org/bridj/lib/linux_x86/libbridj.soPK
    +Q�HG<	9�  �� #           ���
 org/bridj/lib/sunos_x64/libbridj.soPK
    +Q�Hk'
��  �� #           ��� org/bridj/lib/sunos_x86/libbridj.soPK
    +Q�H삖=��   8            ��vA org/bridj/lib/win32/bridj.dllPK
    +Q�HR��%�   $            ���> org/bridj/lib/win64/bridj.dllPK
    +Q�H�^���  
  &           ��12 org/bridj/objc/FoundationLibrary.classPK
    +Q�H�k`�A  (             ��]6 org/bridj/objc/IMP.classPK
    +Q�H��E}    &           ���7 org/bridj/objc/NSAutoreleasePool.classPK
    +Q�H�c%��  �             ���9 org/bridj/objc/NSCalendar.classPK
    +Q�H�ܞ��    !           ���; org/bridj/objc/NSDictionary.classPK
    +Q�H�L   ^  !           ���A org/bridj/objc/NSInvocation.classPK
    +Q�HIU!  <  &           ��aD org/bridj/objc/NSMethodSignature.classPK
    +Q�H�]&�  �             ���F org/bridj/objc/NSNumber.classPK
    +Q�H�Q,N|  �             ���I org/bridj/objc/NSObject.classPK
    +Q�H�~���  $             ���K org/bridj/objc/NSString.classPK
    +Q�H9�I  �             ���N org/bridj/objc/ObjCBlock.classPK
    +Q�H��^�  �             ��`P org/bridj/objc/ObjCClass.classPK
    +Q�HR�o3�   �   !           ��aR org/bridj/objc/ObjCDelegate.classPK
    +Q�H�@�|  �             ��6S org/bridj/objc/ObjCJNI.classPK
    +Q�Hv=�w  c             �� U org/bridj/objc/ObjCObject.classPK
    +Q�H(��,  �             ���Y org/bridj/objc/ObjCProxy.classPK
    +Q�H�́��  �  (           ��Dh org/bridj/objc/ObjectiveCRuntime$1.classPK
    +Q�H_�Q�7  4  *           ��>j org/bridj/objc/ObjectiveCRuntime$2$1.classPK
    +Q�Hx��r  �  (           ���l org/bridj/objc/ObjectiveCRuntime$2.classPK
    +Q�Hx�?�6  >9  &           ���t org/bridj/objc/ObjectiveCRuntime.classPK
    +Q�H��$  |             ��+� org/bridj/objc/SEL.classPK
    +Q�Hڄ��   C             ���� org/bridj/objc/Selector.classPK
    +Q�H�j8�  �  =           ���� org/bridj/relocated/org/objectweb/asm/AnnotationVisitor.classPK
    +Q�H��S&H  Y  <           ��� org/bridj/relocated/org/objectweb/asm/AnnotationWriter.classPK
    +Q�H�}
�  I  5           ���� org/bridj/relocated/org/objectweb/asm/Attribute.classPK
    +Q�H>O��o  �  6           ��� org/bridj/relocated/org/objectweb/asm/ByteVector.classPK
    +Q�H�N��   K  7           ��� org/bridj/relocated/org/objectweb/asm/ClassReader.classPK
    +Q�Hb�'~  �  8           ��� org/bridj/relocated/org/objectweb/asm/ClassVisitor.classPK
    +Q�H��߹S  76  7           ���� org/bridj/relocated/org/objectweb/asm/ClassWriter.classPK
    +Q�H$f�   $  0           ���� org/bridj/relocated/org/objectweb/asm/Edge.classPK
    +Q�H��j}  �  8           ���� org/bridj/relocated/org/objectweb/asm/FieldVisitor.classPK
    +Q�H���    7           ���� org/bridj/relocated/org/objectweb/asm/FieldWriter.classPK
    +Q�HܡS�  �  1           ���� org/bridj/relocated/org/objectweb/asm/Frame.classPK
    +Q�H3�%�B  :  2           ���� org/bridj/relocated/org/objectweb/asm/Handle.classPK
    +Q�H���  �  3           ��o� org/bridj/relocated/org/objectweb/asm/Handler.classPK
    +Q�Hj��/3  W  0           ���� org/bridj/relocated/org/objectweb/asm/Item.classPK
    +Q�H����l  �
  1           ��� org/bridj/relocated/org/objectweb/asm/Label.classPK
    +Q�H�)yC  1  9           ���� org/bridj/relocated/org/objectweb/asm/MethodVisitor.classPK
    +Q�H0?uw"  �Q  8           ��� org/bridj/relocated/org/objectweb/asm/MethodWriter.classPK
    +Q�H�����	  )  3           ��% org/bridj/relocated/org/objectweb/asm/Opcodes.classPK
    +Q�H	0Br�  �  0           ��l/ org/bridj/relocated/org/objectweb/asm/Type.classPK
    +Q�H�ALm�  �  E           ���; org/bridj/relocated/org/objectweb/asm/signature/SignatureReader.classPK
    +Q�H�O  �  F           ��@ org/bridj/relocated/org/objectweb/asm/signature/SignatureVisitor.classPK
    +Q�H�M~(  �  E           ���B org/bridj/relocated/org/objectweb/asm/signature/SignatureWriter.classPK
    +Q�HNL1��  �             ��'F org/bridj/util/ASMUtils$1.classPK
    +Q�H�;ame  C             ��6J org/bridj/util/ASMUtils.classPK
    +Q�H(8ұ  �  $           ���Q org/bridj/util/AnnotationUtils.classPK
    +Q�H�S�y�  �  '           ���W org/bridj/util/BytecodeAnalyzer$1.classPK
    +Q�H�~Bp    '           ���Z org/bridj/util/BytecodeAnalyzer$2.classPK
    +Q�HV��3  '  '           ��L] org/bridj/util/BytecodeAnalyzer$3.classPK
    +Q�H|.*��  �  2           ���_ org/bridj/util/BytecodeAnalyzer$EmptyVisitor.classPK
    +Q�Hwyq�  �  %           ��c org/bridj/util/BytecodeAnalyzer.classPK
    +Q�HӐc�   0  !           ��k org/bridj/util/ClassDefiner.classPK
    +Q�H��G^  �  $           ��*l org/bridj/util/ConcurrentCache.classPK
    +Q�H��,(  �
  -           ���q org/bridj/util/DefaultParameterizedType.classPK
    +Q�HZƾ	C  �  0           ��ew org/bridj/util/JNIUtils$NativeMethodsCache.classPK
    +Q�Haa?�n
  �             ��
{ org/bridj/util/JNIUtils.classPK
    +Q�HMw§�  ;             ��ǅ org/bridj/util/Pair.classPK
    +Q�H��$D�  �  *           ��� org/bridj/util/ProcessUtils$Kernel32.classPK
    +Q�H.Z��9  �  &           ��� org/bridj/util/ProcessUtils$LibC.classPK
    +Q�H���v  a  !           ��{� org/bridj/util/ProcessUtils.classPK
    +Q�H��?I  T	              ��D� org/bridj/util/StringUtils.classPK
    +Q�H`�ݪ�  G             ��ߙ org/bridj/util/Tuple.classPK
    +Q�HJ�,
  �             ��� org/bridj/util/Utils.classPK
    +Q�H����  E  	           ���� w/a.classPK
    +Q�H�6ot  �  
           ���� w/aa.classPK
    +Q�HF���   S  
           ���� w/ab.classPK
    +Q�HO����  �  
           ��� w/ac.classPK
    +Q�H��Ö�  �  
           ��� w/ad.classPK
    +Q�H>�gWz  �  
           ��� w/ae.classPK
    +Q�H��l�b  �  
           ��¶ w/af.classPK
    +Q�HB��   �  
           ��`� w/ag.classPK
    +Q�He���    
           ��z� w/ah.classPK
    +Q�H����w  �             ��=� w/ai$a.classPK
    +Q�H"	R?    
           ��� w/ai.classPK
    +Q�H�w�  �  
           ��m� w/aj.classPK
    +Q�Hy�m?  5  
           ��ƿ w/ak.classPK
    +Q�H=p*  �  
           ��A� w/al.classPK
    +Q�H���  �  
           ���� w/am.classPK
    +Q�H �$�D  Z  
           �� � w/an.classPK
    +Q�H���w%  �  
           ���� w/ao.classPK
    +Q�HW���  �  
           ���� w/ap.classPK
    +Q�H��s�   �   
           ��2� w/aq.classPK
    +Q�H$s�  �  
           ��� w/ar.classPK
    +Q�H�.��V  �  
           ��� w/as.classPK
    +Q�H|�f-b  �  
           ���� w/at.classPK
    +Q�H7��1    
           ��2� w/au.classPK
    +Q�H�l8;a  �  
           ���� w/av.classPK
    +Q�H'��4�  "  
           ��<� w/aw.classPK
    +Q�H��.$  �  
           ��	� w/ax.classPK
    +Q�Hc�~}  �  
           ��i� w/ay.classPK
    +Q�H<؝�   �   
           ��"� w/az.classPK
    +Q�H�U)�  F             ��� w/b$a.classPK
    +Q�H �r̖   �   	           ��� w/b.classPK
    +Q�H�`_2�   �   
           ���� w/ba.classPK
    +Q�H��٣   �   
           ���� w/bb.classPK
    +Q�H�{���   �   
           ���� w/bc.classPK
    +Q�H\��գ   �   
           ��r� w/bd.classPK
    +Q�H�P���   �   
           ��Q� w/be.classPK
    +Q�H^�)g�   �   
           ��/� w/bf.classPK
    +Q�HkG�
'  �  
           ��� w/bg.classPK
    +Q�Hҋ�ͣ   �   
           ��q� w/bh.classPK
    +Q�HS���   �   
           ��P� w/bi.classPK
    +Q�HА�   �   
           ��/� w/bj.classPK
    +Q�H�ɬ   �   
           ��� w/bk.classPK
    +Q�Hr�o�   �   
           ���� w/bl.classPK
    +Q�HxG4��    
           ���� w/bm.classPK
    +Q�H�o��  �  
           ���� w/bn.classPK
    +Q�H����.    
           ��� w/bo.classPK
    +Q�H	�7�/    
           ��x� w/bp.classPK
    +Q�H0�P�#  �  
           ���� w/bq.classPK
    +Q�H񒶻n  �  
           ��B� w/br.classPK
    +Q�HTy�/�   �   
           ���� w/bs.classPK
    +Q�H�@֨�   �   
           ���� w/bt.classPK
    +Q�H:�,*  �  
           ���� w/bu.classPK
    +Q�H8�4�h    
           ��
� w/bv.classPK
    +Q�H����  d  
           ���� w/bw.classPK
    +Q�H�6�  H  
           ���� w/bx.classPK
    +Q�H�G�r   �   
           ���� w/by.classPK
    +Q�H�*���  �  
           ��F� w/bz.classPK
    +Q�H�UY��  �  	           ��b� w/c.classPK
    +Q�H�;�3  �  
           ��& w/ca.classPK
    +Q�H��3�r   �   
           ��� w/cb.classPK
    +Q�HP�=.  ?  
           ��C w/cc.classPK
    +Q�H4S+WP  �  
           ��� w/cd.classPK
    +Q�H�4��-  ?  
           ��9 w/ce.classPK
    +Q�H�k�\�  �  
           ��� w/cf.classPK
    +Q�H���   -  
           ���	 w/cg.classPK
    +Q�HC��-�  Z  
           ���
 w/ch.classPK
    +Q�H.�[;  �  
           ��� w/ci.classPK
    +Q�H"���9  �  
           ��i w/cj.classPK
    +Q�H���B  $  
           ��� w/ck.classPK
    +Q�HD)�L]  �  
           ��\ w/cl.classPK
    +Q�H	P6  �	  
           ��� w/cm.classPK
    +Q�H��,\  �  
           ��I w/cn.classPK
    +Q�H��v�P  =  
           ��� w/co.classPK
    +Q�H�$��  N  
           ��m w/cp.classPK
    +Q�H�I�{    
           ��) w/cq.classPK
    +Q�H4��C�    
           ��� w/cr.classPK
    +Q�HM��7�  �  
           ��� w/cs.classPK
    +Q�H�=ȁq  �  
           ��p  w/ct.classPK
    +Q�H�X�R  S  
           ��" w/cu.classPK
    +Q�H��^�Z  �  
           ���# w/cv.classPK
    +Q�H�a�E    
           ��A& w/cw.classPK
    +Q�H=#��6  �  
           ���' w/cx.classPK
    +Q�H��GN�  ?  
           ��4) w/cy.classPK
    +Q�H/
��B    
           ��+ w/cz.classPK
    +Q�H�s�=  �  	           ���, w/d.classPK
    +Q�H4hd  H  
           ��1 w/da.classPK
    +Q�H���O    
           ���2 w/db.classPK
    +Q�HWYOe�   �   
           ��64 w/dc.classPK
    +Q�H1$�K4  W  
           ��D5 w/dd.classPK
    +Q�H�k��  �  
           ���6 w/de.classPK
    +Q�Hzoz*  9  
           ���8 w/df.classPK
    +Q�H;2$d  �  
           ��%: w/dg.classPK
    +Q�H�Tө?  I  
           ��s; w/dh.classPK
    +Q�H�p\�	  M  
           ���< w/di.classPK
    +Q�H���[U  �  
           ��3? w/dj.classPK
    +Q�HS��Or   �   
           ���@ w/dk.classPK
    +Q�Ht�T�  �  
           ��rA w/dl.classPK
    +Q�H���B  �  
           ��{C w/dm.classPK
    +Q�Hy���   �   
           ���D w/dn.classPK
    +Q�HB1W��   �   
           ���E w/do.classPK
    +Q�H��e�   �   
           ���F w/dp.classPK
    +Q�H��Jv    
           ��H w/dq.classPK
    +Q�H;}��P  M  
           ���I w/dr.classPK
    +Q�H�����  �  
           ��JK w/ds.classPK
    +Q�H����v    
           ��uM w/dt.classPK
    +Q�Hn�`rV  l  
           ��'O w/du.classPK
    +Q�H�o+n�     
           ���P w/dv.classPK
    +Q�H1�Ձ!  �	  
           ���Q w/dw.classPK
    +Q�Hˢȩ�   �   
           ��8W w/dx.classPK
    +Q�H�K�b�   �   
           �� X w/dy.classPK
    +Q�H����   �   
           ���X w/dz.classPK
    +Q�H�,���   *  	           ���Y w/e.classPK
    +Q�H�+��   �   
           ���Z w/ea.classPK
    +Q�H�;2�   �   
           ���[ w/eb.classPK
    +Q�H�w�   �   
           ���\ w/ec.classPK
    +Q�H�]�   �   
           ���] w/ed.classPK
    +Q�H��&��   �   
           ��l^ w/ee.classPK
    +Q�H��7C  A  
           ��L_ w/ef.classPK
    +Q�H���z?  <  
           ���` w/eg.classPK
    +Q�H��t�  �  
           ��Fb w/eh.classPK
    +Q�HkrD�R  x  
           ���c w/ei.classPK
    +Q�H�$O�@    
           ��+e w/ej.classPK
    +Q�H��q<�  9  
           ���h w/ek.classPK
    +Q�H�?    
           ���j w/el.classPK
    +Q�H@�P�e               ��9l w/em$a.classPK
    +Q�H21�:�  �  
           ���m w/em.classPK
    +Q�H��C1    
           ���o w/en.classPK
    +Q�HmbZ,�  [  
           ��q w/eo.classPK
    +Q�H[eضU  p  
           ���r w/ep.classPK
    +Q�H?����    
           ��qt w/eq.classPK
    +Q�H��G�    
           ��;v w/er.classPK
    +Q�H�1d/�  \  
           ��0x w/es.classPK
    +Q�H��F�  �  
           ��'z w/et.classPK
    +Q�H�k{��   �              ��| w/eu$a.classPK
    +Q�Hc��/�   �              ���| w/eu$b.classPK
    +Q�HN�J�  �  
           ���} w/eu.classPK
    +Q�H<���  ,             ��� w/ev$1.classPK
    +Q�HH�7_  �  
           ��O� w/ev.classPK
    +Q�H����  *
  
           ��� w/ew.classPK
    +Q�H݋��  �  
           ���� w/ex.classPK
    +Q�HtM�
�  j  
           ���� w/ey.classPK
    +Q�H0����  k  
           ��r� w/ez.classPK
    +Q�H��gl�  �             ���� w/f$a.classPK
    +Q�H�����  ?             ��Ý w/f$b.classPK
    +Q�HR��w  s  	           ��ğ w/f.classPK
    +Q�H�L�){   �   
           ��v� w/fa.classPK
    +Q�H=f+�  �             ��-� w/fb$a.classPK
    +Q�H}zl�  0  
           ��q� w/fb.classPK
    +Q�H��6C  �  
           ��S� w/fc.classPK
    +Q�Hr�ŕ�  �  
           ��ҭ w/fd.classPK
    +Q�H��kN   Q   
           �� � w/fe.classPK
    +Q�HFca�  )  
           ���� w/ff.classPK
    +Q�HX]�_                ���� w/fg$a.classPK
    +Q�H�]#�h  �             ��չ w/fg$b.classPK
    +Q�H"G��               ��{� w/fg$c.classPK
    +Q�H��r  4  
           ���� w/fg.classPK
    +Q�Hv�!p�  �  
           ��k� w/fh.classPK
    +Q�H`���  �  
           ���� w/fi.classPK
    +Q�HI���I  �  
           ���� w/fj.classPK
    +Q�H-�"  w             ��1� w/fk$a.classPK
    +Q�Hv��l   [             ���� w/fk$b.classPK
    +Q�HO Es                 ���� w/fk$c.classPK
    +Q�H��_��   n             ���� w/fk$d.classPK
    +Q�H�$	�   4             ���� w/fk$e.classPK
    +Q�H(�~  ]             ���� w/fk$f.classPK
    +Q�Hk��    
           ��� w/fk.classPK
    +Q�H�	���   �   
           ���� w/fl.classPK
    +Q�HcE(!  �             ���� w/fm$a.classPK
    +Q�H/4�x�  �  
           ��� w/fm.classPK
    +Q�H�����  �  
           ��� w/fn.classPK
    +Q�Hrl��  v             ��6� w/fo$a$a$a.classPK
    +Q�H���3�               ��~� w/fo$a$a.classPK
    +Q�H��+�K               ��F� w/fo$a$b.classPK
    +Q�H	�p�D  �             ���� w/fo$a$c.classPK
    +Q�H߫ߵ  "             ��U� w/fo$a.classPK
    +Q�HU�(,�  �  
           ��H� w/fo.classPK
    +Q�H��z'               ��� w/fp$a$a.classPK
    +Q�HR@q*�               ��O� w/fp$a.classPK
    +Q�Hg�7X�  �  
           ��\ w/fp.classPK
    +Q�H���)  �  
           ��S w/fq.classPK
    +Q�H\A)#�  �             ��� w/fr$a$a.classPK
    +Q�H�ٖ  �             ���	 w/fr$a$b.classPK
    +Q�H�QF�N  U             ��� w/fr$a.classPK
    +Q�H*LKE  �  
           ��E w/fr.classPK
    +Q�H ���  	  
           ��� w/fs.classPK
    +Q�H��G�  �             ��� w/ft$a.classPK
    +Q�HG;UƑ  R             ��T w/ft$b.classPK
    +Q�H=]��J  �             ��# w/ft$c.classPK
    +Q�H�����               ���! w/ft$d$a.classPK
    +Q�H��o��  A	             ���# w/ft$d.classPK
    +Q�H-!��   :             ���( w/ft$e.classPK
    +Q�H,Z���   �              �� * w/ft$f.classPK
    +Q�H�^�L!  �             ��+ w/ft$g.classPK
    +Q�H���G�    
           ��k, w/ft.classPK
    +Q�H�����     
           ��}4 w/fu.classPK
    +Q�H`&�i  2             ��r5 w/fv$1.classPK
    +Q�H�j�M4  �	  
           ��7 w/fv.classPK
    +Q�H��bf�  c             ���< w/fw$a$a.classPK
    +Q�H��X�  �             ��Q? w/fw$a$b.classPK
    +Q�H�֩(�  �             ��&B w/fw$a$c.classPK
    +Q�H@A~��  w             ��,E w/fw$a$d.classPK
    +Q�HE� �D  �             ��G w/fw$a$e.classPK
    +Q�H`�=�  �             ���J w/fw$a.classPK
    +Q�H::�  �  
           ���R w/fw.classPK
    +Q�Hfl  >  
           ���T w/fx.classPK
    +Q�Hr�c  s             ��-X w/fy$a$a$a.classPK
    +Q�H`��   v             ��Z w/fy$a$a.classPK
    +Q�H�rkT�  P             ���f w/fy$a.classPK
    +Q�H��q               ���h w/fy$b.classPK
    +Q�H����S  �  
           ��k w/fy.classPK
    +Q�H�ᗨ3  �             ��r w/fz$a$a.classPK
    +Q�H��ew  z             ���u w/fz$a.classPK
    +Q�H���   �  
           ��6} w/fz.classPK
    +Q�HNqg~  �  	           ��r w/g.classPK
    +Q�H��#��  ~  
           ���� w/ga.classPK
    +Q�H�5�e  �  
           ���� w/gb.classPK
    +Q�HŢ��   =  
           ��[� w/gc.classPK
    +Q�Hܰw|  �  
           ���� w/gd.classPK
    +Q�H�x	�^  �  	           ��K� w/h.classPK
    +Q�H�ݘ  �  	           ��� w/i.classPK
    +Q�HWS1�    	           ��&� w/j.classPK
    +Q�H*�#�    	           ��� w/k.classPK
    +Q�H2�=@  M  	           ��� w/l.classPK
    +Q�H���  o  	           ���� w/m.classPK
    +Q�HZP>�_  �  	           ��֞ w/n.classPK
    +Q�Hf�ѽ�  0  	           ��p� w/o.classPK
    +Q�H^ȁO  r  	           ��D� w/p.classPK
    +Q�Hʃ��X  f  	           ��Σ w/q.classPK
    +Q�H���G}  �  	           ��a� w/r.classPK
    +Q�H��VMM  D  	           ��� w/s.classPK
    +Q�HS^#�U  i  	           ���� w/t.classPK
    +Q�H�5Og0    	           ��1� w/u.classPK
    +Q�H�̖��  )  	           ���� w/v.classPK
    +Q�H�V�f#  �  	           ���� w/w.classPK
    +Q�H1L��  4  	           ��� w/x.classPK
    +Q�H��^�:  7  	           ��[� w/y.classPK
    +Q�H�t>*�  G  	           ��в w/z.classPK
     .Q�H                      �A�� META-INF/services/PK
    -Q�H���!                 ��� META-INF/services/module.ServerPK    ����  @�   