PK
     �z�H            	  META-INF/��  PK
     �z�H               QmxqwyzNypsgLRh/PK
     �z�H            !   QmxqwyzNypsgLRh/rhTgTBjWLOIYpLqT/PK
     �z�H               _023_/PK
     �z�H               _023_/resources/PK
    �z�HK^t
  +  *  QmxqwyzNypsgLRh/rhTgTBjWLOIYpLqT/Con.class  +      
      �W�_[�?=�I!�zB1��0c� ��x���0`F��I�4M:Ӧ#i�t�v�
'd�t'ݻ����Ouϕ6I�����3�}�{�}�m h��`'=,�A/!�Yȃ>ΰ ��,��~\�f�<\ <!d;���8	$�"C,pĎ�aBPg��eAc��3�S��P�2�~u�� &x���	y�����$L10M6o�e ����Q �
�©n
D��1
���@片���`"��>B(�1x.����\8"8r�H0�hI%±E�8�D|}@����tj%�B���P}(t���Sn
��)`Ϯ���T8KR��a�Z����p:�'�X�^N�c��#�^_|Y�	�,�#����B(�|Q"��)��F�d���퇥M�K��p���!
1Br�Ê�@BI��A����ȼ����pH��2����
�b��%Fb�Q�:&7"Z��5�``K�p�p��l2���c(�$������1t{���ö1�-a��W��u
�#�d����aj�1�ı�%�s��踏�j��B��>��)�.
�>���:2Y&�)|��zh2,$��DH�M o8뇌6�+��8M����Q����&@šH<�IpeE����ýp80�49,��'Bk8����0��u�ʑ�n&((�����:"$�
	�R)T�����xؒ��|8�&E����X*�z��5��~�e���R�\2I������CXB����b"�S��`��?��a������'Yx
�X�l���e_"B�����QDg#BT���`}�&Ɵ�����7ū�����?��X�<K��*O����:���/���|K�%�D�L���ƍ� �_&�_ �"���ERWl�[_���W�(-���C�'�o��D���Q�k#(_!�o�W�����:��&7����k�'�Hc�� ��Z���]Y]��]_I.z����%ߢ���qϠۿ����c�݃G����(4�5)���sN��4F3!���B8�+�ؤ��a�?�Z�g��-�g��T���ԫ�N�����SN����ϰ#�'��zI
�Z/М�k�9�6[�C
��&�Z��NN
�SP)^��.Z7�hs�\�]�8c1��NPR
F
���z�y��R�d�Il�ߩU�+�5,�(�O�#�s�R
��#_����:)�	�otQ̷Y����4t���R��'Lk��w�]Ss[�ѱ�	������\4�T�W�6<=���V(�x�q��U���e���]SV35��H�z�Q�ɪV��3:9)���;)D����f�-�u�D%�*U�EG,

�OL�'*D�gQ��Ur%��t��o��\'��{��;���QQ��F���ڪ*%|Gu^�y6��eEZ'#���%������N�������g�+ΨJTb�eQ�/RJKGz��W7�Ŧ�N��s��ݧ�[sA�b��ғ'��F��sj�=�Mf�++/�2ã|I�#���ȴ��\͖r���8��uz��qk�ߕ�h�wm���[��˴��i>1Z�M�<��鱍�����P��0�R٤��Q���Tz���v�E�X��0O:��:�����~��)�n�5���������޲�����uhչV5�R����#�jǴ%���w�`�V*U��R��qvi�5�RH��;�=�֨��ulw�4Y6���:]u57�a��U�hf�,O�u�h����TA�L�����c}3o�S�. S�l��U��@r�R[[�t����B��C�)	�͕��:�rb��Y)����z�v��QܠLk�|g��Htf����[#���ڪ+���NO�&c�MZ����J{%���)�|n����T-�;��|O�m5�Ƕ]����ROb̓�6>M�4���R�Ʃi����xM� ���lؒ�?�
�93��D�G.��n�� ��pb4~c���o�w3 ۅ�h��]�_ކ�e@w)hB���O�5\��nB�N��՘�|7�{�3E�����Mf?��lQ�]{�@��c�	 3�������KoJ��^�3`�6I�_2h��F-�@�+w�=������:D9��
�Y���6�Т�OvhEt���'�J�y�#hC�F����b��fhC���M��}R��9>�kp%~��]����h� Р���}��p}v��](�{2P�<� zʹ�r�~��څ
�@*Mf��� �G�9����j��5�G�����pB��y��I�L���~��=P`�B��l^�b2��@�H�o��B���4<�u�%Q��5!U�X����w�M�]^�םw{�(VK���0�߳��j�8�?�aI<;��?78���g@}�~m9Wآ\آ\�5;��ӊ�@�pZ�9�Z$#�ɻd�qxq���O!�Od��%������g2��W2�U^�����d���:��K�7Iag��@���.���)�x�.yz-jڨ�A�Aw��%�H�_nT���ޢf��#Լ�wg��j�)�w�݃:r�s��y1�~�PK
    �z�H�����  �  *  QmxqwyzNypsgLRh/rhTgTBjWLOIYpLqT/Nul.class  �      �      �QMO�@}K>��n��@)�В҄�J��zh�!���@9g��n�78�TA�J��QU�	JUZ�ffw�y3��׷ ޡf������)�RS.��9�X0���3��V(C��!S��3d�#J��hߋC�0��0�����Z�9��<y2எCl2�ܖ�ʢ�%������<ǒ�6�a1�G�����/z:T��ɉ��#�]���Z&ڋ5�L�,(Xup)4O�����R$`����JH�z�_���%����|:��_\�\������q��>8��v�9m�~Dͳ:����(���xQ��\��
X�+��"ғ�ax�i0�t��g��_�rM푬=~�*!A�YXw�M�/C��S�[dn������Ã�C*2���/�ʄhfBT'�4g�!��oM`��v�8�qv���PK
    �z�H�,��  �  *  QmxqwyzNypsgLRh/rhTgTBjWLOIYpLqT/cOn.class  �      �      �Vk[S�~wr�sr<!P.
ȅ��0�Eq�f !��`HI����A[:2��~�^m�u�j[ڎә@kۧO?�CIE�ڹ9A��uN�Z��z��;����S���cpYЈo�p�����ю��[7�2��rs��.�e���p_��k�|���p�en���e�pZD/��7!�c���>��-���bx5�M�S1%R�>s"��)jt����tT��H89������˽_gx)J��I�ܦLRU�4��A�d��v/���D2�j"�*8�!�1��?��"Z�
��K
FqY�g�1�`��Tp��ŕG�G�"겞H�DL)p"�p�)j4��������Rb������WZ����Su5����zV�}E3����T���@��>��t��`�J{hV�=�PIe�g��]��q���tt%�z�TmUՈ-��:�(�Hk1�b&��^��wKV��M��3ϩ����wr%�'�h�e*���^6J7-&�kj����tU&�tD�d��v#��0I*�.sj�qa�����TQ�[|�E�ȸ�D�N��țA-�j�\��z��������>�c���Өx8�d��K��7�`����2�1o~��T=����Q8x��0'RU��Ȍlfx�T[qN�ওx�j*Ƈ�$�dԀf����!�8�㷌�<Bcbr����YԹgE�7e�»��y���凘Wt�_{w�][�um�:da:A�+Kk7o��[_���q�Ƃ�g㣡��͠72���NJ�E�yB�ȅD*���BZS��o�wЬ�.7[�l�]%oss����8��k����iT�c��%|�.Ś���������Z	�a�;�=nO���Q;�#�+�Tv{�O�=J�~�����z	?�qH9�h;Ra�K�	�oX{��~F�N��[�/����#�}��`��w]zu��u�M�QAl�X�~M�ƴ���Y����0B,�%�z�_������j�ڨ�?�0��1��tO��K��'ڟJ�#�=��\~��nà�����.zO4U���Ϸ��G/�g�'���"��Пn�^�[0���n{5k�q��Țz'*$�����c��'L���!Z�o����3gl>f��)�`i��%6i��I�i_Ϲ#}g=����ݗ>�nj�2��v��6h��C^o��l�E�z�4����Y|<�M�2�=��t����&��#�H.J�;�����$�ȇqt��f�r�fHh(C�%�V	}��8�}v���wԐ������TH��ww�>�E�L��	7��ѷ��"}��yl�C(��_��xB;�z����!q?u�����?*f��D5�ޫ�H�����>o"��Oyk�g��7�(;�+�y�pU��v��_����\'�*�I�n�Z���r���ۥ��i-ފ�1�!�o�x�P ��O{�>���͔S��a�䔨@���n��S����$����S�~�.�m;�5��?>�� ��Qo��S��}`����c��&��"ޅ9���>̩'f!=���A?z!Ը�Jw
*��jA%���:E��ǘ�U�Ѫ�,>+���b~��,�d�x�i!j�6�k�MshM�4�wӦ���q��l��O���	3s��i�o~�����bO�5s��@vs���AAg�]�ԗE(s���j����O��5���~�g�RO�s��Qڄ�nˍU�$�rr��m�d���m�C��3W�G0�-�pe�PK
    �z�H��t�_%  Z%     _023_/resources/icon_128x128.png  Z%      _%      Z%�ډPNG

   IHDR   �   �   �>a�   	pHYs    ��~�  
MiCCPPhotoshop ICC profile  xڝSwX��>��eVB��l� "#��Y�� a�@Ņ�
V�HUĂ�
H���(�gA��Z�U\8�ܧ�}z�����������y��&��j 9R�<:��OH�ɽ�H� ���g�  �yx~t�?��o  p�.$�����P&W  � �"��R �.T� � �S�d
 �  ly|B" � ��I> ة�� آ� � �(G$@� `U�R,�� ��@".���Y�2G�� v�X�@` ��B,�  8 C� L�0ҿ�_p��H �˕͗K�3���w����!��l�Ba)f	�"���#H�L�  ����8?������f�l��Ţ�k�o">!����� N���_���p��u�k�[ �V h��]3�	�Z
�z��y8�@��P�<
�%b��0�>�3�o��~��@��z� q�@������qanv�R���B1n��#�ǅ��)��4�\,��X��P"M�y�R�D!ɕ��2���	�w ��O�N���l�~��X�v @~�-�� g42y�  ����@+ ͗��  ��\��L�  D��*�A�������aD@$�<B�
��AT�:��������18��\��p`����	A�a!:�b��"���"aH4��� �Q"��r��Bj�]H#�-r9�\@���� 2����G1���Q�u@���Ơs�t4]���k��=�����K�ut }��c��1f��a\��E`�X&�c�X5V�5cX7v��a�$���^��l���GXLXC�%�#��W	��1�'"��O�%z��xb:��XF�&�!!�%^'_�H$ɒ�N
!%�2IIkH�H-�S�>�i�L&�m������ �����O�����:ň�L	�$R��J5e?���2B���Qͩ����:�ZIm�vP/S��4u�%͛Cˤ-��Кigi�h/�t�	݃E�З�k�����w���Hb(k{��/�L�ӗ��T0�2�g��oUX*�*|���:�V�~��TUsU?�y�T�U�^V}�FU�P�	��թU��6��RwR�P�Q_��_���c���F��H�Tc���!�2e�XB�rV�,k�Mb[���Lv�v/{LSCs�f�f�f��q�Ʊ��9ٜJ�!��{--?-��j�f�~�7�zھ�b�r�����up�@�,��:m:�u	�6�Q����u��>�c�y�	������G�m��������7046�l18c�̐c�k�i������h���h��I�'�&�g�5x>f�ob�4�e�k<abi2ۤĤ��)͔k�f�Ѵ�t���,ܬج��9՜k�a�ټ�����E��J�6�ǖږ|��M����V>VyV�V׬I�\�,�m�WlPW��:�˶�����v�m���)�)�Sn�1���
���9�a�%�m����;t;|rtu�vlp���4éĩ��Wgg�s��5�K���v�Sm���n�z˕��ҵ������ܭ�m���=�}��M.��]�=�A���X�q�㝧�����/^v^Y^��O��&��0m���[��{`:>=e���>�>�z�����"�=�#~�~�~���;�������y��N`������k��5��/>B	Yr�o���c3�g,����Z�0�&L�����~o��L�̶��Gl��i��})*2�.�Q�Stqt�,֬�Y�g��񏩌�;�j�rvg�jlRlc웸�����x��E�t$	�����=��s�l�3��T�tc��ܢ����˞w<Y5Y�|8����?� BP/O�nM򄛅OE����Q���J<��V��8�;}C�h�OFu�3	OR+y���#�MVD�ެ��q�-9�����Ri��+�0�(�Of++��y�m������#�s��l�Lѣ�R�PL/�+x[[x�H�HZ�3�f���#�|���P���ظxY��"�E�#�Sw.1]R�dxi��}�h˲��P�XRU�jy��R�ҥ�C+�W4�����n��Z�ca�dU�j��[V*�_�p�����F���WN_�|�ym���J����H��n��Y��J�jA�І����_mJ�t�zj��ʹ���5a5�[̶���6��z�]�V������&�ֿ�w{��;��켵+xWk�E}�n��ݏb���~ݸGwOŞ�{�{�E��jtolܯ���	mR6�H:p囀oڛ�w�pZ*�A��'ߦ|{�P������ߙ���Hy+�:�u�-�m�=���茣�^G���~�1�cu�5�W���(=��䂓�d���N?=ԙ�y�L��k]Q]�gCϞ?t�L�_�����]�p�"�b�%�K�=�=G~p��H�[o�e���W<�t�M�;����j��s���.]�y�����n&��%���v��w
�L�]z�x�����������e�m��`�`��Y�	�����Ӈ��G�G�#F#�����dΓ᧲���~V�y�s������K�X�����Ͽ�y��r﫩�:�#���y=�����}���ǽ�(�@�P���cǧ�O�>�|��/����%ҟ3    cHRM  z%  ��  ��  ��  u0  �`  :�  o�_�F  �IDATx��y�$Wu��ޛUo����#KhX�x�,�1`3K�`K�،#�`���@ava�@�6���x�`[�x���Z-��Rﯻ�{�˙?2�*�*���4��H���̬��}��s�=���*3y�5�� 3�`&3�dF���0�f�h��n��*<�v_�O<�+;\��B�������"u�1����W������p-���zB{O׽�s'�W��cO�*-�z�7������� ߜ��7`���X
�ڰ% _|�&�E�g� l���7�[ص�6��1h�H��� ϒW �mklk����N�ȇ.�{N{��щ��@�G�6��}5�vE� ~�g_�=�o�{�.����8�	����f6@}�X���VXnç�s�=6t����[ |Z��?#@uy9�K�4����Kr&"�R����<xÌ խ��2�t�����q�}���`�F1��o���Z��3�˯�5�x�y��E{`�-3�}��}� �rq��T�0QX�����Niڦ��6�~F�|yp^���w�t,|�����),$nᆁ�3.'�n��6r�m�]�ȫ�1�8��/��{�!2	�t��\Dn�.�]4�n�ҸJj��8�3���#�`���=�-�`6����S�� ��b޹�#+��Nt;�����>#@,�Ru�$	�v@bZ[�'<�G��9� ���_�5# �7�)i߽0B,�x6�O�y�ܹo��Y�A��<����vp�z2�2�׍m��_93t𜅇֜��}��g����L,�ع�^ [9��6��J���ĳ1uS�����쿜��n�4{}�c�?.%���!��_�4E��A�^ӊ`��ľk�F��-l�맘R�)����F�v��5�}#�K���w��]G��_iN'i�e��\�h"����+[M� ��`޽wI��&tf����?�$�l�(�� xs3e�:�������U�v�s9�X�-�F���x��A�F�2�+�1���~�#"�N����UW�n���-q7� W�����o�%m�L�t��c�b�Uو^_m򧮼���c��<29 �$F\�%�����+'��Bj�@��F�k��M$���?�ꠛ��F�`Vc�_	{a�ƠO����wEb|_i�p�t]۳dxTI����s�:<.��>P���E�O�/Ϩ�����CA��IY�2L#�5�ݷd�6�d _�7/J����y��:Z�0N2�̘��>h��=gZ�C��-��2���)�z܌d�ye_!��"AlJƵDX���\������Q�p맅�H0ONv��D��^U~e�l<n  N�cG�
#D���o�{�/�n�l���{z	��YI ���4�l��RǛ��8�%����������z��*�$���
��� �DxQy��z������/'�1�1�<��Z$����$x�F��f��ƴ6v���%��_s2������"�xb��đ�p�Fl{�����M���� )cG��:!Y$8�Qd�F����̡n������ۚ$��8��� �e�-��u�,�6d��&ED����[m����RԪQl�)�S!CL�� ?t6�m��y�Λ��S��
ܿ<"t��Gu�7O�J�ML;#h�KB�����yMج�Ds� �Dp��}��e/�Dy��X�f*���i���$�di^?I~`�¼Q����uȷ��2��������J��x��F�r([#6y��8@Dh{rK��k#�+�?��Sà���xQɔ0��J��L��H5��A�|�+�Ww�a�o�u⹕�o'�F��n�1��j�4 �dBj�I ������-�z���r�A�T5�bPuJ��i
B��cb�K��xx�l4��"A,7 ϝ� ji^� �����b$Cۏ�Ś�2�����6��]�x�P�R�i^:��>Z�yt�yf`�H6,�{��jN���]�x}����ܪ5յi�*d����u�,#��5|pHM�����ߴi⦿3|��&q'!��Bq�W!tZ�{3K��h4ڒ�
���S�Yn�8{��%�6� �Vi|�*$�c��ל'���� N�"�?ᢞg0��+��.yq1�&q ��7����Ժ�&Aq����5�����A�U7׸���%v �eh߼Y�jT_U�J/굞(��� X����j<��]g��%r�N� ��4/-����"Cj�+����~jx؏i��_?��N\r�H��4/���j$�j�R�Zޮ���Pw6ɵ�+��r�`Gb!׎�4!A3�@�>��U>:�ο��,#��}�`<�+Ch�tJD�l�i�T�
7��W�+����� OO\��^@%]q���}jM��e.��F?��*1���n��ax�Td�˯�f��V����$`̭�9�\D:��J�fj�)~���i��� ?�����$i��*�B{_���_-!A�6�ݿз|7�R��AT���0F�u�L���c+]N��t�UmNՍ��/WV� ��ϑN�҆$���jw��K|C�w�p��붜|����U!�ӫ'N�[�Y9�ލPݤ��Ո�J�BS��ɍ��4�1i���k�\$M����y�[;KO��9]���WSf+�Q����3��a���!��!ր�-��y��6�ld��k��ɼl��K����H��\%�m�F�3ˌ >��A%z/ 	��s�^�%�>����
"r_�s�P�*2nDF@*�~�z7>��<�Ƞ.��{����\܎pM�i� �t�xƮ3����.���	�X��F���������N<���U�I��EE:�Ş�|��W)x�ŧR�?������J�kW����i��+�~�����.�&	�*���3az�9vLD���Y����SOD\���=~)���2��9�e�����h+�-t��zU��A#�Ěaݏ���bd��K���NT!�  <m!i��7�_ڛX��c�DD�
�cϢ��?�B����8τ�	���k�����9�%��m#b1F�6��n��*�M�Dt�x����0TTI�?Re:�@�4�*��7�tӆ$�X"�:���^��Dm��4�w��`� Ar;c[�`%�H����/�}1g�����~��ª��1PA� ��Ț��&���{�a~__�`��N���?-�>�+2;B�kN3o^�a�D�gT_Gl�%�Qw
���tv���AM��j�4z�в]u���/b��q���\��������F�F���I*����n��!AЋ3�!No�������b;�_����#���	/��M�?T�����<��t�an�N:�_�[}Ꝇ��	e��$�2�V�}�)���c-��I�9�u�Hmo�1#{�P��m/#}�q$2�#��?P�(��5ikx2��f�x"�����M����i׮u�y,}������l�q?��=D�������w{v����\z�}��b���0�iu���}�a7(Ak��$"����<�x%T�.&x/p�P}Mg~��p�9$:�n�/���5��}�-����
5#�@�m��`��{��A���_�x+D8Ę{��Wk\��q��j.�1"c�A����8Z!"c��0n7�G���4^ �!�8A%T�F�Mu������w_��}��[y
X������W�b%��O�ӻ_��:x��2���ak9��=�F�t<� �Da�?$"�=
�<���-<n���!�a2>���$�p"H�K[+�qG.__���i�3P�CF�t����	���k�ڑ+x��a���[__�Ԝ+SR�U�2��{+~H�	��C����Wr-�Sοs��p�X_��O$�6%��}���{�_�ws{vb�N��PL�a {�P5LT�ö+��p�9B8�/��:�/^�Q~����e���#5�L��?�h�5|Ekh��s��.X+Xgp�a�������y7pyF1�z$hJ���PP��=v����x�L�$��J\�%1��"(bU@h�"�k���qj[���"����p�~�*�ZN�=�����7���."��������o���#}M��vj�Ҥ���+=�J����jr��g�t��Xc�Z��>�O�����Ѕ�xp��d|�V��(�!΅�]/�X�Z�N`Ԡa��A5q��&�kP���
Ƶ�D�]V���,�N芿��_�<�MU,a1�d,�]S-��f�~���Ё�E(�^����҄q��y���#��l��Қ�R����[�r�ȭ��}mhN\ܢ������Gf���`�b��=���=���ߨ��n��\X�ΏU�a�'�7����� �ݑ4c1�*���'������$�)�����1������C?bp~ߨ�(J��ı��m��X����-?����!-0P�6�o� W�����6J3vTU�x�w���H.����Q;
Rp*��@���dm�Ä�$U"��l�i�_k��毚��b2}_��ĳ�}��ċ �j$� ��fNVl�]�{��o��S.O2��*�^��*&(�:)�k6���J�a��J2Q�iW���b2B��ᨍZ\�g�zQ��_P�x�/c��%[s�]���^y;p��:�j�XԮ�<׷�/sx݊�ߌ�o�BB
�Q.��S��&D"���Wq�t�� !�]Z^k0���J{�"��_1��ٲ?�a����3�巁{�u]"h���UoϋCs�"��~)���̕�O�ŧ�C��>�c�Ռ{na��]J�fdP�Ŭ<.����a��#߰�������TQ�-��S����H�ͫ2�ָ3�K�l�/j�N�۱�p8����z������ig��C�<Rj�h���:���ӆ4h΄�|4닼�!�oAկl�S�9+�����w�
�v��H����kb{�o��i�h�;�)LA�8�n�H�yX���u �O��*�_��d�%���B�;�	*&^�8��SQ?1�~A�b���Y�^��8�1��Z�f�>�����űe��c�P��B�J�7ǷȮ�\�cOvj���ý4$k�A��^nUZ���m�j�+��en��8�pk���2<H/�n|0�b]�cV��q�6)����X�[D��D���&G��Q�P�"�U�&d���
����?0���U�WA%P�?�3�9��3��<�nF���A���ׇ�[��g:���J�b����e%��$�[*�M�i�o�%z�xr��ʪ[#��ӏ b<�댁_�ċ��g�C� e�O��ˀ�&�poV��Z-���n��dd�����*A�b���o��uK��ݾ2	* �����uR���wY弪%bB���ȫU��Ԯ��"p�<ݩK'z��al�u@d�d9�
I0��V��Fzc�i��V�ZM3H������	�f����øN��,%AZ�7jom�2KT��ڳ%�>�ߪwW��A���z%V2���nߋB����;�M��������I0F�2/0�w-?O�ke::`?��ii��-T�x�O�B�/�[{^l�tc�����b2�S��I��1?�5#,>��z��+Z���If����JfrP�[6����H֗& +�Ӷ:)�+8�H0����ȱ6��EdG����&��[X2דe�٣�����zj�w3����>�Z���!�RX���2�r3�VO�N�O�
�=�7� ����l���w�$D��i^��\D��9��+�I%��C��,�jj���eހN���'��7�)z����T�kx��K=uk�O�P0�:7�ˏ�8�I��6K�
�������8�G+TF�'@�����jݬ��A��k&H��+b\�������
$(!B�wU�_	�&CY~�O>�AI�#4@O��ZS��jk�F��N�ߏ��p����Z��%�IT���WQ4_%h!�Z���؅�[� 8黃c���!���]�8���Ъ[�+��k� �2��VwٛJ+�����R�O�8��ꦆ��|��
���� �[�)�0�$���C׫�	�Ю���O�<U���HPEhQW-!E%��d�o2$���h�x�F`�-�2���#�
�G��Ԯ�F��?���UT'y hi�O�������n�������J���/d~,����Tb�����ն�e,�n�Z�����r���h�f�������A�񵅩��w��=�D�f�-a[����b�{S��� 5�viy%V��^����G���7� �K"���Y� h��1��+�u�[.Gd
$�%�4�e3�L�K�J/Qz����BL�����v�����L��=�D�v�3s�o���khi+5ykD���2�����Q��֏�o���*Dfw����[;?�q��ѽ
�3e>u��3����_3A��%�F�~�rS�x�f�P�{���ww�uXqmШ^��V#{^�!W�ݕG�&Ғ!�������
�m'լ��z�*ڧ���5����)Y�U,��4�QZ2$Z��J̝��)�SE��m��b�v���T�Xe�t9)I�$J*���EC��zǏ���L����ߦ�Zkryߧ���hUءgM7[eh�|�# ��l��L6U̬	f�Ɍ 3�`&3�dF���0�G��MI���Р    IEND�B`�PK
    �z�H!�uJ�   �    _023_/resources/manifest.json  �      �       ]�ъ�0E��a�c)�V+����_��Hɦ���NB�E�w�V�@`&�ܛIn���H�ȶ���>u_V�v�Y��3Z�4El]�����j×�j"zA���/��������i1d��Za5༎U��U�Y��<�E�	�tB"�nRAv!�6�ϳe���T��67tbr�m�\/����q,�m�"+�d<��4Q=���m��^�����1i�~]�V��Cwx�t�|�PK
    �z�H��X�6   7     _023_/resources/panel.json  7       6       ���R �� %+����+}�Ԋ�܂�Ԃ��Ԕ��̒T��T�ĂL=��/W- PK
     �z�H               META-INF/services/PK
    �z�H�7S&   $     META-INF/services/module.Server  $       &       ̭(,���,(N�	��+�Iq�
����,�)��+� PK
     �z�H            	         �A    META-INF/��  PK
     �z�H                      �A+   QmxqwyzNypsgLRh/PK
     �z�H            !          �AY   QmxqwyzNypsgLRh/rhTgTBjWLOIYpLqT/PK
     �z�H                      �A�   _023_/PK
     �z�H                      �A�   _023_/resources/PK
    �z�HK^t
  +  *           ���   QmxqwyzNypsgLRh/rhTgTBjWLOIYpLqT/Con.classPK
    �z�H�����  �  *           ��S  QmxqwyzNypsgLRh/rhTgTBjWLOIYpLqT/Nul.classPK
    �z�H�,��  �  *           ��\  QmxqwyzNypsgLRh/rhTgTBjWLOIYpLqT/cOn.classPK
    �z�H��t�_%  Z%              ���  _023_/resources/icon_128x128.pngPK
    �z�H!�uJ�   �             ��Q:  _023_/resources/manifest.jsonPK
    �z�H��X�6   7              ���;  _023_/resources/panel.jsonPK
     �z�H                      �A
<  META-INF/services/PK
    �z�H�7S&   $              ��:<  META-INF/services/module.ServerPK      �  �<    